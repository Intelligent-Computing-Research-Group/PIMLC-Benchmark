module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 ;
  assign n262 = x8 & x9 ;
  assign n254 = ~x4 ;
  assign n48 = n254 & n262 ;
  assign n255 = ~x5 ;
  assign n349 = n255 & x8 ;
  assign n350 = x14 | x15 ;
  assign n25 = x13 | n350 ;
  assign n26 = x12 | n25 ;
  assign n27 = x11 | n26 ;
  assign n256 = ~x7 ;
  assign n28 = n256 & x10 ;
  assign n29 = n27 | n28 ;
  assign n30 = n255 & n262 ;
  assign n31 = n29 | n30 ;
  assign n32 = n256 & x9 ;
  assign n33 = x10 | n27 ;
  assign n34 = n32 | n33 ;
  assign n257 = ~n34 ;
  assign n35 = x8 & n257 ;
  assign n258 = ~n35 ;
  assign n36 = x6 & n258 ;
  assign n37 = x9 | n349 ;
  assign n259 = ~n36 ;
  assign n38 = n259 & n37 ;
  assign n39 = n31 | n38 ;
  assign n260 = ~x6 ;
  assign n276 = n260 & n262 ;
  assign n40 = n276 & n257 ;
  assign n261 = ~n40 ;
  assign n41 = n39 & n261 ;
  assign n22 = ~n41 ;
  assign n43 = n349 & n22 ;
  assign n42 = x8 & n22 ;
  assign n263 = ~n42 ;
  assign n44 = x5 & n263 ;
  assign n45 = n43 | n44 ;
  assign n46 = n254 & x8 ;
  assign n47 = x9 | n46 ;
  assign n264 = ~n45 ;
  assign n49 = n264 & n47 ;
  assign n50 = n48 | n49 ;
  assign n265 = ~n31 ;
  assign n51 = n265 & n37 ;
  assign n266 = ~n51 ;
  assign n52 = n36 & n266 ;
  assign n53 = n40 & n51 ;
  assign n54 = n52 | n53 ;
  assign n267 = ~x10 ;
  assign n55 = n267 & n54 ;
  assign n268 = ~n29 ;
  assign n56 = x10 & n268 ;
  assign n57 = n39 & n56 ;
  assign n58 = n55 | n57 ;
  assign n269 = ~n50 ;
  assign n65 = n269 & n58 ;
  assign n270 = ~n54 ;
  assign n59 = x10 & n270 ;
  assign n60 = n50 | n59 ;
  assign n271 = ~n55 ;
  assign n61 = n271 & n60 ;
  assign n287 = x7 & x11 ;
  assign n272 = ~n26 ;
  assign n62 = n287 & n272 ;
  assign n273 = ~n62 ;
  assign n63 = n27 & n273 ;
  assign n64 = n61 | n63 ;
  assign n66 = n54 & n64 ;
  assign n67 = n65 | n66 ;
  assign n94 = n61 & n62 ;
  assign n68 = n256 & n26 ;
  assign n274 = ~x3 ;
  assign n76 = n274 & n262 ;
  assign n275 = ~n57 ;
  assign n69 = n275 & n64 ;
  assign n21 = ~n69 ;
  assign n70 = x8 & n21 ;
  assign n277 = ~n70 ;
  assign n71 = x4 & n277 ;
  assign n72 = n46 & n21 ;
  assign n73 = n71 | n72 ;
  assign n74 = n274 & x8 ;
  assign n75 = x9 | n74 ;
  assign n278 = ~n73 ;
  assign n77 = n278 & n75 ;
  assign n78 = n76 | n77 ;
  assign n80 = x10 | n78 ;
  assign n79 = x10 & n78 ;
  assign n279 = ~n48 ;
  assign n81 = n47 & n279 ;
  assign n82 = n21 & n81 ;
  assign n280 = ~n82 ;
  assign n83 = n45 & n280 ;
  assign n84 = n264 & n82 ;
  assign n85 = n83 | n84 ;
  assign n281 = ~n79 ;
  assign n86 = n281 & n85 ;
  assign n282 = ~n86 ;
  assign n87 = n80 & n282 ;
  assign n88 = x11 & n87 ;
  assign n91 = n25 | n88 ;
  assign n90 = x11 | n87 ;
  assign n283 = ~n67 ;
  assign n92 = n283 & n90 ;
  assign n93 = n91 | n92 ;
  assign n95 = n68 | n93 ;
  assign n284 = ~n94 ;
  assign n96 = n284 & n95 ;
  assign n285 = ~x11 ;
  assign n89 = n285 & n87 ;
  assign n286 = ~n87 ;
  assign n99 = x11 & n286 ;
  assign n100 = n89 | n99 ;
  assign n20 = ~n96 ;
  assign n101 = n20 & n100 ;
  assign n102 = n67 & n101 ;
  assign n103 = n67 | n101 ;
  assign n288 = ~n102 ;
  assign n104 = n288 & n103 ;
  assign n325 = n256 & x13 ;
  assign n136 = n325 | n350 ;
  assign n289 = ~x2 ;
  assign n108 = n289 & n262 ;
  assign n97 = n74 & n20 ;
  assign n98 = x8 & n20 ;
  assign n290 = ~n98 ;
  assign n105 = x3 & n290 ;
  assign n106 = n97 | n105 ;
  assign n302 = n289 & x8 ;
  assign n107 = x9 | n302 ;
  assign n291 = ~n106 ;
  assign n109 = n291 & n107 ;
  assign n110 = n108 | n109 ;
  assign n111 = x10 | n110 ;
  assign n292 = ~n76 ;
  assign n112 = n75 & n292 ;
  assign n113 = n20 & n112 ;
  assign n114 = n278 & n113 ;
  assign n293 = ~n113 ;
  assign n115 = n73 & n293 ;
  assign n116 = n114 | n115 ;
  assign n117 = x10 & n110 ;
  assign n294 = ~n117 ;
  assign n118 = n116 & n294 ;
  assign n295 = ~n118 ;
  assign n119 = n111 & n295 ;
  assign n120 = x11 & n119 ;
  assign n121 = x11 | n119 ;
  assign n122 = n80 & n20 ;
  assign n123 = n86 & n122 ;
  assign n124 = n281 & n122 ;
  assign n125 = n85 | n124 ;
  assign n296 = ~n123 ;
  assign n126 = n296 & n125 ;
  assign n297 = ~n126 ;
  assign n127 = n121 & n297 ;
  assign n128 = n120 | n127 ;
  assign n129 = x12 & n128 ;
  assign n298 = ~n129 ;
  assign n130 = n104 & n298 ;
  assign n131 = x7 & n93 ;
  assign n299 = ~x13 ;
  assign n132 = x12 & n299 ;
  assign n133 = n131 & n132 ;
  assign n134 = x12 | n128 ;
  assign n300 = ~n133 ;
  assign n135 = n300 & n134 ;
  assign n301 = ~n130 ;
  assign n137 = n301 & n135 ;
  assign n138 = n136 | n137 ;
  assign n147 = n298 & n134 ;
  assign n19 = ~n138 ;
  assign n148 = n19 & n147 ;
  assign n303 = ~n104 ;
  assign n149 = n303 & n148 ;
  assign n304 = ~n148 ;
  assign n150 = n104 & n304 ;
  assign n151 = n149 | n150 ;
  assign n305 = ~x15 ;
  assign n143 = n305 & n131 ;
  assign n144 = n26 & n143 ;
  assign n306 = ~x14 ;
  assign n145 = n306 & n144 ;
  assign n146 = n137 & n145 ;
  assign n152 = x8 & n19 ;
  assign n153 = n289 & n152 ;
  assign n307 = ~n152 ;
  assign n154 = x2 & n307 ;
  assign n155 = n153 | n154 ;
  assign n308 = ~x1 ;
  assign n156 = n308 & x8 ;
  assign n157 = x9 | n156 ;
  assign n309 = ~n155 ;
  assign n158 = n309 & n157 ;
  assign n159 = n308 & n262 ;
  assign n160 = n158 | n159 ;
  assign n161 = x10 | n160 ;
  assign n310 = ~n108 ;
  assign n162 = n107 & n310 ;
  assign n163 = n19 & n162 ;
  assign n164 = n291 & n163 ;
  assign n311 = ~n163 ;
  assign n165 = n106 & n311 ;
  assign n166 = n164 | n165 ;
  assign n167 = x10 & n160 ;
  assign n312 = ~n167 ;
  assign n168 = n166 & n312 ;
  assign n313 = ~n168 ;
  assign n169 = n161 & n313 ;
  assign n170 = x11 | n169 ;
  assign n171 = x11 & n169 ;
  assign n172 = n111 & n19 ;
  assign n174 = n118 & n172 ;
  assign n173 = n294 & n172 ;
  assign n175 = n116 | n173 ;
  assign n314 = ~n174 ;
  assign n176 = n314 & n175 ;
  assign n315 = ~n171 ;
  assign n177 = n315 & n176 ;
  assign n316 = ~n177 ;
  assign n178 = n170 & n316 ;
  assign n179 = x12 | n178 ;
  assign n180 = x12 & n178 ;
  assign n317 = ~n120 ;
  assign n181 = n317 & n121 ;
  assign n182 = n19 & n181 ;
  assign n183 = n126 & n182 ;
  assign n184 = n126 | n182 ;
  assign n318 = ~n183 ;
  assign n185 = n318 & n184 ;
  assign n319 = ~n180 ;
  assign n186 = n319 & n185 ;
  assign n320 = ~n186 ;
  assign n187 = n179 & n320 ;
  assign n189 = x13 | n187 ;
  assign n321 = ~n151 ;
  assign n190 = n321 & n189 ;
  assign n188 = x13 & n187 ;
  assign n322 = ~n143 ;
  assign n191 = n350 & n322 ;
  assign n192 = n188 | n191 ;
  assign n193 = n190 | n192 ;
  assign n323 = ~n146 ;
  assign n194 = n323 & n193 ;
  assign n324 = ~n188 ;
  assign n239 = n324 & n189 ;
  assign n18 = ~n194 ;
  assign n240 = n18 & n239 ;
  assign n241 = n321 & n240 ;
  assign n326 = ~n240 ;
  assign n242 = n151 & n326 ;
  assign n243 = n241 | n242 ;
  assign n327 = ~n243 ;
  assign n244 = x14 & n327 ;
  assign n328 = ~n131 ;
  assign n248 = x15 & n328 ;
  assign n249 = n244 | n248 ;
  assign n196 = n161 & n312 ;
  assign n197 = n18 & n196 ;
  assign n198 = n166 | n197 ;
  assign n199 = n166 & n197 ;
  assign n329 = ~n199 ;
  assign n200 = n198 & n329 ;
  assign n330 = ~n200 ;
  assign n219 = x11 & n330 ;
  assign n331 = ~x0 ;
  assign n208 = n331 & n262 ;
  assign n202 = x8 & n18 ;
  assign n203 = n308 & n202 ;
  assign n332 = ~x9 ;
  assign n205 = x0 & n332 ;
  assign n204 = n308 & n157 ;
  assign n206 = n202 | n204 ;
  assign n333 = ~n205 ;
  assign n207 = n333 & n206 ;
  assign n334 = ~n203 ;
  assign n209 = n334 & n207 ;
  assign n210 = n208 | n209 ;
  assign n212 = x10 | n210 ;
  assign n211 = x10 & n210 ;
  assign n335 = ~n159 ;
  assign n213 = n157 & n335 ;
  assign n214 = n18 & n213 ;
  assign n215 = n309 & n214 ;
  assign n336 = ~n214 ;
  assign n216 = n155 & n336 ;
  assign n217 = n215 | n216 ;
  assign n337 = ~n211 ;
  assign n218 = n337 & n217 ;
  assign n338 = ~n218 ;
  assign n220 = n212 & n338 ;
  assign n221 = n219 | n220 ;
  assign n201 = n285 & n200 ;
  assign n222 = n170 & n315 ;
  assign n223 = n18 & n222 ;
  assign n224 = n176 | n223 ;
  assign n225 = n176 & n223 ;
  assign n339 = ~n225 ;
  assign n226 = n224 & n339 ;
  assign n340 = ~x12 ;
  assign n227 = n340 & n226 ;
  assign n228 = n201 | n227 ;
  assign n341 = ~n228 ;
  assign n229 = n221 & n341 ;
  assign n230 = n179 & n319 ;
  assign n231 = n18 & n230 ;
  assign n342 = ~n185 ;
  assign n232 = n342 & n231 ;
  assign n343 = ~n231 ;
  assign n233 = n185 & n343 ;
  assign n234 = n232 | n233 ;
  assign n344 = ~n234 ;
  assign n235 = x13 & n344 ;
  assign n345 = ~n226 ;
  assign n236 = x12 & n345 ;
  assign n237 = n235 | n236 ;
  assign n238 = n229 | n237 ;
  assign n245 = n299 & n234 ;
  assign n246 = n306 & n243 ;
  assign n247 = n245 | n246 ;
  assign n346 = ~n247 ;
  assign n250 = n238 & n346 ;
  assign n251 = n249 | n250 ;
  assign n195 = n138 & n144 ;
  assign n252 = n194 & n195 ;
  assign n347 = ~n252 ;
  assign n253 = n251 & n347 ;
  assign n348 = n260 & x8 ;
  assign n142 = n348 | n34 ;
  assign n139 = n256 & x8 ;
  assign n140 = x9 | n139 ;
  assign n141 = n33 | n140 ;
  assign n17 = ~n253 ;
  assign n23 = ~n142 ;
  assign n24 = ~n141 ;
  assign y0 = n17 ;
  assign y1 = n18 ;
  assign y2 = n19 ;
  assign y3 = n20 ;
  assign y4 = n21 ;
  assign y5 = n22 ;
  assign y6 = n23 ;
  assign y7 = n24 ;
endmodule
