module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 ;
  assign n29877 = x14 & x15 ;
  assign n37294 = x14 | x15 ;
  assign n30013 = ~n29877 ;
  assign n37297 = n30013 & n37294 ;
  assign n29898 = x16 & x17 ;
  assign n37298 = x16 | x17 ;
  assign n30014 = ~n29898 ;
  assign n37299 = n30014 & n37298 ;
  assign n37300 = n37297 & n37299 ;
  assign n37301 = x5 | x6 ;
  assign n65 = x7 | n37301 ;
  assign n29880 = x5 & x6 ;
  assign n30015 = ~n29880 ;
  assign n67 = n30015 & n37301 ;
  assign n30016 = ~n37301 ;
  assign n66 = x7 & n30016 ;
  assign n30017 = ~x7 ;
  assign n68 = n30017 & n29880 ;
  assign n69 = n66 | n68 ;
  assign n70 = n67 | n69 ;
  assign n71 = x8 & n70 ;
  assign n30018 = ~n71 ;
  assign n72 = n65 & n30018 ;
  assign n73 = x24 | x25 ;
  assign n30019 = ~x26 ;
  assign n74 = x23 & n30019 ;
  assign n30020 = ~n73 ;
  assign n75 = n30020 & n74 ;
  assign n30021 = ~x28 ;
  assign n76 = x27 & n30021 ;
  assign n77 = x29 | x30 ;
  assign n30022 = ~n77 ;
  assign n79 = n76 & n30022 ;
  assign n80 = n75 & n79 ;
  assign n30023 = ~x30 ;
  assign n81 = x29 & n30023 ;
  assign n82 = n76 & n81 ;
  assign n83 = n75 & n82 ;
  assign n30024 = ~x29 ;
  assign n84 = n30024 & x30 ;
  assign n86 = n76 & n84 ;
  assign n30025 = ~x25 ;
  assign n87 = x24 & n30025 ;
  assign n88 = x23 | x26 ;
  assign n30026 = ~n88 ;
  assign n89 = n87 & n30026 ;
  assign n90 = n86 & n89 ;
  assign n91 = n83 | n90 ;
  assign n92 = n80 | n91 ;
  assign n30027 = ~x27 ;
  assign n93 = n30027 & x28 ;
  assign n94 = n81 & n93 ;
  assign n30028 = ~x24 ;
  assign n95 = n30028 & x25 ;
  assign n96 = n74 & n95 ;
  assign n97 = n94 & n96 ;
  assign n98 = x27 | x28 ;
  assign n30029 = ~n98 ;
  assign n99 = n84 & n30029 ;
  assign n30030 = ~x23 ;
  assign n100 = n30030 & x26 ;
  assign n101 = n95 & n100 ;
  assign n103 = n99 & n101 ;
  assign n104 = n97 | n103 ;
  assign n105 = n87 & n100 ;
  assign n107 = n79 & n105 ;
  assign n29900 = x29 & x30 ;
  assign n109 = n29900 & n93 ;
  assign n110 = n74 & n87 ;
  assign n112 = n109 & n110 ;
  assign n113 = n107 | n112 ;
  assign n114 = x23 | n73 ;
  assign n30031 = ~n114 ;
  assign n115 = x26 & n30031 ;
  assign n116 = n79 & n115 ;
  assign n117 = n113 | n116 ;
  assign n118 = n104 | n117 ;
  assign n119 = n92 | n118 ;
  assign n120 = n29900 & n76 ;
  assign n29910 = x24 & x25 ;
  assign n122 = x23 & n29910 ;
  assign n123 = x26 & n122 ;
  assign n124 = n120 & n123 ;
  assign n125 = n29900 & n30029 ;
  assign n126 = n75 & n125 ;
  assign n127 = n84 & n93 ;
  assign n29911 = x23 & x24 ;
  assign n128 = n30025 & x26 ;
  assign n129 = n29911 & n128 ;
  assign n130 = n127 & n129 ;
  assign n131 = n126 | n130 ;
  assign n132 = n30026 & n95 ;
  assign n133 = n94 & n132 ;
  assign n134 = n131 | n133 ;
  assign n135 = n124 | n134 ;
  assign n136 = n29910 & n30026 ;
  assign n138 = n109 & n136 ;
  assign n139 = n86 & n96 ;
  assign n140 = n138 | n139 ;
  assign n137 = n75 | n136 ;
  assign n141 = n99 & n137 ;
  assign n142 = n77 | n98 ;
  assign n143 = n73 | n88 ;
  assign n145 = n142 | n143 ;
  assign n30032 = ~n141 ;
  assign n146 = n30032 & n145 ;
  assign n30033 = ~n140 ;
  assign n147 = n30033 & n146 ;
  assign n30034 = ~n135 ;
  assign n148 = n30034 & n147 ;
  assign n30035 = ~n119 ;
  assign n149 = n30035 & n148 ;
  assign n150 = n79 & n123 ;
  assign n151 = n79 & n110 ;
  assign n152 = n150 | n151 ;
  assign n30007 = x27 & x28 ;
  assign n154 = n30007 & n84 ;
  assign n155 = x23 & n30028 ;
  assign n156 = n128 & n155 ;
  assign n157 = n154 & n156 ;
  assign n158 = n82 & n129 ;
  assign n159 = n96 & n99 ;
  assign n160 = n158 | n159 ;
  assign n161 = n157 | n160 ;
  assign n162 = n125 & n129 ;
  assign n163 = n89 & n120 ;
  assign n164 = n162 | n163 ;
  assign n165 = n161 | n164 ;
  assign n166 = n152 | n165 ;
  assign n167 = n101 & n120 ;
  assign n30036 = ~n143 ;
  assign n168 = n94 & n30036 ;
  assign n169 = n81 & n30029 ;
  assign n171 = n75 & n169 ;
  assign n172 = n168 | n171 ;
  assign n173 = n167 | n172 ;
  assign n174 = n105 & n127 ;
  assign n175 = n29900 & n30007 ;
  assign n176 = n105 & n175 ;
  assign n177 = n174 | n176 ;
  assign n37283 = x25 & x26 ;
  assign n178 = n37283 & n155 ;
  assign n179 = n127 & n178 ;
  assign n180 = n30022 & n93 ;
  assign n181 = n136 & n180 ;
  assign n182 = n179 | n181 ;
  assign n183 = n177 | n182 ;
  assign n184 = n173 | n183 ;
  assign n30037 = ~n142 ;
  assign n185 = n115 & n30037 ;
  assign n186 = n178 & n180 ;
  assign n187 = n154 & n178 ;
  assign n188 = n186 | n187 ;
  assign n189 = n185 | n188 ;
  assign n190 = n110 & n120 ;
  assign n191 = n30019 & n29910 ;
  assign n192 = n30007 & n30022 ;
  assign n194 = n191 & n192 ;
  assign n195 = n30030 & n194 ;
  assign n196 = n190 | n195 ;
  assign n197 = n189 | n196 ;
  assign n198 = n184 | n197 ;
  assign n199 = n123 & n154 ;
  assign n200 = n86 & n132 ;
  assign n201 = n199 | n200 ;
  assign n202 = n127 & n156 ;
  assign n203 = n75 & n86 ;
  assign n204 = n202 | n203 ;
  assign n205 = n115 & n125 ;
  assign n206 = n204 | n205 ;
  assign n207 = n201 | n206 ;
  assign n208 = n29910 & n74 ;
  assign n212 = n154 & n208 ;
  assign n213 = n30007 & n81 ;
  assign n214 = n105 & n213 ;
  assign n215 = n212 | n214 ;
  assign n216 = n105 & n180 ;
  assign n217 = n79 & n208 ;
  assign n218 = n216 | n217 ;
  assign n219 = n215 | n218 ;
  assign n220 = n156 & n175 ;
  assign n221 = n156 & n169 ;
  assign n222 = n220 | n221 ;
  assign n223 = n96 & n125 ;
  assign n224 = n169 & n178 ;
  assign n225 = n223 | n224 ;
  assign n226 = n222 | n225 ;
  assign n227 = n219 | n226 ;
  assign n228 = n207 | n227 ;
  assign n229 = n198 | n228 ;
  assign n230 = n166 | n229 ;
  assign n30038 = ~n230 ;
  assign n231 = n149 & n30038 ;
  assign n232 = n125 & n178 ;
  assign n233 = n109 & n115 ;
  assign n234 = n232 | n233 ;
  assign n235 = n75 & n30037 ;
  assign n236 = n99 & n105 ;
  assign n237 = n235 | n236 ;
  assign n238 = n234 | n237 ;
  assign n239 = n115 & n127 ;
  assign n240 = n94 & n101 ;
  assign n241 = n110 & n175 ;
  assign n242 = n240 | n241 ;
  assign n243 = n239 | n242 ;
  assign n244 = n96 & n175 ;
  assign n245 = n175 & n178 ;
  assign n247 = n244 | n245 ;
  assign n248 = n82 & n30036 ;
  assign n249 = n178 & n192 ;
  assign n250 = n248 | n249 ;
  assign n251 = n247 | n250 ;
  assign n252 = n243 | n251 ;
  assign n253 = n127 & n30036 ;
  assign n254 = n86 & n191 ;
  assign n255 = x23 & n254 ;
  assign n256 = n253 | n255 ;
  assign n257 = n79 & n132 ;
  assign n258 = n79 & n129 ;
  assign n259 = n30030 & x24 ;
  assign n261 = n37283 & n259 ;
  assign n263 = n86 & n261 ;
  assign n264 = n258 | n263 ;
  assign n265 = n257 | n264 ;
  assign n266 = n256 | n265 ;
  assign n267 = n252 | n266 ;
  assign n268 = n238 | n267 ;
  assign n269 = n82 & n101 ;
  assign n270 = n75 & n127 ;
  assign n271 = n269 | n270 ;
  assign n272 = n89 & n154 ;
  assign n273 = n125 & n132 ;
  assign n274 = n272 | n273 ;
  assign n275 = n271 | n274 ;
  assign n276 = n89 & n175 ;
  assign n277 = n175 & n261 ;
  assign n278 = n276 | n277 ;
  assign n279 = n120 & n156 ;
  assign n280 = n125 & n261 ;
  assign n281 = n279 | n280 ;
  assign n282 = n110 & n180 ;
  assign n283 = n75 & n94 ;
  assign n285 = n282 | n283 ;
  assign n286 = n281 | n285 ;
  assign n287 = n278 | n286 ;
  assign n288 = n275 | n287 ;
  assign n289 = n105 & n120 ;
  assign n290 = n86 & n123 ;
  assign n291 = n289 | n290 ;
  assign n292 = n99 & n115 ;
  assign n293 = n109 & n132 ;
  assign n294 = n292 | n293 ;
  assign n295 = n291 | n294 ;
  assign n296 = n127 & n261 ;
  assign n297 = n169 & n191 ;
  assign n298 = x23 & n297 ;
  assign n299 = n296 | n298 ;
  assign n300 = n120 & n129 ;
  assign n301 = n89 & n99 ;
  assign n302 = n129 & n169 ;
  assign n303 = n301 | n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = n299 | n304 ;
  assign n306 = n295 | n305 ;
  assign n307 = n288 | n306 ;
  assign n308 = n268 | n307 ;
  assign n309 = n79 & n96 ;
  assign n310 = n105 & n30037 ;
  assign n311 = n309 | n310 ;
  assign n312 = n89 & n30037 ;
  assign n313 = n82 & n156 ;
  assign n314 = n86 & n178 ;
  assign n315 = n313 | n314 ;
  assign n316 = n312 | n315 ;
  assign n317 = n311 | n316 ;
  assign n318 = n125 & n208 ;
  assign n319 = n132 & n213 ;
  assign n320 = n110 & n154 ;
  assign n321 = n319 | n320 ;
  assign n322 = n318 | n321 ;
  assign n323 = n120 & n30036 ;
  assign n324 = n208 & n213 ;
  assign n325 = n323 | n324 ;
  assign n326 = n75 & n154 ;
  assign n327 = n79 & n101 ;
  assign n328 = n326 | n327 ;
  assign n329 = n325 | n328 ;
  assign n330 = n322 | n329 ;
  assign n331 = n75 & n109 ;
  assign n332 = n136 & n30037 ;
  assign n333 = n331 | n332 ;
  assign n334 = n82 & n132 ;
  assign n335 = n75 & n192 ;
  assign n336 = n334 | n335 ;
  assign n337 = n94 & n261 ;
  assign n338 = n94 & n110 ;
  assign n339 = n337 | n338 ;
  assign n340 = n336 | n339 ;
  assign n341 = n333 | n340 ;
  assign n342 = n330 | n341 ;
  assign n343 = n317 | n342 ;
  assign n344 = n86 & n115 ;
  assign n345 = n132 & n154 ;
  assign n346 = n82 & n178 ;
  assign n347 = n345 | n346 ;
  assign n348 = n127 & n136 ;
  assign n349 = n105 & n125 ;
  assign n350 = n348 | n349 ;
  assign n351 = n347 | n350 ;
  assign n352 = n344 | n351 ;
  assign n353 = n101 & n192 ;
  assign n354 = n101 & n125 ;
  assign n355 = n101 & n127 ;
  assign n356 = n354 | n355 ;
  assign n357 = n353 | n356 ;
  assign n358 = n30036 & n192 ;
  assign n359 = n82 & n105 ;
  assign n360 = n120 & n178 ;
  assign n361 = n359 | n360 ;
  assign n362 = n358 | n361 ;
  assign n363 = n357 | n362 ;
  assign n364 = n352 | n363 ;
  assign n365 = n125 & n136 ;
  assign n366 = n115 & n175 ;
  assign n367 = n365 | n366 ;
  assign n368 = n180 & n208 ;
  assign n369 = n30036 & n169 ;
  assign n370 = n368 | n369 ;
  assign n371 = n86 & n110 ;
  assign n372 = n82 & n208 ;
  assign n373 = n371 | n372 ;
  assign n374 = n370 | n373 ;
  assign n375 = n367 | n374 ;
  assign n376 = n105 & n169 ;
  assign n377 = n96 & n180 ;
  assign n378 = n376 | n377 ;
  assign n379 = n89 & n169 ;
  assign n380 = n79 & n89 ;
  assign n381 = n379 | n380 ;
  assign n382 = n378 | n381 ;
  assign n383 = n99 & n178 ;
  assign n384 = n30030 & n254 ;
  assign n385 = n383 | n384 ;
  assign n386 = n382 | n385 ;
  assign n387 = n375 | n386 ;
  assign n388 = n364 | n387 ;
  assign n389 = n343 | n388 ;
  assign n390 = n308 | n389 ;
  assign n30039 = ~n390 ;
  assign n391 = n231 & n30039 ;
  assign n30040 = ~n72 ;
  assign n392 = n30040 & n391 ;
  assign n30041 = ~n391 ;
  assign n393 = n72 & n30041 ;
  assign n394 = n392 | n393 ;
  assign n395 = n109 & n208 ;
  assign n396 = n99 & n30036 ;
  assign n397 = n90 | n396 ;
  assign n398 = n395 | n397 ;
  assign n399 = n127 & n132 ;
  assign n400 = n99 & n129 ;
  assign n401 = n94 & n156 ;
  assign n402 = n400 | n401 ;
  assign n403 = n399 | n402 ;
  assign n404 = n398 | n403 ;
  assign n405 = n96 & n192 ;
  assign n406 = n176 | n405 ;
  assign n407 = n132 & n180 ;
  assign n408 = n244 | n407 ;
  assign n409 = n406 | n408 ;
  assign n410 = n129 & n154 ;
  assign n411 = n277 | n410 ;
  assign n412 = n115 & n154 ;
  assign n413 = n411 | n412 ;
  assign n414 = n409 | n413 ;
  assign n415 = n404 | n414 ;
  assign n416 = n94 & n123 ;
  assign n417 = n109 & n156 ;
  assign n418 = n79 & n136 ;
  assign n419 = n417 | n418 ;
  assign n420 = n416 | n419 ;
  assign n421 = n253 | n420 ;
  assign n422 = n82 & n96 ;
  assign n423 = n276 | n312 ;
  assign n424 = n422 | n423 ;
  assign n425 = n196 | n424 ;
  assign n426 = n421 | n425 ;
  assign n427 = n415 | n426 ;
  assign n428 = n94 & n115 ;
  assign n429 = n240 | n428 ;
  assign n430 = n120 & n136 ;
  assign n431 = n300 | n430 ;
  assign n432 = n120 & n208 ;
  assign n433 = n30036 & n154 ;
  assign n434 = n86 & n101 ;
  assign n435 = n433 | n434 ;
  assign n436 = n432 | n435 ;
  assign n437 = n431 | n436 ;
  assign n438 = n429 | n437 ;
  assign n439 = n96 & n213 ;
  assign n440 = n82 & n89 ;
  assign n441 = n129 & n180 ;
  assign n442 = n440 | n441 ;
  assign n443 = n439 | n442 ;
  assign n444 = n291 | n443 ;
  assign n445 = n136 & n213 ;
  assign n446 = n96 & n127 ;
  assign n447 = n445 | n446 ;
  assign n448 = n122 & n169 ;
  assign n449 = n151 | n448 ;
  assign n450 = n447 | n449 ;
  assign n451 = n94 & n178 ;
  assign n452 = n75 & n99 ;
  assign n453 = n154 & n261 ;
  assign n454 = n452 | n453 ;
  assign n455 = n451 | n454 ;
  assign n456 = n450 | n455 ;
  assign n457 = n444 | n456 ;
  assign n458 = n438 | n457 ;
  assign n459 = n427 | n458 ;
  assign n460 = n105 & n154 ;
  assign n461 = n89 & n180 ;
  assign n462 = n358 | n461 ;
  assign n463 = n460 | n462 ;
  assign n464 = n99 & n208 ;
  assign n465 = n301 | n464 ;
  assign n466 = n270 | n377 ;
  assign n467 = n465 | n466 ;
  assign n468 = n463 | n467 ;
  assign n469 = n30037 & n178 ;
  assign n470 = n82 & n115 ;
  assign n471 = n348 | n470 ;
  assign n472 = n469 | n471 ;
  assign n473 = n79 & n30036 ;
  assign n474 = n213 & n261 ;
  assign n475 = n473 | n474 ;
  assign n476 = n82 & n110 ;
  assign n477 = n99 & n110 ;
  assign n478 = n476 | n477 ;
  assign n479 = n180 & n261 ;
  assign n480 = n110 & n127 ;
  assign n481 = n479 | n480 ;
  assign n482 = n478 | n481 ;
  assign n483 = n475 | n482 ;
  assign n484 = n472 | n483 ;
  assign n485 = n468 | n484 ;
  assign n486 = n129 & n192 ;
  assign n487 = n129 & n30037 ;
  assign n488 = n486 | n487 ;
  assign n489 = n156 & n213 ;
  assign n490 = n283 | n489 ;
  assign n491 = n96 & n30037 ;
  assign n492 = n186 | n491 ;
  assign n493 = n490 | n492 ;
  assign n494 = n488 | n493 ;
  assign n495 = n30037 & n261 ;
  assign n496 = n353 | n495 ;
  assign n497 = n132 & n30037 ;
  assign n498 = n223 | n497 ;
  assign n499 = n496 | n498 ;
  assign n500 = n75 & n180 ;
  assign n501 = n109 & n30036 ;
  assign n502 = n162 | n501 ;
  assign n503 = n500 | n502 ;
  assign n504 = n499 | n503 ;
  assign n505 = n494 | n504 ;
  assign n506 = n99 & n156 ;
  assign n507 = n103 | n506 ;
  assign n508 = n101 & n169 ;
  assign n509 = n89 & n127 ;
  assign n510 = n508 | n509 ;
  assign n511 = n507 | n510 ;
  assign n512 = n192 & n261 ;
  assign n513 = n171 | n512 ;
  assign n514 = n138 | n513 ;
  assign n515 = n511 | n514 ;
  assign n516 = n75 & n175 ;
  assign n517 = n86 & n105 ;
  assign n518 = n516 | n517 ;
  assign n519 = n124 | n518 ;
  assign n520 = n125 & n30036 ;
  assign n521 = n365 | n520 ;
  assign n522 = n326 | n371 ;
  assign n523 = n521 | n522 ;
  assign n524 = n519 | n523 ;
  assign n525 = n515 | n524 ;
  assign n526 = n505 | n525 ;
  assign n527 = n485 | n526 ;
  assign n528 = n105 & n109 ;
  assign n529 = n89 & n192 ;
  assign n530 = n528 | n529 ;
  assign n531 = n255 | n530 ;
  assign n532 = n89 & n213 ;
  assign n533 = n369 | n532 ;
  assign n534 = n96 & n120 ;
  assign n535 = n248 | n534 ;
  assign n536 = n533 | n535 ;
  assign n537 = n531 | n536 ;
  assign n538 = n109 & n261 ;
  assign n539 = n116 | n538 ;
  assign n540 = n125 & n156 ;
  assign n541 = n359 | n540 ;
  assign n542 = n156 & n180 ;
  assign n543 = n120 & n261 ;
  assign n544 = n542 | n543 ;
  assign n545 = n541 | n544 ;
  assign n546 = n539 | n545 ;
  assign n547 = n537 | n546 ;
  assign n548 = n99 & n132 ;
  assign n549 = n217 | n548 ;
  assign n550 = n120 & n132 ;
  assign n551 = n366 | n550 ;
  assign n552 = n549 | n551 ;
  assign n553 = n115 & n120 ;
  assign n554 = n101 & n180 ;
  assign n555 = n553 | n554 ;
  assign n556 = n313 | n555 ;
  assign n557 = n552 | n556 ;
  assign n558 = n547 | n557 ;
  assign n559 = n112 | n133 ;
  assign n560 = n156 & n192 ;
  assign n561 = n331 | n560 ;
  assign n562 = n559 | n561 ;
  assign n563 = n347 | n562 ;
  assign n564 = n110 & n192 ;
  assign n565 = n150 | n564 ;
  assign n566 = n139 | n384 ;
  assign n567 = n565 | n566 ;
  assign n568 = n82 & n261 ;
  assign n569 = n319 | n568 ;
  assign n570 = n293 | n338 ;
  assign n571 = n569 | n570 ;
  assign n572 = n187 | n318 ;
  assign n573 = n129 & n175 ;
  assign n574 = n269 | n573 ;
  assign n575 = n572 | n574 ;
  assign n576 = n571 | n575 ;
  assign n577 = n567 | n576 ;
  assign n578 = n563 | n577 ;
  assign n579 = n558 | n578 ;
  assign n580 = n527 | n579 ;
  assign n581 = n459 | n580 ;
  assign n582 = n394 & n581 ;
  assign n583 = n394 | n581 ;
  assign n30042 = ~n582 ;
  assign n584 = n30042 & n583 ;
  assign n585 = n337 | n379 ;
  assign n586 = n528 | n534 ;
  assign n587 = n245 | n480 ;
  assign n588 = n586 | n587 ;
  assign n589 = n585 | n588 ;
  assign n590 = n277 | n319 ;
  assign n591 = n75 & n213 ;
  assign n592 = n500 | n591 ;
  assign n593 = n590 | n592 ;
  assign n594 = x23 & n194 ;
  assign n595 = n217 | n594 ;
  assign n596 = n331 | n334 ;
  assign n597 = n432 | n596 ;
  assign n598 = n595 | n597 ;
  assign n599 = n593 | n598 ;
  assign n600 = n589 | n599 ;
  assign n601 = n185 | n520 ;
  assign n602 = n179 | n491 ;
  assign n603 = n318 | n407 ;
  assign n604 = n434 | n506 ;
  assign n605 = n603 | n604 ;
  assign n606 = n602 | n605 ;
  assign n607 = n601 | n606 ;
  assign n608 = n82 & n136 ;
  assign n609 = n538 | n608 ;
  assign n610 = n89 & n94 ;
  assign n611 = n212 | n610 ;
  assign n612 = n609 | n611 ;
  assign n613 = n187 | n258 ;
  assign n614 = n376 | n508 ;
  assign n615 = n613 | n614 ;
  assign n616 = n612 | n615 ;
  assign n617 = n433 | n501 ;
  assign n618 = n488 | n617 ;
  assign n619 = n291 | n618 ;
  assign n620 = n255 | n292 ;
  assign n621 = n123 & n192 ;
  assign n622 = n178 & n213 ;
  assign n623 = n621 | n622 ;
  assign n624 = n620 | n623 ;
  assign n625 = n619 | n624 ;
  assign n626 = n616 | n625 ;
  assign n627 = n607 | n626 ;
  assign n628 = n600 | n627 ;
  assign n30043 = ~n195 ;
  assign n629 = n145 & n30043 ;
  assign n630 = n136 & n154 ;
  assign n631 = n517 | n543 ;
  assign n632 = n630 | n631 ;
  assign n30044 = ~n632 ;
  assign n633 = n629 & n30044 ;
  assign n634 = n369 | n460 ;
  assign n635 = n94 & n208 ;
  assign n636 = n132 & n169 ;
  assign n637 = n635 | n636 ;
  assign n638 = n417 | n441 ;
  assign n639 = n637 | n638 ;
  assign n640 = n634 | n639 ;
  assign n641 = n271 | n293 ;
  assign n642 = n83 | n296 ;
  assign n643 = n344 | n642 ;
  assign n644 = n641 | n643 ;
  assign n645 = n640 | n644 ;
  assign n30045 = ~n645 ;
  assign n646 = n633 & n30045 ;
  assign n647 = n175 & n208 ;
  assign n648 = n232 | n348 ;
  assign n649 = n647 | n648 ;
  assign n650 = n263 | n400 ;
  assign n651 = n101 & n154 ;
  assign n652 = n560 | n651 ;
  assign n653 = n650 | n652 ;
  assign n654 = n235 | n474 ;
  assign n655 = n285 | n654 ;
  assign n656 = n653 | n655 ;
  assign n657 = n649 | n656 ;
  assign n658 = n110 & n30037 ;
  assign n659 = n312 | n658 ;
  assign n660 = n94 & n136 ;
  assign n661 = n368 | n660 ;
  assign n662 = n214 | n554 ;
  assign n663 = n661 | n662 ;
  assign n664 = n659 | n663 ;
  assign n665 = n223 | n469 ;
  assign n666 = n115 & n213 ;
  assign n667 = n665 | n666 ;
  assign n668 = n105 & n192 ;
  assign n669 = n461 | n668 ;
  assign n670 = n126 | n440 ;
  assign n671 = n669 | n670 ;
  assign n672 = n667 | n671 ;
  assign n673 = n664 | n672 ;
  assign n674 = n657 | n673 ;
  assign n30046 = ~n674 ;
  assign n675 = n646 & n30046 ;
  assign n676 = n94 & n129 ;
  assign n677 = n115 & n169 ;
  assign n678 = n676 | n677 ;
  assign n679 = n86 & n30036 ;
  assign n680 = n244 | n679 ;
  assign n681 = n678 | n680 ;
  assign n682 = n75 & n120 ;
  assign n683 = n405 | n682 ;
  assign n684 = n110 & n169 ;
  assign n685 = n199 | n684 ;
  assign n686 = n683 | n685 ;
  assign n687 = n79 & n178 ;
  assign n688 = n479 | n687 ;
  assign n689 = n372 | n422 ;
  assign n690 = n396 | n464 ;
  assign n691 = n689 | n690 ;
  assign n692 = n688 | n691 ;
  assign n693 = n686 | n692 ;
  assign n694 = n681 | n693 ;
  assign n695 = n127 & n208 ;
  assign n696 = n371 | n695 ;
  assign n697 = n310 | n696 ;
  assign n698 = n123 & n175 ;
  assign n699 = n395 | n698 ;
  assign n700 = n107 | n380 ;
  assign n701 = n239 | n700 ;
  assign n702 = n699 | n701 ;
  assign n703 = n697 | n702 ;
  assign n704 = n86 & n129 ;
  assign n705 = n216 | n512 ;
  assign n706 = n704 | n705 ;
  assign n707 = n327 | n353 ;
  assign n708 = n97 | n453 ;
  assign n709 = n707 | n708 ;
  assign n710 = n706 | n709 ;
  assign n711 = n123 & n180 ;
  assign n712 = n203 | n711 ;
  assign n713 = n109 & n178 ;
  assign n714 = n358 | n365 ;
  assign n715 = n713 | n714 ;
  assign n716 = n712 | n715 ;
  assign n717 = n710 | n716 ;
  assign n718 = n174 | n359 ;
  assign n719 = n412 | n718 ;
  assign n720 = n161 | n719 ;
  assign n721 = n30037 & n208 ;
  assign n722 = n123 & n125 ;
  assign n723 = n721 | n722 ;
  assign n724 = n385 | n723 ;
  assign n725 = n720 | n724 ;
  assign n726 = n717 | n725 ;
  assign n727 = n703 | n726 ;
  assign n728 = n694 | n727 ;
  assign n30047 = ~n728 ;
  assign n729 = n675 & n30047 ;
  assign n30048 = ~n628 ;
  assign n730 = n30048 & n729 ;
  assign n732 = n581 | n730 ;
  assign n733 = x0 | x1 ;
  assign n30049 = ~x2 ;
  assign n734 = n30049 & n733 ;
  assign n29884 = x2 & x3 ;
  assign n735 = x4 & n29884 ;
  assign n736 = x2 | x3 ;
  assign n30050 = ~n29884 ;
  assign n738 = n30050 & n736 ;
  assign n30051 = ~n736 ;
  assign n737 = x4 & n30051 ;
  assign n30052 = ~x4 ;
  assign n739 = n30052 & n29884 ;
  assign n740 = n737 | n739 ;
  assign n741 = n738 | n740 ;
  assign n30053 = ~x5 ;
  assign n742 = n30053 & n741 ;
  assign n743 = n735 | n742 ;
  assign n744 = n734 | n743 ;
  assign n745 = n734 & n743 ;
  assign n747 = n171 | n249 ;
  assign n748 = n489 | n528 ;
  assign n749 = n747 | n748 ;
  assign n750 = n30036 & n175 ;
  assign n751 = n217 | n750 ;
  assign n752 = n348 | n412 ;
  assign n753 = n751 | n752 ;
  assign n754 = n749 | n753 ;
  assign n755 = n433 | n713 ;
  assign n756 = n186 | n326 ;
  assign n757 = n722 | n756 ;
  assign n758 = n755 | n757 ;
  assign n759 = n344 | n487 ;
  assign n760 = n338 | n380 ;
  assign n761 = n676 | n760 ;
  assign n762 = n759 | n761 ;
  assign n763 = n758 | n762 ;
  assign n764 = n136 & n175 ;
  assign n765 = n110 & n213 ;
  assign n766 = n764 | n765 ;
  assign n767 = n79 & n261 ;
  assign n768 = n360 | n767 ;
  assign n769 = n766 | n768 ;
  assign n770 = n123 & n169 ;
  assign n771 = n682 | n770 ;
  assign n772 = n190 | n372 ;
  assign n773 = n658 | n772 ;
  assign n774 = n771 | n773 ;
  assign n775 = n769 | n774 ;
  assign n776 = n763 | n775 ;
  assign n777 = n754 | n776 ;
  assign n778 = n216 | n550 ;
  assign n779 = n347 | n778 ;
  assign n780 = n337 | n473 ;
  assign n781 = n491 | n704 ;
  assign n782 = n780 | n781 ;
  assign n783 = n779 | n782 ;
  assign n784 = n500 | n711 ;
  assign n785 = n195 | n273 ;
  assign n786 = n784 | n785 ;
  assign n787 = n783 | n786 ;
  assign n788 = n115 & n180 ;
  assign n789 = n301 | n379 ;
  assign n790 = n401 | n469 ;
  assign n791 = n789 | n790 ;
  assign n792 = n788 | n791 ;
  assign n793 = n110 & n125 ;
  assign n794 = n138 | n793 ;
  assign n795 = n30036 & n213 ;
  assign n796 = n283 | n795 ;
  assign n797 = n30030 & n297 ;
  assign n798 = n796 | n797 ;
  assign n799 = n794 | n798 ;
  assign n800 = n792 | n799 ;
  assign n801 = n787 | n800 ;
  assign n802 = n331 | n460 ;
  assign n803 = n508 | n802 ;
  assign n804 = n90 | n313 ;
  assign n805 = n199 | n804 ;
  assign n806 = n803 | n805 ;
  assign n807 = n272 | n668 ;
  assign n808 = n99 & n136 ;
  assign n809 = n553 | n808 ;
  assign n810 = n807 | n809 ;
  assign n811 = n96 & n154 ;
  assign n812 = n270 | n548 ;
  assign n813 = n811 | n812 ;
  assign n814 = n109 & n129 ;
  assign n815 = n543 | n814 ;
  assign n816 = n89 & n125 ;
  assign n817 = n815 | n816 ;
  assign n818 = n813 | n817 ;
  assign n819 = n810 | n818 ;
  assign n820 = n806 | n819 ;
  assign n821 = n801 | n820 ;
  assign n822 = n777 | n821 ;
  assign n823 = n174 | n532 ;
  assign n824 = n232 | n292 ;
  assign n825 = n823 | n824 ;
  assign n826 = n310 | n501 ;
  assign n827 = n101 & n175 ;
  assign n828 = n509 | n827 ;
  assign n829 = n826 | n828 ;
  assign n830 = n167 | n245 ;
  assign n831 = n104 | n830 ;
  assign n832 = n829 | n831 ;
  assign n833 = n123 & n30037 ;
  assign n834 = n396 | n833 ;
  assign n30054 = ~n416 ;
  assign n835 = n145 & n30054 ;
  assign n30055 = ~n834 ;
  assign n836 = n30055 & n835 ;
  assign n30056 = ~n832 ;
  assign n837 = n30056 & n836 ;
  assign n30057 = ~n825 ;
  assign n838 = n30057 & n837 ;
  assign n839 = n89 & n109 ;
  assign n840 = n223 | n839 ;
  assign n841 = n94 & n105 ;
  assign n842 = n452 | n841 ;
  assign n843 = n840 | n842 ;
  assign n844 = n130 | n477 ;
  assign n845 = n101 & n30037 ;
  assign n846 = n258 | n845 ;
  assign n847 = n844 | n846 ;
  assign n848 = n332 | n349 ;
  assign n849 = n358 | n534 ;
  assign n850 = n848 | n849 ;
  assign n851 = n847 | n850 ;
  assign n852 = n843 | n851 ;
  assign n853 = n395 | n666 ;
  assign n854 = n320 | n853 ;
  assign n855 = n355 | n486 ;
  assign n856 = n564 | n855 ;
  assign n857 = n101 & n213 ;
  assign n858 = n474 | n857 ;
  assign n859 = n133 | n176 ;
  assign n860 = n858 | n859 ;
  assign n861 = n856 | n860 ;
  assign n862 = n854 | n861 ;
  assign n863 = n852 | n862 ;
  assign n864 = n159 | n517 ;
  assign n865 = n30036 & n180 ;
  assign n866 = n695 | n865 ;
  assign n867 = n864 | n866 ;
  assign n868 = n323 | n461 ;
  assign n869 = n369 | n422 ;
  assign n870 = n253 | n335 ;
  assign n871 = n869 | n870 ;
  assign n872 = n868 | n871 ;
  assign n873 = n867 | n872 ;
  assign n874 = n376 | n542 ;
  assign n875 = n212 | n221 ;
  assign n876 = n445 | n875 ;
  assign n877 = n874 | n876 ;
  assign n878 = n429 | n877 ;
  assign n879 = n873 | n878 ;
  assign n880 = n863 | n879 ;
  assign n30058 = ~n880 ;
  assign n881 = n838 & n30058 ;
  assign n30059 = ~n822 ;
  assign n882 = n30059 & n881 ;
  assign n884 = n745 | n882 ;
  assign n885 = n744 & n884 ;
  assign n887 = n581 | n885 ;
  assign n886 = n581 & n885 ;
  assign n30060 = ~n886 ;
  assign n888 = n30060 & n887 ;
  assign n30061 = ~n29900 ;
  assign n108 = n30061 & n77 ;
  assign n889 = x31 & n108 ;
  assign n37284 = x26 & x27 ;
  assign n890 = x26 | x27 ;
  assign n30062 = ~n37284 ;
  assign n891 = n30062 & n890 ;
  assign n37285 = x28 & x29 ;
  assign n892 = x28 | x29 ;
  assign n30063 = ~n37285 ;
  assign n893 = n30063 & n892 ;
  assign n895 = n891 & n893 ;
  assign n896 = n220 | n369 ;
  assign n897 = n221 | n550 ;
  assign n898 = n807 | n897 ;
  assign n899 = n896 | n898 ;
  assign n900 = n99 & n123 ;
  assign n901 = n679 | n900 ;
  assign n30064 = ~n590 ;
  assign n902 = n145 & n30064 ;
  assign n30065 = ~n901 ;
  assign n903 = n30065 & n902 ;
  assign n904 = n366 | n432 ;
  assign n905 = n123 & n127 ;
  assign n906 = n174 | n905 ;
  assign n907 = n904 | n906 ;
  assign n30066 = ~n907 ;
  assign n908 = n903 & n30066 ;
  assign n30067 = ~n899 ;
  assign n909 = n30067 & n908 ;
  assign n910 = n407 | n695 ;
  assign n911 = n358 | n910 ;
  assign n912 = n318 | n540 ;
  assign n913 = n130 | n348 ;
  assign n914 = n912 | n913 ;
  assign n915 = n911 | n914 ;
  assign n916 = n292 | n666 ;
  assign n917 = n185 | n512 ;
  assign n918 = n916 | n917 ;
  assign n919 = n915 | n918 ;
  assign n920 = n296 | n359 ;
  assign n921 = n224 | n473 ;
  assign n922 = n480 | n921 ;
  assign n923 = n920 | n922 ;
  assign n924 = n176 | n827 ;
  assign n925 = n79 & n156 ;
  assign n926 = n721 | n925 ;
  assign n927 = n269 | n399 ;
  assign n928 = n926 | n927 ;
  assign n929 = n924 | n928 ;
  assign n30068 = ~n75 ;
  assign n144 = n30068 & n143 ;
  assign n30069 = ~n144 ;
  assign n930 = n94 & n30069 ;
  assign n193 = n79 | n192 ;
  assign n931 = n89 & n193 ;
  assign n932 = n930 | n931 ;
  assign n262 = n101 | n261 ;
  assign n933 = n99 & n262 ;
  assign n934 = n232 | n765 ;
  assign n935 = n933 | n934 ;
  assign n936 = n932 | n935 ;
  assign n937 = n929 | n936 ;
  assign n938 = n923 | n937 ;
  assign n939 = n919 | n938 ;
  assign n30070 = ~n939 ;
  assign n940 = n909 & n30070 ;
  assign n941 = n190 | n273 ;
  assign n942 = n447 | n941 ;
  assign n943 = n510 | n942 ;
  assign n944 = n398 | n678 ;
  assign n945 = n943 | n944 ;
  assign n946 = n489 | n568 ;
  assign n947 = n711 | n793 ;
  assign n948 = n946 | n947 ;
  assign n949 = n298 | n520 ;
  assign n950 = n245 | n270 ;
  assign n951 = n949 | n950 ;
  assign n952 = n948 | n951 ;
  assign n953 = n945 | n952 ;
  assign n954 = n400 | n622 ;
  assign n955 = n233 | n954 ;
  assign n956 = n660 | n865 ;
  assign n957 = n495 | n497 ;
  assign n958 = n487 | n957 ;
  assign n959 = n956 | n958 ;
  assign n960 = n955 | n959 ;
  assign n961 = n132 & n192 ;
  assign n962 = n255 | n961 ;
  assign n963 = n126 | n517 ;
  assign n964 = n554 | n560 ;
  assign n965 = n963 | n964 ;
  assign n966 = n428 | n683 ;
  assign n967 = n965 | n966 ;
  assign n968 = n962 | n967 ;
  assign n969 = n960 | n968 ;
  assign n970 = n953 | n969 ;
  assign n971 = n167 | n289 ;
  assign n972 = n469 | n704 ;
  assign n973 = n97 | n845 ;
  assign n974 = n972 | n973 ;
  assign n975 = n971 | n974 ;
  assign n976 = n365 | n553 ;
  assign n977 = n181 | n532 ;
  assign n978 = n169 & n261 ;
  assign n979 = n635 | n978 ;
  assign n980 = n977 | n979 ;
  assign n981 = n976 | n980 ;
  assign n982 = n416 | n713 ;
  assign n983 = n199 | n422 ;
  assign n984 = n982 | n983 ;
  assign n985 = n981 | n984 ;
  assign n986 = n975 | n985 ;
  assign n987 = n163 | n324 ;
  assign n988 = n338 | n987 ;
  assign n989 = n109 & n123 ;
  assign n990 = n636 | n989 ;
  assign n991 = n379 | n687 ;
  assign n992 = n276 | n461 ;
  assign n993 = n991 | n992 ;
  assign n994 = n990 | n993 ;
  assign n995 = n988 | n994 ;
  assign n996 = n96 & n109 ;
  assign n997 = n310 | n474 ;
  assign n998 = n996 | n997 ;
  assign n999 = n249 | n608 ;
  assign n1000 = n647 | n999 ;
  assign n1001 = n998 | n1000 ;
  assign n1002 = n542 | n767 ;
  assign n1003 = n171 | n327 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = n80 | n372 ;
  assign n1006 = n814 | n1005 ;
  assign n1007 = n1004 | n1006 ;
  assign n1008 = n1001 | n1007 ;
  assign n1009 = n150 | n384 ;
  assign n1010 = n132 & n175 ;
  assign n1011 = n323 | n1010 ;
  assign n1012 = n368 | n410 ;
  assign n1013 = n1011 | n1012 ;
  assign n1014 = n1009 | n1013 ;
  assign n1015 = n212 | n240 ;
  assign n1016 = n478 | n1015 ;
  assign n1017 = n549 | n1016 ;
  assign n1018 = n1014 | n1017 ;
  assign n1019 = n1008 | n1018 ;
  assign n1020 = n995 | n1019 ;
  assign n1021 = n986 | n1020 ;
  assign n1022 = n970 | n1021 ;
  assign n30071 = ~n1022 ;
  assign n1023 = n940 & n30071 ;
  assign n1025 = n130 | n433 ;
  assign n1026 = n460 | n528 ;
  assign n1027 = n1025 | n1026 ;
  assign n1028 = n179 | n241 ;
  assign n1029 = n302 | n540 ;
  assign n1030 = n1028 | n1029 ;
  assign n1031 = n1027 | n1030 ;
  assign n1032 = n263 | n594 ;
  assign n1033 = n203 | n651 ;
  assign n1034 = n470 | n1033 ;
  assign n1035 = n440 | n610 ;
  assign n1036 = n407 | n795 ;
  assign n1037 = n1035 | n1036 ;
  assign n1038 = n1034 | n1037 ;
  assign n1039 = n1032 | n1038 ;
  assign n1040 = n1031 | n1039 ;
  assign n1041 = n186 | n833 ;
  assign n1042 = n464 | n486 ;
  assign n1043 = n1041 | n1042 ;
  assign n1044 = n500 | n765 ;
  assign n1045 = n141 | n807 ;
  assign n1046 = n1044 | n1045 ;
  assign n1047 = n123 & n213 ;
  assign n1048 = n930 | n1047 ;
  assign n1049 = n30037 & n156 ;
  assign n1050 = n235 | n1049 ;
  assign n1051 = n202 | n430 ;
  assign n1052 = n1050 | n1051 ;
  assign n1053 = n1048 | n1052 ;
  assign n1054 = n1046 | n1053 ;
  assign n1055 = n1043 | n1054 ;
  assign n1056 = n258 | n280 ;
  assign n1057 = n441 | n1056 ;
  assign n1058 = n158 | n529 ;
  assign n1059 = n151 | n401 ;
  assign n1060 = n550 | n1059 ;
  assign n1061 = n1058 | n1060 ;
  assign n1062 = n1057 | n1061 ;
  assign n1063 = n279 | n538 ;
  assign n1064 = n921 | n1063 ;
  assign n1065 = n901 | n1064 ;
  assign n1066 = n797 | n925 ;
  assign n1067 = n721 | n770 ;
  assign n1068 = n1066 | n1067 ;
  assign n1069 = n1065 | n1068 ;
  assign n1070 = n1062 | n1069 ;
  assign n1071 = n1055 | n1070 ;
  assign n1072 = n1040 | n1071 ;
  assign n1073 = n389 | n970 ;
  assign n1074 = n1072 | n1073 ;
  assign n1077 = n1023 & n1074 ;
  assign n1081 = n1023 | n1074 ;
  assign n30072 = ~n1077 ;
  assign n1082 = n30072 & n1081 ;
  assign n1083 = n418 | n486 ;
  assign n1084 = n811 | n1083 ;
  assign n1085 = n168 | n293 ;
  assign n1086 = n300 | n319 ;
  assign n1087 = n1085 | n1086 ;
  assign n1088 = n683 | n1087 ;
  assign n1089 = n1084 | n1088 ;
  assign n1090 = n556 | n1089 ;
  assign n1091 = n101 & n109 ;
  assign n1092 = n150 | n1091 ;
  assign n1093 = n241 | n497 ;
  assign n1094 = n564 | n1093 ;
  assign n1095 = n432 | n489 ;
  assign n1096 = n239 | n1095 ;
  assign n1097 = n1094 | n1096 ;
  assign n1098 = n1092 | n1097 ;
  assign n1099 = n115 & n192 ;
  assign n1100 = n501 | n1099 ;
  assign n1101 = n433 | n684 ;
  assign n1102 = n359 | n1101 ;
  assign n1103 = n1100 | n1102 ;
  assign n1104 = n97 | n608 ;
  assign n1105 = n126 | n1104 ;
  assign n1106 = n290 | n349 ;
  assign n1107 = n1105 | n1106 ;
  assign n1108 = n1103 | n1107 ;
  assign n1109 = n212 | n380 ;
  assign n1110 = n445 | n476 ;
  assign n1111 = n377 | n422 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n1109 | n1112 ;
  assign n1114 = n399 | n534 ;
  assign n1115 = n139 | n280 ;
  assign n1116 = n371 | n464 ;
  assign n1117 = n1115 | n1116 ;
  assign n1118 = n1114 | n1117 ;
  assign n1119 = n1113 | n1118 ;
  assign n1120 = n1108 | n1119 ;
  assign n1121 = n1098 | n1120 ;
  assign n1122 = n1090 | n1121 ;
  assign n1123 = n383 | n1047 ;
  assign n1124 = n358 | n376 ;
  assign n1125 = n610 | n1124 ;
  assign n1126 = n337 | n621 ;
  assign n1127 = n1125 | n1126 ;
  assign n1128 = n1123 | n1127 ;
  assign n1129 = n82 & n123 ;
  assign n1130 = n298 | n344 ;
  assign n1131 = n1129 | n1130 ;
  assign n1132 = n591 | n721 ;
  assign n1133 = n491 | n1049 ;
  assign n1134 = n1132 | n1133 ;
  assign n1135 = n309 | n538 ;
  assign n1136 = n658 | n795 ;
  assign n1137 = n1135 | n1136 ;
  assign n1138 = n1134 | n1137 ;
  assign n1139 = n1131 | n1138 ;
  assign n1140 = n1128 | n1139 ;
  assign n1141 = n195 | n630 ;
  assign n1142 = n216 | n312 ;
  assign n1143 = n687 | n978 ;
  assign n1144 = n1142 | n1143 ;
  assign n1145 = n1141 | n1144 ;
  assign n1146 = n171 | n257 ;
  assign n1147 = n348 | n827 ;
  assign n1148 = n560 | n1147 ;
  assign n1149 = n1146 | n1148 ;
  assign n1150 = n825 | n1149 ;
  assign n1151 = n1145 | n1150 ;
  assign n111 = n105 | n110 ;
  assign n1152 = n94 & n111 ;
  assign n1153 = n202 | n326 ;
  assign n1154 = n1152 | n1153 ;
  assign n1155 = n157 | n379 ;
  assign n1156 = n417 | n517 ;
  assign n1157 = n1155 | n1156 ;
  assign n1158 = n955 | n1157 ;
  assign n1159 = n1154 | n1158 ;
  assign n1160 = n335 | n446 ;
  assign n1161 = n430 | n865 ;
  assign n1162 = n244 | n410 ;
  assign n1163 = n1161 | n1162 ;
  assign n1164 = n1160 | n1163 ;
  assign n1165 = n237 | n594 ;
  assign n1166 = n528 | n839 ;
  assign n1167 = n263 | n314 ;
  assign n1168 = n1166 | n1167 ;
  assign n1169 = n1165 | n1168 ;
  assign n1170 = n1164 | n1169 ;
  assign n1171 = n1159 | n1170 ;
  assign n1172 = n1151 | n1171 ;
  assign n1173 = n1140 | n1172 ;
  assign n1174 = n345 | n543 ;
  assign n1175 = n222 | n666 ;
  assign n1176 = n1174 | n1175 ;
  assign n1177 = n185 | n996 ;
  assign n1178 = n249 | n272 ;
  assign n1179 = n129 & n213 ;
  assign n1180 = n508 | n1179 ;
  assign n1181 = n1178 | n1180 ;
  assign n1182 = n1177 | n1181 ;
  assign n1183 = n660 | n833 ;
  assign n1184 = n441 | n573 ;
  assign n1185 = n788 | n1184 ;
  assign n1186 = n1183 | n1185 ;
  assign n1187 = n1182 | n1186 ;
  assign n1188 = n1176 | n1187 ;
  assign n1189 = n279 | n434 ;
  assign n1190 = n647 | n816 ;
  assign n1191 = n1189 | n1190 ;
  assign n1192 = n116 | n961 ;
  assign n1193 = n550 | n635 ;
  assign n1194 = n858 | n1193 ;
  assign n1195 = n1192 | n1194 ;
  assign n1196 = n1191 | n1195 ;
  assign n1197 = n372 | n679 ;
  assign n1198 = n713 | n1197 ;
  assign n1199 = n99 & n261 ;
  assign n1200 = n179 | n1199 ;
  assign n1201 = n186 | n273 ;
  assign n1202 = n1200 | n1201 ;
  assign n1203 = n1198 | n1202 ;
  assign n1204 = n256 | n922 ;
  assign n1205 = n1203 | n1204 ;
  assign n1206 = n520 | n764 ;
  assign n1207 = n613 | n1206 ;
  assign n1208 = n429 | n1207 ;
  assign n1209 = n310 | n334 ;
  assign n1210 = n103 | n223 ;
  assign n1211 = n190 | n323 ;
  assign n1212 = n1210 | n1211 ;
  assign n1213 = n1209 | n1212 ;
  assign n1214 = n1208 | n1213 ;
  assign n1215 = n1205 | n1214 ;
  assign n1216 = n1196 | n1215 ;
  assign n1217 = n1188 | n1216 ;
  assign n1218 = n1173 | n1217 ;
  assign n1219 = n1122 | n1218 ;
  assign n30073 = ~n1219 ;
  assign n1220 = n1023 & n30073 ;
  assign n30074 = ~n1023 ;
  assign n1225 = n30074 & n1219 ;
  assign n1226 = n1220 | n1225 ;
  assign n1227 = n163 | n622 ;
  assign n1228 = n1010 | n1227 ;
  assign n1229 = n795 | n1091 ;
  assign n1230 = n353 | n538 ;
  assign n1231 = n1229 | n1230 ;
  assign n1232 = n1228 | n1231 ;
  assign n1233 = n214 | n564 ;
  assign n1234 = n271 | n1233 ;
  assign n1235 = n367 | n1004 ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = n1232 | n1236 ;
  assign n1238 = n358 | n428 ;
  assign n1239 = n322 | n1066 ;
  assign n1240 = n1238 | n1239 ;
  assign n1241 = n241 | n276 ;
  assign n1242 = n433 | n816 ;
  assign n1243 = n501 | n764 ;
  assign n1244 = n1242 | n1243 ;
  assign n1245 = n1241 | n1244 ;
  assign n1246 = n240 | n434 ;
  assign n1247 = n1200 | n1246 ;
  assign n1248 = n159 | n331 ;
  assign n1249 = n181 | n407 ;
  assign n1250 = n1248 | n1249 ;
  assign n1251 = n1247 | n1250 ;
  assign n1252 = n96 & n169 ;
  assign n1253 = n290 | n1252 ;
  assign n1254 = n344 | n683 ;
  assign n1255 = n1253 | n1254 ;
  assign n1256 = n1251 | n1255 ;
  assign n1257 = n1245 | n1256 ;
  assign n1258 = n1240 | n1257 ;
  assign n1259 = n1237 | n1258 ;
  assign n1260 = n573 | n957 ;
  assign n1261 = n1259 | n1260 ;
  assign n30075 = ~n469 ;
  assign n1262 = n145 & n30075 ;
  assign n30076 = ~n811 ;
  assign n1263 = n30076 & n1262 ;
  assign n30077 = ~n255 ;
  assign n1264 = n30077 & n1263 ;
  assign n1265 = n225 | n314 ;
  assign n1266 = n510 | n1265 ;
  assign n1267 = n239 | n334 ;
  assign n1268 = n678 | n1267 ;
  assign n1269 = n1266 | n1268 ;
  assign n30078 = ~n1269 ;
  assign n1270 = n1264 & n30078 ;
  assign n1271 = n133 | n292 ;
  assign n1272 = n103 | n309 ;
  assign n1273 = n368 | n412 ;
  assign n1274 = n1272 | n1273 ;
  assign n1275 = n1271 | n1274 ;
  assign n1276 = n400 | n1129 ;
  assign n1277 = n263 | n289 ;
  assign n1278 = n608 | n1277 ;
  assign n1279 = n150 | n865 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = n1276 | n1280 ;
  assign n1282 = n460 | n478 ;
  assign n1283 = n722 | n1282 ;
  assign n1284 = n452 | n610 ;
  assign n1285 = n815 | n1284 ;
  assign n1286 = n788 | n793 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = n1283 | n1287 ;
  assign n1289 = n1281 | n1288 ;
  assign n1290 = n1275 | n1289 ;
  assign n30079 = ~n1290 ;
  assign n1291 = n1270 & n30079 ;
  assign n1292 = n900 | n1099 ;
  assign n1293 = n491 | n1179 ;
  assign n1294 = n360 | n516 ;
  assign n1295 = n1293 | n1294 ;
  assign n1296 = n1292 | n1295 ;
  assign n1297 = n451 | n651 ;
  assign n1298 = n721 | n1297 ;
  assign n1300 = n245 | n369 ;
  assign n1301 = n698 | n1300 ;
  assign n1302 = n1298 | n1301 ;
  assign n1303 = n983 | n1302 ;
  assign n1304 = n1296 | n1303 ;
  assign n1305 = n258 | n470 ;
  assign n1306 = n279 | n395 ;
  assign n1307 = n1305 | n1306 ;
  assign n1308 = n205 | n695 ;
  assign n1309 = n83 | n839 ;
  assign n1310 = n833 | n1309 ;
  assign n1311 = n216 | n441 ;
  assign n1312 = n232 | n827 ;
  assign n1313 = n1311 | n1312 ;
  assign n1314 = n1310 | n1313 ;
  assign n1315 = n1308 | n1314 ;
  assign n1316 = n1307 | n1315 ;
  assign n1317 = n190 | n560 ;
  assign n1318 = n978 | n1317 ;
  assign n1319 = n116 | n1318 ;
  assign n1320 = n349 | n550 ;
  assign n1321 = n97 | n1049 ;
  assign n1322 = n1320 | n1321 ;
  assign n1323 = n277 | n548 ;
  assign n1324 = n512 | n750 ;
  assign n1325 = n1323 | n1324 ;
  assign n1326 = n1322 | n1325 ;
  assign n1327 = n253 | n345 ;
  assign n1328 = n500 | n1327 ;
  assign n1329 = n250 | n823 ;
  assign n1330 = n1328 | n1329 ;
  assign n1331 = n1326 | n1330 ;
  assign n1332 = n1319 | n1331 ;
  assign n1333 = n1316 | n1332 ;
  assign n1334 = n1304 | n1333 ;
  assign n30080 = ~n1334 ;
  assign n1335 = n1291 & n30080 ;
  assign n30081 = ~n1261 ;
  assign n1336 = n30081 & n1335 ;
  assign n1337 = n30073 & n1336 ;
  assign n30082 = ~n1336 ;
  assign n1342 = n1219 & n30082 ;
  assign n1343 = n1337 | n1342 ;
  assign n1344 = n422 | n500 ;
  assign n1345 = n554 | n1344 ;
  assign n1346 = n171 | n346 ;
  assign n284 = n236 | n283 ;
  assign n1347 = n376 | n516 ;
  assign n1348 = n284 | n1347 ;
  assign n1349 = n1346 | n1348 ;
  assign n1350 = n1345 | n1349 ;
  assign n1351 = n1275 | n1350 ;
  assign n1352 = n150 | n377 ;
  assign n1354 = n216 | n320 ;
  assign n1355 = n360 | n1354 ;
  assign n1356 = n232 | n240 ;
  assign n1357 = n1029 | n1356 ;
  assign n1358 = n1355 | n1357 ;
  assign n1359 = n1352 | n1358 ;
  assign n1360 = n138 | n290 ;
  assign n1361 = n116 | n399 ;
  assign n1362 = n167 | n651 ;
  assign n1363 = n925 | n1362 ;
  assign n1364 = n1361 | n1363 ;
  assign n1365 = n1360 | n1364 ;
  assign n209 = n115 | n208 ;
  assign n210 = n110 | n209 ;
  assign n1366 = n175 & n210 ;
  assign n1367 = n358 | n489 ;
  assign n1368 = n379 | n476 ;
  assign n1369 = n1367 | n1368 ;
  assign n1370 = n591 | n765 ;
  assign n1371 = n112 | n354 ;
  assign n1372 = n1370 | n1371 ;
  assign n1373 = n1369 | n1372 ;
  assign n1374 = n1366 | n1373 ;
  assign n1375 = n1365 | n1374 ;
  assign n1376 = n1359 | n1375 ;
  assign n1377 = n1351 | n1376 ;
  assign n1378 = n300 | n538 ;
  assign n1379 = n327 | n407 ;
  assign n1380 = n797 | n1379 ;
  assign n1381 = n1378 | n1380 ;
  assign n1382 = n532 | n698 ;
  assign n1383 = n809 | n1382 ;
  assign n1384 = n168 | n542 ;
  assign n1385 = n780 | n858 ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = n1383 | n1386 ;
  assign n1388 = n1381 | n1387 ;
  assign n1389 = n722 | n1047 ;
  assign n1390 = n205 | n430 ;
  assign n1391 = n848 | n1035 ;
  assign n1392 = n1390 | n1391 ;
  assign n1393 = n1389 | n1392 ;
  assign n1394 = n217 | n416 ;
  assign n1395 = n450 | n1394 ;
  assign n1396 = n641 | n1102 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = n1393 | n1397 ;
  assign n1399 = n1388 | n1398 ;
  assign n1400 = n1188 | n1399 ;
  assign n1401 = n402 | n634 ;
  assign n1402 = n905 | n989 ;
  assign n1403 = n1401 | n1402 ;
  assign n1404 = n509 | n795 ;
  assign n1405 = n793 | n1404 ;
  assign n1406 = n83 | n97 ;
  assign n1407 = n365 | n405 ;
  assign n1408 = n1406 | n1407 ;
  assign n1409 = n1405 | n1408 ;
  assign n1410 = n1403 | n1409 ;
  assign n1411 = n384 | n695 ;
  assign n1412 = n301 | n1411 ;
  assign n1413 = n312 | n961 ;
  assign n1414 = n668 | n764 ;
  assign n1415 = n282 | n372 ;
  assign n1416 = n1414 | n1415 ;
  assign n1417 = n1413 | n1416 ;
  assign n1418 = n1412 | n1417 ;
  assign n1419 = n1410 | n1418 ;
  assign n1420 = n497 | n870 ;
  assign n1421 = n635 | n687 ;
  assign n1422 = n158 | n608 ;
  assign n1423 = n200 | n464 ;
  assign n1424 = n1422 | n1423 ;
  assign n1425 = n1421 | n1424 ;
  assign n1426 = n1420 | n1425 ;
  assign n1427 = n139 | n841 ;
  assign n1428 = n978 | n1427 ;
  assign n1429 = n124 | n1129 ;
  assign n1430 = n477 | n548 ;
  assign n1431 = n434 | n512 ;
  assign n1432 = n1430 | n1431 ;
  assign n1433 = n1429 | n1432 ;
  assign n1434 = n1428 | n1433 ;
  assign n1435 = n80 | n244 ;
  assign n1436 = n214 | n1435 ;
  assign n1437 = n174 | n235 ;
  assign n1438 = n380 | n1437 ;
  assign n1439 = n1267 | n1438 ;
  assign n1440 = n1436 | n1439 ;
  assign n1441 = n1434 | n1440 ;
  assign n1442 = n1426 | n1441 ;
  assign n1443 = n1419 | n1442 ;
  assign n1444 = n1400 | n1443 ;
  assign n1445 = n1377 | n1444 ;
  assign n30083 = ~n1445 ;
  assign n1446 = n1336 & n30083 ;
  assign n1450 = n30082 & n1445 ;
  assign n1451 = n1446 | n1450 ;
  assign n1452 = n497 | n554 ;
  assign n1453 = n124 | n1452 ;
  assign n1454 = n133 | n337 ;
  assign n1455 = n439 | n1252 ;
  assign n1456 = n1454 | n1455 ;
  assign n1457 = n1453 | n1456 ;
  assign n1458 = n159 | n279 ;
  assign n1459 = n630 | n1458 ;
  assign n1460 = n1125 | n1459 ;
  assign n1461 = n1177 | n1460 ;
  assign n1462 = n1457 | n1461 ;
  assign n1463 = n441 | n470 ;
  assign n1464 = n174 | n293 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = n150 | n383 ;
  assign n1467 = n1389 | n1466 ;
  assign n1468 = n296 | n365 ;
  assign n1469 = n236 | n841 ;
  assign n1470 = n1468 | n1469 ;
  assign n1471 = n80 | n440 ;
  assign n1472 = n216 | n679 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = n1470 | n1473 ;
  assign n1475 = n1467 | n1474 ;
  assign n1476 = n1465 | n1475 ;
  assign n1477 = n239 | n961 ;
  assign n1478 = n171 | n647 ;
  assign n1479 = n1091 | n1478 ;
  assign n1480 = n900 | n1479 ;
  assign n1481 = n1477 | n1480 ;
  assign n1482 = n222 | n278 ;
  assign n1483 = n300 | n310 ;
  assign n1485 = n1166 | n1483 ;
  assign n1486 = n1482 | n1485 ;
  assign n1487 = n90 | n698 ;
  assign n1488 = n369 | n380 ;
  assign n1489 = n1049 | n1488 ;
  assign n1490 = n1487 | n1489 ;
  assign n1491 = n1486 | n1490 ;
  assign n1492 = n1481 | n1491 ;
  assign n1493 = n1476 | n1492 ;
  assign n1494 = n1462 | n1493 ;
  assign n1495 = n301 | n529 ;
  assign n1496 = n202 | n548 ;
  assign n1497 = n83 | n461 ;
  assign n1498 = n1496 | n1497 ;
  assign n1499 = n1495 | n1498 ;
  assign n1500 = n313 | n795 ;
  assign n1501 = n495 | n1500 ;
  assign n1502 = n217 | n793 ;
  assign n1503 = n978 | n1502 ;
  assign n1504 = n955 | n1503 ;
  assign n1505 = n1501 | n1504 ;
  assign n1506 = n1499 | n1505 ;
  assign n1507 = n1100 | n1234 ;
  assign n1508 = n158 | n335 ;
  assign n1509 = n621 | n1508 ;
  assign n1510 = n354 | n384 ;
  assign n1511 = n1509 | n1510 ;
  assign n1512 = n1507 | n1511 ;
  assign n1513 = n476 | n573 ;
  assign n1514 = n1162 | n1370 ;
  assign n1515 = n1513 | n1514 ;
  assign n1516 = n203 | n225 ;
  assign n1517 = n344 | n488 ;
  assign n1518 = n1516 | n1517 ;
  assign n1519 = n1515 | n1518 ;
  assign n1520 = n1512 | n1519 ;
  assign n1521 = n1506 | n1520 ;
  assign n1522 = n319 | n452 ;
  assign n1523 = n532 | n687 ;
  assign n1524 = n1522 | n1523 ;
  assign n1525 = n292 | n1524 ;
  assign n1526 = n157 | n273 ;
  assign n1527 = n473 | n1526 ;
  assign n1528 = n283 | n418 ;
  assign n1529 = n989 | n1528 ;
  assign n1530 = n1527 | n1529 ;
  assign n1531 = n253 | n635 ;
  assign n1532 = n348 | n543 ;
  assign n1533 = n104 | n1532 ;
  assign n1534 = n1531 | n1533 ;
  assign n1535 = n1530 | n1534 ;
  assign n1536 = n1525 | n1535 ;
  assign n1537 = n320 | n407 ;
  assign n1538 = n200 | n272 ;
  assign n1539 = n1011 | n1538 ;
  assign n1540 = n1537 | n1539 ;
  assign n1541 = n258 | n770 ;
  assign n1542 = n116 | n682 ;
  assign n1543 = n1541 | n1542 ;
  assign n1544 = n1540 | n1543 ;
  assign n1545 = n249 | n451 ;
  assign n1546 = n695 | n1545 ;
  assign n1547 = n797 | n1129 ;
  assign n1548 = n186 | n658 ;
  assign n1549 = n30031 & n175 ;
  assign n1550 = n1548 | n1549 ;
  assign n1551 = n1547 | n1550 ;
  assign n1552 = n1546 | n1551 ;
  assign n1553 = n1544 | n1552 ;
  assign n1554 = n1536 | n1553 ;
  assign n1555 = n1521 | n1554 ;
  assign n1556 = n1494 | n1555 ;
  assign n1562 = n1445 | n1556 ;
  assign n1559 = n30083 & n1556 ;
  assign n30084 = ~n1556 ;
  assign n1563 = n1445 & n30084 ;
  assign n1564 = n1559 | n1563 ;
  assign n1565 = n181 | n445 ;
  assign n1566 = n978 | n1565 ;
  assign n1567 = n151 | n622 ;
  assign n1568 = n695 | n925 ;
  assign n1569 = n1567 | n1568 ;
  assign n1570 = n1438 | n1569 ;
  assign n1571 = n1566 | n1570 ;
  assign n1572 = n253 | n722 ;
  assign n1573 = n433 | n1572 ;
  assign n1574 = n460 | n750 ;
  assign n1575 = n334 | n865 ;
  assign n1576 = n661 | n1575 ;
  assign n1577 = n1574 | n1576 ;
  assign n1578 = n1573 | n1577 ;
  assign n1579 = n1571 | n1578 ;
  assign n1580 = n905 | n971 ;
  assign n1581 = n1147 | n1580 ;
  assign n1582 = n440 | n486 ;
  assign n1583 = n1179 | n1582 ;
  assign n1584 = n162 | n432 ;
  assign n1585 = n540 | n1584 ;
  assign n1586 = n1583 | n1585 ;
  assign n1587 = n1581 | n1586 ;
  assign n30085 = ~n244 ;
  assign n1588 = n145 & n30085 ;
  assign n30086 = ~n338 ;
  assign n1589 = n30086 & n1588 ;
  assign n30087 = ~n593 ;
  assign n1590 = n30087 & n1589 ;
  assign n1591 = n354 | n658 ;
  assign n1592 = n439 | n1591 ;
  assign n1593 = n215 | n704 ;
  assign n1594 = n1592 | n1593 ;
  assign n30088 = ~n1594 ;
  assign n1595 = n1590 & n30088 ;
  assign n1596 = n249 | n479 ;
  assign n1597 = n241 | n314 ;
  assign n1598 = n453 | n1597 ;
  assign n1599 = n1596 | n1598 ;
  assign n1600 = n135 | n1599 ;
  assign n30089 = ~n1600 ;
  assign n1601 = n1595 & n30089 ;
  assign n30090 = ~n1587 ;
  assign n1602 = n30090 & n1601 ;
  assign n30091 = ~n1579 ;
  assign n1603 = n30091 & n1602 ;
  assign n1604 = n159 | n176 ;
  assign n1605 = n300 | n1604 ;
  assign n1606 = n548 | n845 ;
  assign n1607 = n1347 | n1606 ;
  assign n1608 = n1605 | n1607 ;
  assign n1609 = n185 | n594 ;
  assign n1610 = n1041 | n1106 ;
  assign n1611 = n1609 | n1610 ;
  assign n1612 = n1608 | n1611 ;
  assign n30092 = ~n1612 ;
  assign n1613 = n1603 & n30092 ;
  assign n1614 = n517 | n528 ;
  assign n1615 = n713 | n811 ;
  assign n1616 = n1614 | n1615 ;
  assign n1617 = n785 | n1616 ;
  assign n1618 = n360 | n677 ;
  assign n1619 = n171 | n245 ;
  assign n1620 = n1538 | n1619 ;
  assign n1621 = n1618 | n1620 ;
  assign n1622 = n1617 | n1621 ;
  assign n1623 = n203 | n365 ;
  assign n1624 = n535 | n1623 ;
  assign n1625 = n224 | n538 ;
  assign n1626 = n276 | n1049 ;
  assign n1627 = n1625 | n1626 ;
  assign n1628 = n1624 | n1627 ;
  assign n1629 = n1307 | n1628 ;
  assign n1630 = n107 | n297 ;
  assign n1631 = n335 | n480 ;
  assign n1632 = n1252 | n1631 ;
  assign n1633 = n1630 | n1632 ;
  assign n1634 = n179 | n711 ;
  assign n1635 = n355 | n808 ;
  assign n1636 = n532 | n1635 ;
  assign n1637 = n1634 | n1636 ;
  assign n1638 = n1633 | n1637 ;
  assign n1639 = n1629 | n1638 ;
  assign n1640 = n1622 | n1639 ;
  assign n1641 = n384 | n1099 ;
  assign n1642 = n858 | n1641 ;
  assign n1643 = n233 | n651 ;
  assign n1644 = n451 | n469 ;
  assign n1645 = n529 | n765 ;
  assign n1646 = n1644 | n1645 ;
  assign n1647 = n1643 | n1646 ;
  assign n1648 = n325 | n621 ;
  assign n1649 = n897 | n1648 ;
  assign n1650 = n1647 | n1649 ;
  assign n1651 = n1642 | n1650 ;
  assign n1652 = n495 | n608 ;
  assign n1653 = n610 | n1652 ;
  assign n1654 = n157 | n506 ;
  assign n1655 = n509 | n1654 ;
  assign n1656 = n1185 | n1655 ;
  assign n1657 = n1653 | n1656 ;
  assign n1658 = n477 | n512 ;
  assign n1659 = n636 | n767 ;
  assign n1660 = n1658 | n1659 ;
  assign n1661 = n916 | n1660 ;
  assign n1662 = n564 | n961 ;
  assign n1663 = n446 | n1199 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n400 | n900 ;
  assign n1666 = n1664 | n1665 ;
  assign n1667 = n1661 | n1666 ;
  assign n1668 = n1657 | n1667 ;
  assign n1669 = n1651 | n1668 ;
  assign n1670 = n1640 | n1669 ;
  assign n30093 = ~n1670 ;
  assign n1671 = n1613 & n30093 ;
  assign n1676 = n30084 & n1671 ;
  assign n1675 = n1556 & n1671 ;
  assign n1677 = n1556 | n1671 ;
  assign n30094 = ~n1675 ;
  assign n1678 = n30094 & n1677 ;
  assign n1679 = n418 | n573 ;
  assign n1680 = n628 | n1679 ;
  assign n1681 = n257 | n833 ;
  assign n1682 = n857 | n1681 ;
  assign n1683 = n167 | n417 ;
  assign n1684 = n439 | n839 ;
  assign n1685 = n722 | n1684 ;
  assign n1686 = n1683 | n1685 ;
  assign n1687 = n684 | n816 ;
  assign n1688 = n220 | n542 ;
  assign n1689 = n181 | n327 ;
  assign n1690 = n1688 | n1689 ;
  assign n1691 = n1687 | n1690 ;
  assign n1692 = n1686 | n1691 ;
  assign n1693 = n1682 | n1692 ;
  assign n1694 = n323 | n451 ;
  assign n1695 = n285 | n1129 ;
  assign n1696 = n1694 | n1695 ;
  assign n1697 = n320 | n428 ;
  assign n1698 = n174 | n540 ;
  assign n1699 = n865 | n1698 ;
  assign n1700 = n1697 | n1699 ;
  assign n1701 = n1696 | n1700 ;
  assign n1702 = n139 | n473 ;
  assign n1703 = n1091 | n1702 ;
  assign n1704 = n203 | n309 ;
  assign n1705 = n335 | n1704 ;
  assign n30095 = ~n130 ;
  assign n1706 = n30095 & n145 ;
  assign n30096 = ~n1294 ;
  assign n1707 = n30096 & n1706 ;
  assign n30097 = ~n1705 ;
  assign n1708 = n30097 & n1707 ;
  assign n30098 = ~n1703 ;
  assign n1709 = n30098 & n1708 ;
  assign n30099 = ~n1701 ;
  assign n1710 = n30099 & n1709 ;
  assign n30100 = ~n1693 ;
  assign n1711 = n30100 & n1710 ;
  assign n1712 = n126 | n410 ;
  assign n1713 = n263 | n1712 ;
  assign n1714 = n461 | n711 ;
  assign n1715 = n1643 | n1714 ;
  assign n1716 = n1713 | n1715 ;
  assign n1717 = n163 | n395 ;
  assign n1718 = n269 | n314 ;
  assign n1719 = n430 | n1718 ;
  assign n1720 = n1717 | n1719 ;
  assign n1721 = n565 | n1066 ;
  assign n1722 = n1720 | n1721 ;
  assign n1723 = n1716 | n1722 ;
  assign n1724 = n133 | n190 ;
  assign n1725 = n412 | n1724 ;
  assign n1726 = n326 | n989 ;
  assign n1727 = n901 | n1726 ;
  assign n1728 = n1725 | n1727 ;
  assign n1729 = n448 | n548 ;
  assign n1730 = n244 | n280 ;
  assign n1731 = n168 | n396 ;
  assign n1732 = n1730 | n1731 ;
  assign n1733 = n1729 | n1732 ;
  assign n1734 = n171 | n766 ;
  assign n1735 = n1152 | n1423 ;
  assign n1736 = n1734 | n1735 ;
  assign n1737 = n1733 | n1736 ;
  assign n1738 = n440 | n767 ;
  assign n1739 = n1252 | n1738 ;
  assign n1740 = n794 | n957 ;
  assign n1741 = n1739 | n1740 ;
  assign n1742 = n369 | n446 ;
  assign n1743 = n814 | n1742 ;
  assign n1744 = n279 | n324 ;
  assign n1745 = n344 | n1744 ;
  assign n1746 = n1743 | n1745 ;
  assign n1747 = n1741 | n1746 ;
  assign n1748 = n1737 | n1747 ;
  assign n1749 = n1728 | n1748 ;
  assign n1750 = n1723 | n1749 ;
  assign n30101 = ~n1750 ;
  assign n1751 = n1711 & n30101 ;
  assign n30102 = ~n1680 ;
  assign n1752 = n30102 & n1751 ;
  assign n1753 = n1671 & n1752 ;
  assign n1756 = n1671 | n1752 ;
  assign n30103 = ~n1753 ;
  assign n1757 = n30103 & n1756 ;
  assign n1758 = n255 | n529 ;
  assign n1759 = n107 | n1758 ;
  assign n1760 = n272 | n1199 ;
  assign n1761 = n245 | n591 ;
  assign n1762 = n233 | n1761 ;
  assign n1763 = n1760 | n1762 ;
  assign n1764 = n310 | n487 ;
  assign n1765 = n410 | n441 ;
  assign n1766 = n346 | n434 ;
  assign n1767 = n1765 | n1766 ;
  assign n1768 = n1764 | n1767 ;
  assign n1769 = n1763 | n1768 ;
  assign n1770 = n1759 | n1769 ;
  assign n1771 = n171 | n509 ;
  assign n1772 = n517 | n1771 ;
  assign n1773 = n366 | n924 ;
  assign n1774 = n1772 | n1773 ;
  assign n1775 = n289 | n550 ;
  assign n1776 = n788 | n1775 ;
  assign n1777 = n1141 | n1776 ;
  assign n1778 = n1774 | n1777 ;
  assign n1779 = n1701 | n1778 ;
  assign n1780 = n1770 | n1779 ;
  assign n1781 = n269 | n318 ;
  assign n1782 = n516 | n1781 ;
  assign n1783 = n1592 | n1782 ;
  assign n1784 = n130 | n158 ;
  assign n1785 = n244 | n332 ;
  assign n1786 = n1784 | n1785 ;
  assign n1787 = n86 & n156 ;
  assign n1788 = n376 | n1787 ;
  assign n1789 = n770 | n1788 ;
  assign n1790 = n1786 | n1789 ;
  assign n1791 = n1783 | n1790 ;
  assign n1792 = n162 | n263 ;
  assign n1793 = n402 | n1792 ;
  assign n1794 = n1468 | n1793 ;
  assign n1795 = n207 | n1794 ;
  assign n1796 = n1791 | n1795 ;
  assign n1797 = n112 | n232 ;
  assign n1798 = n845 | n1797 ;
  assign n1799 = n900 | n1798 ;
  assign n1800 = n235 | n277 ;
  assign n1801 = n302 | n1800 ;
  assign n1802 = n1799 | n1801 ;
  assign n1803 = n326 | n721 ;
  assign n1804 = n470 | n1803 ;
  assign n1805 = n496 | n1160 ;
  assign n1806 = n1248 | n1805 ;
  assign n1807 = n1804 | n1806 ;
  assign n1808 = n995 | n1807 ;
  assign n1809 = n1802 | n1808 ;
  assign n1810 = n1796 | n1809 ;
  assign n1811 = n1780 | n1810 ;
  assign n1812 = n1122 | n1811 ;
  assign n30104 = ~n1812 ;
  assign n1813 = n1752 & n30104 ;
  assign n30105 = ~n1752 ;
  assign n1818 = n30105 & n1812 ;
  assign n1819 = n1813 | n1818 ;
  assign n1820 = n181 | n520 ;
  assign n1821 = n90 | n487 ;
  assign n1822 = n300 | n349 ;
  assign n1823 = n205 | n1822 ;
  assign n1824 = n1821 | n1823 ;
  assign n1825 = n354 | n410 ;
  assign n1826 = n1099 | n1825 ;
  assign n1827 = n434 | n529 ;
  assign n1828 = n548 | n1827 ;
  assign n1829 = n1826 | n1828 ;
  assign n1830 = n378 | n406 ;
  assign n1831 = n814 | n1422 ;
  assign n1832 = n1830 | n1831 ;
  assign n1833 = n1829 | n1832 ;
  assign n1834 = n1824 | n1833 ;
  assign n1835 = n272 | n314 ;
  assign n1836 = n480 | n1835 ;
  assign n1837 = n1682 | n1836 ;
  assign n1838 = n717 | n1837 ;
  assign n1839 = n1834 | n1838 ;
  assign n1840 = n1820 | n1839 ;
  assign n1841 = n190 | n416 ;
  assign n1842 = n224 | n446 ;
  assign n1843 = n573 | n1842 ;
  assign n1844 = n1066 | n1843 ;
  assign n1845 = n1841 | n1844 ;
  assign n1846 = n124 | n1787 ;
  assign n1847 = n912 | n1846 ;
  assign n1848 = n202 | n221 ;
  assign n1849 = n241 | n1848 ;
  assign n1850 = n1500 | n1849 ;
  assign n1851 = n1847 | n1850 ;
  assign n1852 = n1845 | n1851 ;
  assign n1853 = n816 | n905 ;
  assign n1854 = n1166 | n1252 ;
  assign n1855 = n1853 | n1854 ;
  assign n1856 = n200 | n961 ;
  assign n1857 = n476 | n495 ;
  assign n1858 = n1856 | n1857 ;
  assign n1859 = n516 | n811 ;
  assign n1860 = n163 | n280 ;
  assign n1861 = n1859 | n1860 ;
  assign n1862 = n1858 | n1861 ;
  assign n1863 = n217 | n309 ;
  assign n1864 = n489 | n1863 ;
  assign n1865 = n334 | n1199 ;
  assign n1866 = n770 | n1865 ;
  assign n1867 = n1864 | n1866 ;
  assign n1868 = n1862 | n1867 ;
  assign n1869 = n1855 | n1868 ;
  assign n1870 = n168 | n292 ;
  assign n1871 = n346 | n500 ;
  assign n1872 = n827 | n1871 ;
  assign n1873 = n112 | n355 ;
  assign n1874 = n151 | n301 ;
  assign n1875 = n1873 | n1874 ;
  assign n1876 = n1872 | n1875 ;
  assign n1877 = n1870 | n1876 ;
  assign n1878 = n253 | n1469 ;
  assign n1879 = n501 | n1129 ;
  assign n1880 = n366 | n1688 ;
  assign n1881 = n1879 | n1880 ;
  assign n1882 = n1878 | n1881 ;
  assign n1883 = n1877 | n1882 ;
  assign n1884 = n1869 | n1883 ;
  assign n1885 = n1852 | n1884 ;
  assign n30106 = ~n1885 ;
  assign n1886 = n675 & n30106 ;
  assign n30107 = ~n1840 ;
  assign n1887 = n30107 & n1886 ;
  assign n1888 = n30104 & n1887 ;
  assign n30108 = ~n1887 ;
  assign n1890 = n1812 & n30108 ;
  assign n1891 = n1888 | n1890 ;
  assign n1892 = n240 | n309 ;
  assign n1893 = n973 | n1892 ;
  assign n1894 = n263 | n405 ;
  assign n1895 = n324 | n676 ;
  assign n1896 = n1894 | n1895 ;
  assign n1897 = n1893 | n1896 ;
  assign n1898 = n827 | n833 ;
  assign n1899 = n1789 | n1898 ;
  assign n1900 = n179 | n368 ;
  assign n1901 = n704 | n1900 ;
  assign n1902 = n528 | n797 ;
  assign n1903 = n1901 | n1902 ;
  assign n1904 = n1899 | n1903 ;
  assign n1905 = n1897 | n1904 ;
  assign n1906 = n253 | n337 ;
  assign n1907 = n417 | n422 ;
  assign n1908 = n1906 | n1907 ;
  assign n211 = n156 | n208 ;
  assign n1909 = n125 & n211 ;
  assign n1910 = n513 | n1909 ;
  assign n1911 = n1908 | n1910 ;
  assign n1912 = n205 | n345 ;
  assign n1913 = n432 | n814 ;
  assign n1914 = n961 | n1913 ;
  assign n1915 = n1912 | n1914 ;
  assign n1916 = n1911 | n1915 ;
  assign n1917 = n236 | n506 ;
  assign n1918 = n839 | n1010 ;
  assign n1919 = n1047 | n1918 ;
  assign n1920 = n1917 | n1919 ;
  assign n30109 = ~n1920 ;
  assign n1921 = n147 & n30109 ;
  assign n1922 = n312 | n418 ;
  assign n1923 = n282 | n430 ;
  assign n1924 = n199 | n1923 ;
  assign n1925 = n1922 | n1924 ;
  assign n1926 = n497 | n1035 ;
  assign n1927 = n353 | n668 ;
  assign n1928 = n320 | n338 ;
  assign n1929 = n1927 | n1928 ;
  assign n1930 = n1926 | n1929 ;
  assign n1931 = n1925 | n1930 ;
  assign n30110 = ~n1931 ;
  assign n1932 = n1921 & n30110 ;
  assign n30111 = ~n1916 ;
  assign n1933 = n30111 & n1932 ;
  assign n30112 = ~n1905 ;
  assign n1934 = n30112 & n1933 ;
  assign n1935 = n186 | n379 ;
  assign n1936 = n660 | n1091 ;
  assign n1937 = n1935 | n1936 ;
  assign n1938 = n475 | n1101 ;
  assign n1939 = n1937 | n1938 ;
  assign n1940 = n151 | n711 ;
  assign n1941 = n1106 | n1940 ;
  assign n1942 = n1939 | n1941 ;
  assign n1943 = n399 | n1252 ;
  assign n1944 = n1574 | n1766 ;
  assign n1945 = n1943 | n1944 ;
  assign n1946 = n1599 | n1945 ;
  assign n1947 = n163 | n279 ;
  assign n1948 = n371 | n1947 ;
  assign n1949 = n257 | n1948 ;
  assign n1950 = n310 | n905 ;
  assign n1951 = n176 | n372 ;
  assign n1952 = n1950 | n1951 ;
  assign n1953 = n1949 | n1952 ;
  assign n1954 = n1946 | n1953 ;
  assign n1955 = n1942 | n1954 ;
  assign n1956 = n1521 | n1955 ;
  assign n30113 = ~n1956 ;
  assign n1957 = n1934 & n30113 ;
  assign n1964 = n1887 & n1957 ;
  assign n30114 = ~n1957 ;
  assign n1959 = n1887 & n30114 ;
  assign n1965 = n30108 & n1957 ;
  assign n1966 = n1959 | n1965 ;
  assign n1967 = n273 | n453 ;
  assign n1968 = n124 | n440 ;
  assign n1969 = n1967 | n1968 ;
  assign n1970 = n349 | n816 ;
  assign n1971 = n553 | n1688 ;
  assign n1972 = n1970 | n1971 ;
  assign n1973 = n249 | n318 ;
  assign n1975 = n396 | n1973 ;
  assign n1976 = n336 | n406 ;
  assign n1977 = n1975 | n1976 ;
  assign n1978 = n1972 | n1977 ;
  assign n1979 = n1969 | n1978 ;
  assign n1980 = n112 | n319 ;
  assign n1981 = n116 | n1980 ;
  assign n1982 = n272 | n548 ;
  assign n1983 = n587 | n1982 ;
  assign n1984 = n1981 | n1983 ;
  assign n1985 = n332 | n400 ;
  assign n1986 = n529 | n1179 ;
  assign n1987 = n1985 | n1986 ;
  assign n1988 = n1177 | n1987 ;
  assign n1989 = n1984 | n1988 ;
  assign n1990 = n159 | n383 ;
  assign n1991 = n839 | n1990 ;
  assign n1992 = n1126 | n1991 ;
  assign n1993 = n1902 | n1992 ;
  assign n1994 = n139 | n795 ;
  assign n1996 = n630 | n1994 ;
  assign n1997 = n962 | n1713 ;
  assign n1998 = n1996 | n1997 ;
  assign n1999 = n1993 | n1998 ;
  assign n2000 = n1989 | n1999 ;
  assign n2001 = n1979 | n2000 ;
  assign n2002 = n162 | n1940 ;
  assign n2003 = n300 | n355 ;
  assign n2004 = n678 | n2003 ;
  assign n2005 = n1465 | n2004 ;
  assign n2006 = n2002 | n2005 ;
  assign n2007 = n216 | n258 ;
  assign n2008 = n371 | n517 ;
  assign n2009 = n2007 | n2008 ;
  assign n2010 = n199 | n412 ;
  assign n2011 = n2009 | n2010 ;
  assign n2012 = n1360 | n2011 ;
  assign n2013 = n301 | n417 ;
  assign n2014 = n345 | n534 ;
  assign n2015 = n2013 | n2014 ;
  assign n2016 = n360 | n1010 ;
  assign n2017 = n244 | n814 ;
  assign n2018 = n2016 | n2017 ;
  assign n2019 = n2015 | n2018 ;
  assign n2020 = n496 | n1694 ;
  assign n2021 = n367 | n2020 ;
  assign n2022 = n2019 | n2021 ;
  assign n2023 = n2012 | n2022 ;
  assign n2024 = n2006 | n2023 ;
  assign n2025 = n447 | n905 ;
  assign n30115 = ~n824 ;
  assign n2026 = n30115 & n835 ;
  assign n30116 = ~n2025 ;
  assign n2027 = n30116 & n2026 ;
  assign n2028 = n479 | n1431 ;
  assign n2029 = n327 | n395 ;
  assign n2030 = n253 | n439 ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = n2028 | n2031 ;
  assign n2033 = n723 | n759 ;
  assign n2034 = n2032 | n2033 ;
  assign n30117 = ~n2034 ;
  assign n2035 = n2027 & n30117 ;
  assign n2036 = n507 | n1591 ;
  assign n2037 = n379 | n540 ;
  assign n2038 = n1928 | n2037 ;
  assign n2039 = n2036 | n2038 ;
  assign n2040 = n543 | n698 ;
  assign n2041 = n282 | n765 ;
  assign n2042 = n225 | n2041 ;
  assign n2043 = n2040 | n2042 ;
  assign n2044 = n2039 | n2043 ;
  assign n2045 = n568 | n1129 ;
  assign n2046 = n845 | n1049 ;
  assign n2047 = n163 | n179 ;
  assign n2048 = n2046 | n2047 ;
  assign n2049 = n2045 | n2048 ;
  assign n2050 = n90 | n212 ;
  assign n2051 = n133 | n857 ;
  assign n2052 = n167 | n331 ;
  assign n2053 = n2051 | n2052 ;
  assign n2054 = n2050 | n2053 ;
  assign n2055 = n1149 | n2054 ;
  assign n2056 = n2049 | n2055 ;
  assign n2057 = n2044 | n2056 ;
  assign n30118 = ~n2057 ;
  assign n2058 = n2035 & n30118 ;
  assign n30119 = ~n2024 ;
  assign n2059 = n30119 & n2058 ;
  assign n30120 = ~n2001 ;
  assign n2060 = n30120 & n2059 ;
  assign n2063 = n1957 & n2060 ;
  assign n2064 = n1957 | n2060 ;
  assign n30121 = ~n2063 ;
  assign n2065 = n30121 & n2064 ;
  assign n2066 = n157 | n487 ;
  assign n2067 = n540 | n2066 ;
  assign n2068 = n570 | n896 ;
  assign n2069 = n2067 | n2068 ;
  assign n2070 = n255 | n480 ;
  assign n2071 = n223 | n355 ;
  assign n2072 = n1967 | n2071 ;
  assign n2073 = n2070 | n2072 ;
  assign n2074 = n2069 | n2073 ;
  assign n2075 = n1113 | n1268 ;
  assign n2076 = n2074 | n2075 ;
  assign n2077 = n1802 | n2076 ;
  assign n2078 = n713 | n1825 ;
  assign n2079 = n1786 | n2078 ;
  assign n2080 = n807 | n924 ;
  assign n2081 = n946 | n2080 ;
  assign n2082 = n2079 | n2081 ;
  assign n2083 = n107 | n464 ;
  assign n2084 = n610 | n2083 ;
  assign n2085 = n199 | n298 ;
  assign n2086 = n2084 | n2085 ;
  assign n2087 = n430 | n507 ;
  assign n2088 = n688 | n2087 ;
  assign n2089 = n2086 | n2088 ;
  assign n2090 = n2082 | n2089 ;
  assign n246 = n168 | n245 ;
  assign n2091 = n359 | n1681 ;
  assign n2092 = n246 | n2091 ;
  assign n2093 = n794 | n1160 ;
  assign n2094 = n1483 | n1574 ;
  assign n2095 = n2093 | n2094 ;
  assign n2096 = n195 | n301 ;
  assign n2097 = n420 | n2096 ;
  assign n2098 = n2095 | n2097 ;
  assign n2099 = n2092 | n2098 ;
  assign n2100 = n2090 | n2099 ;
  assign n2101 = n2077 | n2100 ;
  assign n2102 = n1261 | n2101 ;
  assign n30122 = ~n2102 ;
  assign n2103 = n2060 & n30122 ;
  assign n30123 = ~n2060 ;
  assign n2108 = n30123 & n2102 ;
  assign n2109 = n2103 | n2108 ;
  assign n2110 = n395 | n441 ;
  assign n2111 = n80 | n845 ;
  assign n2112 = n2110 | n2111 ;
  assign n2113 = n162 | n405 ;
  assign n2114 = n103 | n190 ;
  assign n2115 = n2113 | n2114 ;
  assign n2116 = n2112 | n2115 ;
  assign n2117 = n255 | n300 ;
  assign n2118 = n723 | n2117 ;
  assign n2119 = n2116 | n2118 ;
  assign n2120 = n330 | n2119 ;
  assign n2121 = n768 | n815 ;
  assign n2122 = n263 | n827 ;
  assign n2123 = n682 | n1049 ;
  assign n2124 = n2122 | n2123 ;
  assign n2125 = n2121 | n2124 ;
  assign n2126 = n130 | n301 ;
  assign n2127 = n432 | n2126 ;
  assign n2128 = n124 | n344 ;
  assign n2129 = n2127 | n2128 ;
  assign n2130 = n2125 | n2129 ;
  assign n2131 = n187 | n217 ;
  assign n2132 = n839 | n2131 ;
  assign n2133 = n711 | n2132 ;
  assign n2134 = n311 | n418 ;
  assign n2135 = n788 | n2134 ;
  assign n2136 = n2133 | n2135 ;
  assign n2137 = n2130 | n2136 ;
  assign n2138 = n314 | n816 ;
  assign n2139 = n282 | n500 ;
  assign n2140 = n296 | n430 ;
  assign n2141 = n2139 | n2140 ;
  assign n2142 = n2138 | n2141 ;
  assign n2143 = n651 | n1452 ;
  assign n2144 = n649 | n2143 ;
  assign n2145 = n2142 | n2144 ;
  assign n2146 = n480 | n764 ;
  assign n2147 = n1091 | n2146 ;
  assign n2148 = n553 | n696 ;
  assign n2149 = n1664 | n2148 ;
  assign n2150 = n2147 | n2149 ;
  assign n2151 = n2145 | n2150 ;
  assign n2152 = n2137 | n2151 ;
  assign n2153 = n2120 | n2152 ;
  assign n2154 = n83 | n416 ;
  assign n2155 = n359 | n1454 ;
  assign n2156 = n2154 | n2155 ;
  assign n2157 = n660 | n930 ;
  assign n2158 = n470 | n1129 ;
  assign n2159 = n2157 | n2158 ;
  assign n2160 = n97 | n451 ;
  assign n2161 = n1422 | n2160 ;
  assign n2162 = n334 | n568 ;
  assign n2163 = n1152 | n2162 ;
  assign n2164 = n2161 | n2163 ;
  assign n2165 = n2159 | n2164 ;
  assign n2166 = n2156 | n2165 ;
  assign n2167 = n248 | n376 ;
  assign n2168 = n2166 | n2167 ;
  assign n2169 = n277 | n594 ;
  assign n2170 = n167 | n214 ;
  assign n2171 = n280 | n2170 ;
  assign n2172 = n204 | n2171 ;
  assign n2173 = n2169 | n2172 ;
  assign n2174 = n513 | n684 ;
  assign n2175 = n369 | n621 ;
  assign n2176 = n221 | n1252 ;
  assign n2177 = n448 | n2176 ;
  assign n2178 = n2175 | n2177 ;
  assign n2179 = n2174 | n2178 ;
  assign n2180 = n151 | n276 ;
  assign n2181 = n501 | n2180 ;
  assign n2182 = n486 | n491 ;
  assign n2183 = n690 | n2182 ;
  assign n2184 = n2181 | n2183 ;
  assign n2185 = n517 | n1047 ;
  assign n2186 = n205 | n257 ;
  assign n2187 = n2185 | n2186 ;
  assign n2188 = n2184 | n2187 ;
  assign n2189 = n2179 | n2188 ;
  assign n2190 = n2173 | n2189 ;
  assign n2191 = n530 | n870 ;
  assign n2192 = n272 | n520 ;
  assign n2193 = n900 | n2192 ;
  assign n2194 = n2191 | n2193 ;
  assign n2195 = n358 | n793 ;
  assign n2196 = n466 | n2195 ;
  assign n2197 = n291 | n2196 ;
  assign n2198 = n2072 | n2197 ;
  assign n2199 = n2194 | n2198 ;
  assign n2200 = n439 | n905 ;
  assign n2201 = n383 | n452 ;
  assign n2202 = n506 | n2201 ;
  assign n2203 = n112 | n399 ;
  assign n2204 = n345 | n477 ;
  assign n2205 = n2203 | n2204 ;
  assign n2206 = n2202 | n2205 ;
  assign n2207 = n2200 | n2206 ;
  assign n2208 = n116 | n249 ;
  assign n2209 = n220 | n548 ;
  assign n2210 = n2208 | n2209 ;
  assign n2211 = n1145 | n2210 ;
  assign n2212 = n2207 | n2211 ;
  assign n2213 = n2199 | n2212 ;
  assign n2214 = n2190 | n2213 ;
  assign n2215 = n2168 | n2214 ;
  assign n2216 = n2153 | n2215 ;
  assign n2217 = n2102 | n2216 ;
  assign n2222 = n2102 & n2216 ;
  assign n30124 = ~n2222 ;
  assign n2223 = n2217 & n30124 ;
  assign n2224 = n560 | n767 ;
  assign n2225 = n713 | n2224 ;
  assign n2226 = n107 | n989 ;
  assign n2227 = n1618 | n2226 ;
  assign n2228 = n2225 | n2227 ;
  assign n2229 = n157 | n368 ;
  assign n2230 = n263 | n461 ;
  assign n2231 = n280 | n668 ;
  assign n2232 = n2230 | n2231 ;
  assign n2233 = n2229 | n2232 ;
  assign n2234 = n133 | n162 ;
  assign n2235 = n492 | n2234 ;
  assign n2236 = n1477 | n2235 ;
  assign n2237 = n2233 | n2236 ;
  assign n2238 = n2228 | n2237 ;
  assign n2239 = n181 | n324 ;
  assign n2240 = n205 | n2239 ;
  assign n2241 = n464 | n469 ;
  assign n2242 = n875 | n2241 ;
  assign n2243 = n827 | n841 ;
  assign n2244 = n487 | n750 ;
  assign n2245 = n2243 | n2244 ;
  assign n2246 = n2242 | n2245 ;
  assign n2247 = n2240 | n2246 ;
  assign n2248 = n279 | n1384 ;
  assign n2249 = n601 | n1126 ;
  assign n2250 = n2248 | n2249 ;
  assign n2251 = n921 | n973 ;
  assign n2252 = n379 | n679 ;
  assign n2253 = n1760 | n2252 ;
  assign n2254 = n2251 | n2253 ;
  assign n2255 = n516 | n622 ;
  assign n2256 = n636 | n684 ;
  assign n2257 = n2255 | n2256 ;
  assign n2258 = n377 | n460 ;
  assign n2259 = n592 | n2258 ;
  assign n2260 = n2257 | n2259 ;
  assign n2261 = n2254 | n2260 ;
  assign n2262 = n2250 | n2261 ;
  assign n2263 = n2247 | n2262 ;
  assign n2264 = n2238 | n2263 ;
  assign n2265 = n366 | n793 ;
  assign n2266 = n203 | n257 ;
  assign n2267 = n512 | n2266 ;
  assign n2268 = n103 | n200 ;
  assign n2269 = n2123 | n2268 ;
  assign n2270 = n2267 | n2269 ;
  assign n2271 = n2265 | n2270 ;
  assign n2272 = n187 | n808 ;
  assign n2273 = n354 | n676 ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = n1066 | n2274 ;
  assign n2276 = n249 | n319 ;
  assign n2277 = n199 | n2276 ;
  assign n2278 = n2185 | n2277 ;
  assign n2279 = n2275 | n2278 ;
  assign n2280 = n348 | n476 ;
  assign n2281 = n857 | n2280 ;
  assign n2282 = n540 | n660 ;
  assign n2283 = n220 | n293 ;
  assign n2284 = n2282 | n2283 ;
  assign n2285 = n2281 | n2284 ;
  assign n2286 = n150 | n920 ;
  assign n2287 = n327 | n346 ;
  assign n2288 = n630 | n1010 ;
  assign n2289 = n2287 | n2288 ;
  assign n2290 = n2286 | n2289 ;
  assign n2291 = n2285 | n2290 ;
  assign n2292 = n2279 | n2291 ;
  assign n2293 = n2271 | n2292 ;
  assign n2294 = n459 | n2293 ;
  assign n2295 = n2264 | n2294 ;
  assign n2300 = n2216 | n2295 ;
  assign n2301 = n2216 & n2295 ;
  assign n30125 = ~n2301 ;
  assign n2302 = n2300 & n30125 ;
  assign n2303 = n1099 | n1109 ;
  assign n2304 = n1414 | n2303 ;
  assign n2305 = n205 | n369 ;
  assign n30126 = ~n368 ;
  assign n2306 = n145 & n30126 ;
  assign n30127 = ~n573 ;
  assign n2307 = n30127 & n2306 ;
  assign n30128 = ~n2305 ;
  assign n2308 = n30128 & n2307 ;
  assign n30129 = ~n2304 ;
  assign n2309 = n30129 & n2308 ;
  assign n2310 = n282 | n296 ;
  assign n2311 = n122 & n125 ;
  assign n2312 = n630 | n2311 ;
  assign n2313 = n2310 | n2312 ;
  assign n2314 = n398 | n2313 ;
  assign n2315 = n865 | n1825 ;
  assign n2316 = n331 | n658 ;
  assign n2317 = n124 | n2316 ;
  assign n2318 = n2315 | n2317 ;
  assign n2319 = n2314 | n2318 ;
  assign n102 = n96 | n101 ;
  assign n2320 = n82 & n102 ;
  assign n2321 = n273 | n405 ;
  assign n2322 = n2230 | n2321 ;
  assign n2323 = n2320 | n2322 ;
  assign n2324 = n446 | n532 ;
  assign n2325 = n236 | n335 ;
  assign n2326 = n224 | n487 ;
  assign n2327 = n2325 | n2326 ;
  assign n2328 = n2324 | n2327 ;
  assign n2329 = n2323 | n2328 ;
  assign n2330 = n2319 | n2329 ;
  assign n30130 = ~n2330 ;
  assign n2331 = n2309 & n30130 ;
  assign n30131 = ~n1436 ;
  assign n2332 = n30131 & n2331 ;
  assign n2333 = n476 | n925 ;
  assign n2334 = n472 | n2333 ;
  assign n2335 = n377 | n1249 ;
  assign n2336 = n1726 | n2045 ;
  assign n2337 = n2335 | n2336 ;
  assign n2338 = n1989 | n2337 ;
  assign n2339 = n2334 | n2338 ;
  assign n2340 = n292 | n496 ;
  assign n2341 = n1033 | n1413 ;
  assign n2342 = n2340 | n2341 ;
  assign n2343 = n223 | n432 ;
  assign n2344 = n676 | n2343 ;
  assign n2345 = n1238 | n2344 ;
  assign n2346 = n2342 | n2345 ;
  assign n2347 = n221 | n507 ;
  assign n2348 = n808 | n839 ;
  assign n2349 = n220 | n2348 ;
  assign n2350 = n2347 | n2349 ;
  assign n2351 = n277 | n1787 ;
  assign n2352 = n509 | n564 ;
  assign n2353 = n2351 | n2352 ;
  assign n2354 = n133 | n816 ;
  assign n2355 = n83 | n608 ;
  assign n2356 = n2354 | n2355 ;
  assign n2357 = n2353 | n2356 ;
  assign n2358 = n2350 | n2357 ;
  assign n2359 = n2346 | n2358 ;
  assign n2360 = n445 | n677 ;
  assign n2361 = n441 | n682 ;
  assign n2362 = n2360 | n2361 ;
  assign n2363 = n592 | n971 ;
  assign n2364 = n313 | n721 ;
  assign n2365 = n1050 | n2364 ;
  assign n2366 = n2363 | n2365 ;
  assign n2367 = n301 | n543 ;
  assign n2368 = n841 | n2367 ;
  assign n2369 = n233 | n298 ;
  assign n2370 = n2368 | n2369 ;
  assign n2371 = n2366 | n2370 ;
  assign n2372 = n2362 | n2371 ;
  assign n2373 = n2359 | n2372 ;
  assign n2374 = n2339 | n2373 ;
  assign n2375 = n1955 | n2374 ;
  assign n30132 = ~n2375 ;
  assign n2376 = n2332 & n30132 ;
  assign n30133 = ~n2295 ;
  assign n2379 = n30133 & n2376 ;
  assign n2378 = n2295 & n2376 ;
  assign n2380 = n2295 | n2376 ;
  assign n30134 = ~n2378 ;
  assign n2381 = n30134 & n2380 ;
  assign n2569 = n666 | n841 ;
  assign n2570 = n669 | n845 ;
  assign n2571 = n601 | n2570 ;
  assign n2572 = n2569 | n2571 ;
  assign n2573 = n371 | n417 ;
  assign n2574 = n1495 | n2229 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = n248 | n540 ;
  assign n2577 = n1252 | n2576 ;
  assign n2578 = n478 | n662 ;
  assign n2579 = n2577 | n2578 ;
  assign n2580 = n2575 | n2579 ;
  assign n2581 = n2572 | n2580 ;
  assign n2582 = n543 | n621 ;
  assign n2583 = n560 | n2582 ;
  assign n2584 = n324 | n439 ;
  assign n2585 = n971 | n2113 ;
  assign n2586 = n2584 | n2585 ;
  assign n2587 = n704 | n961 ;
  assign n2588 = n104 | n2587 ;
  assign n2589 = n840 | n905 ;
  assign n2590 = n2588 | n2589 ;
  assign n2591 = n2586 | n2590 ;
  assign n2592 = n2583 | n2591 ;
  assign n2593 = n312 | n453 ;
  assign n2594 = n416 | n2593 ;
  assign n2394 = n345 | n1129 ;
  assign n2595 = n1703 | n2394 ;
  assign n2596 = n2594 | n2595 ;
  assign n2597 = n763 | n2596 ;
  assign n2598 = n2592 | n2597 ;
  assign n2599 = n2581 | n2598 ;
  assign n2403 = n765 | n1047 ;
  assign n2404 = n785 | n1501 ;
  assign n2405 = n2403 | n2404 ;
  assign n2406 = n158 | n346 ;
  assign n2407 = n365 | n2406 ;
  assign n2408 = n176 | n221 ;
  assign n2409 = n2407 | n2408 ;
  assign n2410 = n479 | n509 ;
  assign n106 = n101 | n105 ;
  assign n2411 = n79 & n106 ;
  assign n2412 = n236 | n434 ;
  assign n2413 = n2411 | n2412 ;
  assign n2414 = n2410 | n2413 ;
  assign n2415 = n179 | n359 ;
  assign n2416 = n1010 | n2415 ;
  assign n2417 = n586 | n956 ;
  assign n2418 = n2416 | n2417 ;
  assign n2419 = n2414 | n2418 ;
  assign n2420 = n2409 | n2419 ;
  assign n2421 = n2405 | n2420 ;
  assign n2422 = n1304 | n2421 ;
  assign n2600 = n647 | n788 ;
  assign n2601 = n412 | n2600 ;
  assign n2602 = n282 | n1787 ;
  assign n2603 = n2601 | n2602 ;
  assign n2604 = n253 | n480 ;
  assign n2605 = n486 | n2604 ;
  assign n2606 = n220 | n630 ;
  assign n2607 = n470 | n2252 ;
  assign n2608 = n2606 | n2607 ;
  assign n2609 = n2605 | n2608 ;
  assign n2610 = n2603 | n2609 ;
  assign n2611 = n181 | n358 ;
  assign n2612 = n187 | n290 ;
  assign n2613 = n2611 | n2612 ;
  assign n2614 = n163 | n751 ;
  assign n2615 = n1423 | n2614 ;
  assign n2616 = n428 | n513 ;
  assign n2617 = n337 | n622 ;
  assign n2618 = n1421 | n2617 ;
  assign n2619 = n2616 | n2618 ;
  assign n2620 = n2615 | n2619 ;
  assign n2621 = n2613 | n2620 ;
  assign n2622 = n276 | n833 ;
  assign n2623 = n254 | n797 ;
  assign n2624 = n202 | n372 ;
  assign n2625 = n1437 | n2624 ;
  assign n2626 = n2623 | n2625 ;
  assign n2627 = n2622 | n2626 ;
  assign n2628 = n636 | n677 ;
  assign n2629 = n212 | n355 ;
  assign n2630 = n446 | n857 ;
  assign n2631 = n2629 | n2630 ;
  assign n2632 = n141 | n378 ;
  assign n2633 = n2631 | n2632 ;
  assign n2634 = n2628 | n2633 ;
  assign n2635 = n2627 | n2634 ;
  assign n2636 = n2621 | n2635 ;
  assign n2637 = n2610 | n2636 ;
  assign n2638 = n2422 | n2637 ;
  assign n2639 = n2599 | n2638 ;
  assign n2382 = n453 | n1252 ;
  assign n2383 = n141 | n2382 ;
  assign n2384 = n553 | n2052 ;
  assign n2385 = n2383 | n2384 ;
  assign n2386 = n916 | n1238 ;
  assign n2387 = n2385 | n2386 ;
  assign n30135 = ~n2387 ;
  assign n2388 = n1264 & n30135 ;
  assign n2389 = n302 | n508 ;
  assign n2390 = n334 | n407 ;
  assign n2391 = n461 | n2390 ;
  assign n2392 = n2389 | n2391 ;
  assign n2393 = n1057 | n2392 ;
  assign n2395 = n440 | n677 ;
  assign n2396 = n244 | n474 ;
  assign n2397 = n371 | n2396 ;
  assign n2398 = n2395 | n2397 ;
  assign n2399 = n2394 | n2398 ;
  assign n2400 = n2271 | n2399 ;
  assign n2401 = n2393 | n2400 ;
  assign n30136 = ~n2401 ;
  assign n2402 = n2388 & n30136 ;
  assign n2423 = n277 | n538 ;
  assign n2424 = n223 | n320 ;
  assign n2425 = n2423 | n2424 ;
  assign n2426 = n249 | n324 ;
  assign n2427 = n240 | n713 ;
  assign n2428 = n2426 | n2427 ;
  assign n2429 = n2425 | n2428 ;
  assign n2430 = n157 | n711 ;
  assign n2431 = n323 | n489 ;
  assign n2432 = n554 | n684 ;
  assign n2433 = n2431 | n2432 ;
  assign n2434 = n1477 | n2433 ;
  assign n2435 = n2430 | n2434 ;
  assign n2436 = n2429 | n2435 ;
  assign n2437 = n497 | n542 ;
  assign n2438 = n591 | n2437 ;
  assign n2439 = n1718 | n2438 ;
  assign n2440 = x26 | n29910 ;
  assign n2441 = n155 | n2440 ;
  assign n2442 = n73 & n2441 ;
  assign n260 = n155 | n259 ;
  assign n2443 = x25 | x26 ;
  assign n30137 = ~n2443 ;
  assign n2447 = n260 & n30137 ;
  assign n30138 = ~n2447 ;
  assign n2448 = n109 & n30138 ;
  assign n30139 = ~n2442 ;
  assign n2449 = n30139 & n2448 ;
  assign n2450 = n124 | n2449 ;
  assign n2451 = n506 | n668 ;
  assign n2452 = n168 | n621 ;
  assign n2453 = n2451 | n2452 ;
  assign n2454 = n2450 | n2453 ;
  assign n2455 = n2439 | n2454 ;
  assign n2456 = n767 | n978 ;
  assign n2457 = n383 | n2456 ;
  assign n2458 = n310 | n416 ;
  assign n2459 = n283 | n573 ;
  assign n2460 = n608 | n1091 ;
  assign n2461 = n2459 | n2460 ;
  assign n2462 = n2458 | n2461 ;
  assign n2463 = n2457 | n2462 ;
  assign n2464 = n921 | n1909 ;
  assign n2465 = n2140 | n2464 ;
  assign n2466 = n404 | n2465 ;
  assign n2467 = n2463 | n2466 ;
  assign n2468 = n2455 | n2467 ;
  assign n2469 = n2436 | n2468 ;
  assign n2470 = n2422 | n2469 ;
  assign n30140 = ~n2470 ;
  assign n2471 = n2402 & n30140 ;
  assign n2472 = n698 | n1787 ;
  assign n2473 = n324 | n506 ;
  assign n2474 = n2472 | n2473 ;
  assign n2475 = n138 | n346 ;
  assign n2476 = n722 | n2475 ;
  assign n2477 = n86 & n2447 ;
  assign n2478 = n477 | n516 ;
  assign n2479 = n2477 | n2478 ;
  assign n2480 = n2476 | n2479 ;
  assign n2481 = n112 | n473 ;
  assign n2482 = n996 | n2481 ;
  assign n2483 = n678 | n2482 ;
  assign n2484 = n2480 | n2483 ;
  assign n2485 = n2474 | n2484 ;
  assign n2486 = n223 | n1496 ;
  assign n2487 = n555 | n2486 ;
  assign n2488 = n1136 | n1689 ;
  assign n2489 = n660 | n1049 ;
  assign n2490 = n162 | n326 ;
  assign n2491 = n2489 | n2490 ;
  assign n2492 = n2488 | n2491 ;
  assign n2493 = n334 | n380 ;
  assign n2494 = n679 | n2493 ;
  assign n2495 = n384 | n751 ;
  assign n2497 = n2494 | n2495 ;
  assign n2498 = n2492 | n2497 ;
  assign n2499 = n2487 | n2498 ;
  assign n2500 = n157 | n412 ;
  assign n2501 = n853 | n2500 ;
  assign n2502 = n126 | n195 ;
  assign n2503 = n323 | n611 ;
  assign n2504 = n2502 | n2503 ;
  assign n2505 = n2501 | n2504 ;
  assign n2506 = n2334 | n2505 ;
  assign n2507 = n2499 | n2506 ;
  assign n2508 = n2485 | n2507 ;
  assign n2509 = n279 | n320 ;
  assign n2510 = n399 | n2509 ;
  assign n2511 = n550 | n764 ;
  assign n2512 = n337 | n451 ;
  assign n2513 = n2511 | n2512 ;
  assign n2514 = n2510 | n2513 ;
  assign n2515 = n418 | n845 ;
  assign n2516 = n1853 | n2515 ;
  assign n2517 = n961 | n1179 ;
  assign n2518 = n1688 | n2288 ;
  assign n2519 = n2517 | n2518 ;
  assign n2520 = n2516 | n2519 ;
  assign n2521 = n2514 | n2520 ;
  assign n2522 = n428 | n767 ;
  assign n2523 = n1047 | n2522 ;
  assign n2524 = n298 | n1252 ;
  assign n2525 = n190 | n517 ;
  assign n2526 = n1099 | n2525 ;
  assign n2527 = n2524 | n2526 ;
  assign n2528 = n2523 | n2527 ;
  assign n2529 = n479 | n797 ;
  assign n2530 = n1831 | n2529 ;
  assign n2531 = n1200 | n2122 ;
  assign n2532 = n366 | n486 ;
  assign n2533 = n2531 | n2532 ;
  assign n2534 = n2530 | n2533 ;
  assign n2535 = n2528 | n2534 ;
  assign n2536 = n2521 | n2535 ;
  assign n2537 = n104 | n271 ;
  assign n2538 = n510 | n1765 ;
  assign n2539 = n2537 | n2538 ;
  assign n2540 = n416 | n765 ;
  assign n2541 = n282 | n302 ;
  assign n2542 = n355 | n2541 ;
  assign n2543 = n1912 | n2542 ;
  assign n2544 = n2540 | n2543 ;
  assign n2545 = n2539 | n2544 ;
  assign n2546 = n512 | n635 ;
  assign n2547 = n1967 | n2546 ;
  assign n2548 = n1609 | n1879 ;
  assign n2549 = n2547 | n2548 ;
  assign n2550 = n572 | n586 ;
  assign n2551 = n1152 | n1497 ;
  assign n2552 = n2550 | n2551 ;
  assign n2553 = n150 | n300 ;
  assign n2554 = n983 | n2553 ;
  assign n2555 = n2552 | n2554 ;
  assign n30141 = ~n770 ;
  assign n2556 = n145 & n30141 ;
  assign n30142 = ~n2208 ;
  assign n2557 = n30142 & n2556 ;
  assign n2558 = n500 | n636 ;
  assign n170 = n127 | n169 ;
  assign n2559 = n110 & n170 ;
  assign n2560 = n2325 | n2559 ;
  assign n2561 = n2558 | n2560 ;
  assign n30143 = ~n2561 ;
  assign n2562 = n2557 & n30143 ;
  assign n30144 = ~n2555 ;
  assign n2563 = n30144 & n2562 ;
  assign n30145 = ~n2549 ;
  assign n2564 = n30145 & n2563 ;
  assign n30146 = ~n2545 ;
  assign n2565 = n30146 & n2564 ;
  assign n30147 = ~n2536 ;
  assign n2566 = n30147 & n2565 ;
  assign n30148 = ~n2508 ;
  assign n2567 = n30148 & n2566 ;
  assign n2640 = n2471 | n2567 ;
  assign n30149 = ~n2639 ;
  assign n2641 = n30149 & n2640 ;
  assign n2642 = n195 | n1047 ;
  assign n2643 = n1970 | n2412 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = n276 | n372 ;
  assign n2646 = n113 | n2645 ;
  assign n2647 = n455 | n2646 ;
  assign n2648 = n2644 | n2647 ;
  assign n2649 = n1131 | n2648 ;
  assign n2650 = n212 | n489 ;
  assign n2651 = n621 | n2650 ;
  assign n2652 = n2472 | n2651 ;
  assign n2653 = n233 | n594 ;
  assign n2654 = n255 | n396 ;
  assign n2655 = n2653 | n2654 ;
  assign n2656 = n2652 | n2655 ;
  assign n2657 = n200 | n345 ;
  assign n2658 = n841 | n2657 ;
  assign n2659 = n417 | n538 ;
  assign n2660 = n384 | n2659 ;
  assign n2661 = n2658 | n2660 ;
  assign n2662 = n1208 | n2661 ;
  assign n2663 = n2135 | n2662 ;
  assign n2664 = n2656 | n2663 ;
  assign n2665 = n2649 | n2664 ;
  assign n2666 = n688 | n2490 ;
  assign n2667 = n2617 | n2666 ;
  assign n2668 = n217 | n377 ;
  assign n2669 = n630 | n2668 ;
  assign n2670 = n244 | n383 ;
  assign n2671 = n542 | n1091 ;
  assign n2672 = n2670 | n2671 ;
  assign n2673 = n2315 | n2672 ;
  assign n2674 = n2669 | n2673 ;
  assign n2675 = n2667 | n2674 ;
  assign n2676 = n750 | n989 ;
  assign n2677 = n124 | n441 ;
  assign n2678 = n2676 | n2677 ;
  assign n2679 = n248 | n346 ;
  assign n2680 = n491 | n2679 ;
  assign n2681 = n282 | n1252 ;
  assign n2682 = n1430 | n2681 ;
  assign n2683 = n2680 | n2682 ;
  assign n2684 = n2678 | n2683 ;
  assign n2685 = n280 | n1179 ;
  assign n2686 = n273 | n501 ;
  assign n2687 = n151 | n651 ;
  assign n2688 = n2686 | n2687 ;
  assign n2689 = n2685 | n2688 ;
  assign n2690 = n138 | n179 ;
  assign n2691 = n379 | n2690 ;
  assign n2692 = n496 | n661 ;
  assign n2693 = n2691 | n2692 ;
  assign n2694 = n360 | n815 ;
  assign n2695 = n1267 | n2694 ;
  assign n2696 = n2693 | n2695 ;
  assign n2697 = n2689 | n2696 ;
  assign n2698 = n2684 | n2697 ;
  assign n2699 = n2675 | n2698 ;
  assign n30150 = ~n2699 ;
  assign n2700 = n940 & n30150 ;
  assign n30151 = ~n2665 ;
  assign n2701 = n30151 & n2700 ;
  assign n2702 = n2641 | n2701 ;
  assign n2703 = n301 | n954 ;
  assign n2704 = n1423 | n2703 ;
  assign n2705 = n162 | n176 ;
  assign n2706 = n195 | n2705 ;
  assign n2707 = n430 | n476 ;
  assign n2708 = n2160 | n2707 ;
  assign n2709 = n2706 | n2708 ;
  assign n2710 = n513 | n2138 ;
  assign n2711 = n240 | n534 ;
  assign n2712 = n2411 | n2711 ;
  assign n2713 = n2710 | n2712 ;
  assign n2714 = n2709 | n2713 ;
  assign n2715 = n2704 | n2714 ;
  assign n2716 = n344 | n418 ;
  assign n2717 = n187 | n621 ;
  assign n2718 = n540 | n682 ;
  assign n2719 = n610 | n2718 ;
  assign n2720 = n2717 | n2719 ;
  assign n2721 = n2716 | n2720 ;
  assign n2722 = n280 | n770 ;
  assign n2723 = n469 | n473 ;
  assign n2724 = n767 | n2723 ;
  assign n2725 = n2430 | n2724 ;
  assign n2726 = n2722 | n2725 ;
  assign n2727 = n2721 | n2726 ;
  assign n2728 = n2715 | n2727 ;
  assign n2729 = n140 | n811 ;
  assign n2730 = n698 | n2729 ;
  assign n2731 = n571 | n990 ;
  assign n2732 = n150 | n401 ;
  assign n2733 = n292 | n679 ;
  assign n2734 = n2732 | n2733 ;
  assign n2735 = n2731 | n2734 ;
  assign n2736 = n2730 | n2735 ;
  assign n2737 = n520 | n695 ;
  assign n2738 = n796 | n2737 ;
  assign n2739 = n991 | n1865 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n245 | n407 ;
  assign n2742 = n417 | n647 ;
  assign n2743 = n2741 | n2742 ;
  assign n2744 = n2200 | n2743 ;
  assign n2745 = n2740 | n2744 ;
  assign n2746 = n309 | n978 ;
  assign n2747 = n1066 | n2746 ;
  assign n2748 = n126 | n332 ;
  assign n2749 = n452 | n1091 ;
  assign n2750 = n1873 | n2749 ;
  assign n2751 = n2748 | n2750 ;
  assign n2752 = n2747 | n2751 ;
  assign n2753 = n2745 | n2752 ;
  assign n2754 = n2736 | n2753 ;
  assign n2755 = n2728 | n2754 ;
  assign n2756 = n151 | n190 ;
  assign n2757 = n460 | n2756 ;
  assign n2758 = n844 | n2757 ;
  assign n2759 = n103 | n479 ;
  assign n2760 = n2758 | n2759 ;
  assign n2761 = n609 | n2406 ;
  assign n2762 = n2540 | n2761 ;
  assign n2763 = n181 | n594 ;
  assign n2764 = n120 & n209 ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = n2762 | n2765 ;
  assign n2767 = n372 | n564 ;
  assign n2768 = n279 | n313 ;
  assign n2769 = n202 | n376 ;
  assign n2770 = n2768 | n2769 ;
  assign n2771 = n2767 | n2770 ;
  assign n2772 = n235 | n383 ;
  assign n2773 = n492 | n2772 ;
  assign n2774 = n1681 | n2773 ;
  assign n2775 = n2771 | n2774 ;
  assign n2776 = n2766 | n2775 ;
  assign n2777 = n2760 | n2776 ;
  assign n30152 = ~n2777 ;
  assign n2778 = n2331 & n30152 ;
  assign n30153 = ~n2755 ;
  assign n2779 = n30153 & n2778 ;
  assign n2786 = n2702 & n2779 ;
  assign n30154 = ~n2702 ;
  assign n2785 = n30154 & n2779 ;
  assign n30155 = ~n2471 ;
  assign n2794 = n30155 & n2639 ;
  assign n30156 = ~n2794 ;
  assign n2798 = n2701 & n30156 ;
  assign n30157 = ~n2779 ;
  assign n2799 = n30157 & n2798 ;
  assign n2800 = n2785 | n2799 ;
  assign n2801 = n2376 & n2800 ;
  assign n2802 = n2786 | n2801 ;
  assign n30158 = ~n2381 ;
  assign n2804 = n30158 & n2802 ;
  assign n2805 = n2379 | n2804 ;
  assign n2807 = n2302 & n2805 ;
  assign n30159 = ~n2807 ;
  assign n2808 = n2300 & n30159 ;
  assign n30160 = ~n2808 ;
  assign n2810 = n2223 & n30160 ;
  assign n30161 = ~n2810 ;
  assign n2811 = n2217 & n30161 ;
  assign n2812 = n2109 | n2811 ;
  assign n30162 = ~n2103 ;
  assign n2813 = n30162 & n2812 ;
  assign n30163 = ~n2813 ;
  assign n2815 = n2065 & n30163 ;
  assign n2816 = n2063 | n2815 ;
  assign n2817 = n1966 & n2816 ;
  assign n2818 = n1964 | n2817 ;
  assign n30164 = ~n1891 ;
  assign n2821 = n30164 & n2818 ;
  assign n2822 = n1888 | n2821 ;
  assign n30165 = ~n1819 ;
  assign n2823 = n30165 & n2822 ;
  assign n2824 = n1813 | n2823 ;
  assign n2827 = n1757 & n2824 ;
  assign n2828 = n1753 | n2827 ;
  assign n30166 = ~n1678 ;
  assign n2829 = n30166 & n2828 ;
  assign n2830 = n1676 | n2829 ;
  assign n2832 = n1564 & n2830 ;
  assign n30167 = ~n2832 ;
  assign n2833 = n1562 & n30167 ;
  assign n2834 = n1451 | n2833 ;
  assign n30168 = ~n1446 ;
  assign n2835 = n30168 & n2834 ;
  assign n2838 = n1343 | n2835 ;
  assign n30169 = ~n1337 ;
  assign n2839 = n30169 & n2838 ;
  assign n2840 = n1226 | n2839 ;
  assign n30170 = ~n1220 ;
  assign n2841 = n30170 & n2840 ;
  assign n30171 = ~n1082 ;
  assign n2842 = n30171 & n2841 ;
  assign n30172 = ~n2841 ;
  assign n2844 = n1082 & n30172 ;
  assign n2845 = n2842 | n2844 ;
  assign n30173 = ~n2845 ;
  assign n2846 = n895 & n30173 ;
  assign n30174 = ~n893 ;
  assign n894 = n891 & n30174 ;
  assign n1078 = n894 & n1074 ;
  assign n30175 = ~n30007 ;
  assign n153 = n30175 & n98 ;
  assign n30176 = ~n891 ;
  assign n2860 = n30176 & n893 ;
  assign n30177 = ~n153 ;
  assign n2861 = n30177 & n2860 ;
  assign n2864 = n1219 & n2861 ;
  assign n2875 = n1078 | n2864 ;
  assign n2849 = n153 & n30176 ;
  assign n2876 = n30074 & n2849 ;
  assign n2877 = n2875 | n2876 ;
  assign n2878 = n2846 | n2877 ;
  assign n30178 = ~n2878 ;
  assign n2879 = x29 & n30178 ;
  assign n2880 = n30024 & n2878 ;
  assign n2881 = n2879 | n2880 ;
  assign n2882 = n235 | n399 ;
  assign n2883 = n1787 | n2882 ;
  assign n2884 = n1047 | n2883 ;
  assign n2885 = n289 | n529 ;
  assign n2886 = n366 | n2885 ;
  assign n2887 = n163 | n272 ;
  assign n2888 = n2749 | n2887 ;
  assign n2889 = n2886 | n2888 ;
  assign n2890 = n1066 | n2582 ;
  assign n2891 = n2889 | n2890 ;
  assign n2892 = n2884 | n2891 ;
  assign n2893 = n200 | n433 ;
  assign n2894 = n550 | n2893 ;
  assign n2895 = n453 | n507 ;
  assign n2896 = n620 | n2895 ;
  assign n2897 = n2894 | n2896 ;
  assign n2898 = n765 | n996 ;
  assign n2899 = n1857 | n2898 ;
  assign n2900 = n174 | n808 ;
  assign n2901 = n517 | n682 ;
  assign n2902 = n2900 | n2901 ;
  assign n2903 = n2899 | n2902 ;
  assign n2904 = n1731 | n2769 ;
  assign n2905 = n151 | n248 ;
  assign n2906 = n139 | n461 ;
  assign n2907 = n2905 | n2906 ;
  assign n2908 = n2904 | n2907 ;
  assign n2909 = n592 | n788 ;
  assign n2910 = n1146 | n1574 ;
  assign n2911 = n2909 | n2910 ;
  assign n2912 = n2908 | n2911 ;
  assign n2913 = n2903 | n2912 ;
  assign n2914 = n2897 | n2913 ;
  assign n2915 = n2892 | n2914 ;
  assign n2916 = n1037 | n1853 ;
  assign n2917 = n865 | n900 ;
  assign n2918 = n282 | n332 ;
  assign n2919 = n181 | n764 ;
  assign n2920 = n2918 | n2919 ;
  assign n2921 = n2917 | n2920 ;
  assign n2922 = n2916 | n2921 ;
  assign n2923 = n162 | n214 ;
  assign n2924 = n1694 | n2412 ;
  assign n2925 = n2923 | n2924 ;
  assign n2926 = n80 | n319 ;
  assign n2927 = n688 | n2926 ;
  assign n2928 = n696 | n794 ;
  assign n2929 = n2927 | n2928 ;
  assign n2930 = n338 | n395 ;
  assign n2931 = n961 | n2930 ;
  assign n2932 = n983 | n2931 ;
  assign n2933 = n2929 | n2932 ;
  assign n2934 = n2925 | n2933 ;
  assign n2935 = n2922 | n2934 ;
  assign n2936 = n150 | n497 ;
  assign n2937 = n2013 | n2936 ;
  assign n2938 = n203 | n548 ;
  assign n2939 = n1321 | n2938 ;
  assign n2940 = n400 | n1252 ;
  assign n2941 = n126 | n326 ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = n2939 | n2942 ;
  assign n2944 = n220 | n647 ;
  assign n2945 = n658 | n1179 ;
  assign n2946 = n2944 | n2945 ;
  assign n2947 = n849 | n1294 ;
  assign n2948 = n2946 | n2947 ;
  assign n2949 = n2943 | n2948 ;
  assign n2950 = n2937 | n2949 ;
  assign n2951 = n302 | n635 ;
  assign n2952 = n186 | n368 ;
  assign n2953 = n2951 | n2952 ;
  assign n2954 = n668 | n978 ;
  assign n2955 = n331 | n554 ;
  assign n2956 = n2954 | n2955 ;
  assign n2957 = n2953 | n2956 ;
  assign n2958 = n279 | n827 ;
  assign n2959 = n572 | n2958 ;
  assign n2960 = n677 | n1200 ;
  assign n2961 = n2959 | n2960 ;
  assign n2962 = n239 | n560 ;
  assign n2963 = n2669 | n2962 ;
  assign n2964 = n2961 | n2963 ;
  assign n2965 = n2957 | n2964 ;
  assign n2966 = n432 | n477 ;
  assign n2967 = n679 | n2966 ;
  assign n2968 = n487 | n491 ;
  assign n2969 = n157 | n221 ;
  assign n2970 = n2968 | n2969 ;
  assign n2971 = n2967 | n2970 ;
  assign n2972 = n469 | n814 ;
  assign n2973 = n841 | n2972 ;
  assign n2974 = n90 | n989 ;
  assign n2975 = n1390 | n2974 ;
  assign n2976 = n2973 | n2975 ;
  assign n2977 = n2971 | n2976 ;
  assign n2978 = n2965 | n2977 ;
  assign n2979 = n2950 | n2978 ;
  assign n2980 = n2935 | n2979 ;
  assign n2981 = n2915 | n2980 ;
  assign n30179 = ~n2981 ;
  assign n2982 = x11 & n30179 ;
  assign n30180 = ~x11 ;
  assign n2983 = n30180 & n2981 ;
  assign n2984 = n2982 | n2983 ;
  assign n2985 = n107 | n553 ;
  assign n2986 = n235 | n293 ;
  assign n2987 = n326 | n2986 ;
  assign n2988 = n173 | n2987 ;
  assign n2989 = n2985 | n2988 ;
  assign n2990 = n452 | n1635 ;
  assign n2991 = n2364 | n2990 ;
  assign n2992 = n158 | n1047 ;
  assign n2993 = n528 | n651 ;
  assign n2994 = n1970 | n2993 ;
  assign n2995 = n2992 | n2994 ;
  assign n2996 = n2991 | n2995 ;
  assign n2997 = n2989 | n2996 ;
  assign n2998 = n335 | n517 ;
  assign n2999 = n1179 | n2998 ;
  assign n3000 = n476 | n1967 ;
  assign n3001 = n996 | n1787 ;
  assign n3002 = n2252 | n3001 ;
  assign n3003 = n3000 | n3002 ;
  assign n3004 = n2999 | n3003 ;
  assign n3005 = n1544 | n3004 ;
  assign n3006 = n2997 | n3005 ;
  assign n3007 = n2965 | n3006 ;
  assign n3008 = n376 | n636 ;
  assign n3009 = n282 | n520 ;
  assign n3010 = n3008 | n3009 ;
  assign n3011 = n1609 | n3010 ;
  assign n3012 = n1950 | n3011 ;
  assign n3013 = n263 | n410 ;
  assign n3014 = n2412 | n3013 ;
  assign n3015 = n550 | n647 ;
  assign n3016 = n704 | n925 ;
  assign n3017 = n3015 | n3016 ;
  assign n3018 = n3014 | n3017 ;
  assign n3019 = n564 | n622 ;
  assign n3020 = n2966 | n3019 ;
  assign n3021 = n1102 | n3020 ;
  assign n3022 = n610 | n764 ;
  assign n3023 = n216 | n3022 ;
  assign n3024 = n1725 | n3023 ;
  assign n3025 = n3021 | n3024 ;
  assign n3026 = n3018 | n3025 ;
  assign n3027 = n3012 | n3026 ;
  assign n3028 = n297 | n591 ;
  assign n3029 = n465 | n3028 ;
  assign n3030 = n1665 | n3029 ;
  assign n3031 = n202 | n383 ;
  assign n3032 = n1435 | n3031 ;
  assign n3033 = n2651 | n3032 ;
  assign n3034 = n3030 | n3033 ;
  assign n3035 = n1152 | n1860 ;
  assign n3036 = n2140 | n2320 ;
  assign n3037 = n3035 | n3036 ;
  assign n3038 = n2002 | n3037 ;
  assign n3039 = n291 | n1324 ;
  assign n3040 = n460 | n687 ;
  assign n3041 = n2203 | n2489 ;
  assign n3042 = n3040 | n3041 ;
  assign n3043 = n3039 | n3042 ;
  assign n3044 = n3038 | n3043 ;
  assign n3045 = n3034 | n3044 ;
  assign n3046 = n3027 | n3045 ;
  assign n3047 = n3007 | n3046 ;
  assign n30181 = ~n2984 ;
  assign n3048 = n30181 & n3047 ;
  assign n30182 = ~n3047 ;
  assign n3049 = n2984 & n30182 ;
  assign n3050 = n3048 | n3049 ;
  assign n3051 = n479 | n1049 ;
  assign n3052 = n205 | n431 ;
  assign n3053 = n3051 | n3052 ;
  assign n3054 = n354 | n446 ;
  assign n3055 = n647 | n3054 ;
  assign n3056 = n80 | n506 ;
  assign n3057 = n568 | n3056 ;
  assign n3058 = n3055 | n3057 ;
  assign n3059 = n3053 | n3058 ;
  assign n3060 = n513 | n516 ;
  assign n3061 = n410 | n651 ;
  assign n3062 = n767 | n3061 ;
  assign n3063 = n1100 | n3062 ;
  assign n3064 = n3060 | n3063 ;
  assign n3065 = n2092 | n3064 ;
  assign n3066 = n3059 | n3065 ;
  assign n3067 = n214 | n353 ;
  assign n3068 = n486 | n814 ;
  assign n3069 = n3067 | n3068 ;
  assign n3070 = n535 | n3069 ;
  assign n3071 = n929 | n3070 ;
  assign n3072 = n2758 | n3071 ;
  assign n3073 = n1462 | n3072 ;
  assign n3074 = n3066 | n3073 ;
  assign n3075 = n379 | n396 ;
  assign n3076 = n195 | n713 ;
  assign n3077 = n3075 | n3076 ;
  assign n3078 = n808 | n1422 ;
  assign n3079 = n784 | n3078 ;
  assign n3080 = n3077 | n3079 ;
  assign n3081 = n445 | n489 ;
  assign n3082 = n848 | n3081 ;
  assign n3083 = n355 | n417 ;
  assign n3084 = n764 | n3083 ;
  assign n3085 = n3082 | n3084 ;
  assign n3086 = n346 | n704 ;
  assign n3087 = n1101 | n3086 ;
  assign n3088 = n282 | n368 ;
  assign n3089 = n480 | n1179 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = n3087 | n3090 ;
  assign n3092 = n3085 | n3091 ;
  assign n3093 = n405 | n428 ;
  assign n3094 = n360 | n371 ;
  assign n3095 = n912 | n3094 ;
  assign n3096 = n3093 | n3095 ;
  assign n3097 = n1865 | n2411 ;
  assign n3098 = n432 | n560 ;
  assign n3099 = n312 | n636 ;
  assign n3100 = n3098 | n3099 ;
  assign n3101 = n3097 | n3100 ;
  assign n3102 = n3096 | n3101 ;
  assign n3103 = n3092 | n3102 ;
  assign n3104 = n3080 | n3103 ;
  assign n3105 = n1506 | n3104 ;
  assign n3106 = n1554 | n3105 ;
  assign n3107 = n3074 | n3106 ;
  assign n30183 = ~n3107 ;
  assign n3109 = n3047 & n30183 ;
  assign n3108 = n3047 | n3107 ;
  assign n3110 = n3047 & n3107 ;
  assign n30184 = ~n3110 ;
  assign n3111 = n3108 & n30184 ;
  assign n3112 = n80 | n1940 ;
  assign n3113 = n232 | n371 ;
  assign n3114 = n440 | n2311 ;
  assign n3115 = n3113 | n3114 ;
  assign n3116 = n833 | n905 ;
  assign n3117 = n497 | n532 ;
  assign n3118 = n506 | n548 ;
  assign n3119 = n3117 | n3118 ;
  assign n3120 = n3116 | n3119 ;
  assign n3121 = n3115 | n3120 ;
  assign n3122 = n3112 | n3121 ;
  assign n3123 = n921 | n2517 ;
  assign n3124 = n668 | n857 ;
  assign n3125 = n591 | n793 ;
  assign n3126 = n3124 | n3125 ;
  assign n3127 = n3123 | n3126 ;
  assign n3128 = n168 | n277 ;
  assign n3129 = n1510 | n3128 ;
  assign n3130 = n1472 | n2749 ;
  assign n3131 = n269 | n276 ;
  assign n3132 = n377 | n925 ;
  assign n3133 = n3131 | n3132 ;
  assign n3134 = n3130 | n3133 ;
  assign n3135 = n3129 | n3134 ;
  assign n3136 = n3127 | n3135 ;
  assign n3137 = n248 | n367 ;
  assign n3138 = n678 | n3137 ;
  assign n3139 = n610 | n1002 ;
  assign n3140 = n2962 | n3139 ;
  assign n3141 = n236 | n1495 ;
  assign n3142 = n167 | n445 ;
  assign n3143 = n1422 | n3142 ;
  assign n3144 = n3141 | n3143 ;
  assign n3145 = n3140 | n3144 ;
  assign n3146 = n3138 | n3145 ;
  assign n3147 = n3136 | n3146 ;
  assign n3148 = n3122 | n3147 ;
  assign n3149 = n1100 | n1361 ;
  assign n3150 = n241 | n495 ;
  assign n3151 = n797 | n3150 ;
  assign n3152 = n405 | n474 ;
  assign n3153 = n751 | n3152 ;
  assign n3154 = n3151 | n3153 ;
  assign n3155 = n3149 | n3154 ;
  assign n3156 = n848 | n1483 ;
  assign n3157 = n2389 | n3156 ;
  assign n3158 = n313 | n479 ;
  assign n3159 = n622 | n3158 ;
  assign n3160 = n853 | n3159 ;
  assign n3161 = n3157 | n3160 ;
  assign n3162 = n3155 | n3161 ;
  assign n3163 = n157 | n489 ;
  assign n3164 = n416 | n3163 ;
  assign n3165 = n138 | n163 ;
  assign n3166 = n126 | n573 ;
  assign n3167 = n3165 | n3166 ;
  assign n3168 = n3164 | n3167 ;
  assign n3169 = n2654 | n3168 ;
  assign n3170 = n200 | n1575 ;
  assign n3171 = n2968 | n3170 ;
  assign n3172 = n3060 | n3171 ;
  assign n3173 = n3169 | n3172 ;
  assign n3174 = n3162 | n3173 ;
  assign n3175 = n247 | n788 ;
  assign n3176 = n1050 | n1537 ;
  assign n3177 = n3175 | n3176 ;
  assign n3178 = n279 | n360 ;
  assign n3179 = n509 | n635 ;
  assign n3180 = n3178 | n3179 ;
  assign n3181 = n1032 | n3180 ;
  assign n3182 = n2717 | n3181 ;
  assign n3183 = n3177 | n3182 ;
  assign n3184 = n221 | n568 ;
  assign n3185 = n428 | n3184 ;
  assign n3186 = n1012 | n3185 ;
  assign n3187 = n900 | n1166 ;
  assign n3188 = n199 | n470 ;
  assign n3189 = n3187 | n3188 ;
  assign n3190 = n3186 | n3189 ;
  assign n3191 = n139 | n214 ;
  assign n3192 = n257 | n309 ;
  assign n3193 = n3191 | n3192 ;
  assign n3194 = n1123 | n3193 ;
  assign n3195 = n2605 | n2974 ;
  assign n3196 = n3194 | n3195 ;
  assign n3197 = n185 | n659 ;
  assign n3198 = n298 | n933 ;
  assign n3199 = n3197 | n3198 ;
  assign n3200 = n846 | n1497 ;
  assign n3201 = n721 | n1252 ;
  assign n3202 = n2511 | n3201 ;
  assign n3203 = n3200 | n3202 ;
  assign n3204 = n3199 | n3203 ;
  assign n3205 = n3196 | n3204 ;
  assign n3206 = n3190 | n3205 ;
  assign n3207 = n3183 | n3206 ;
  assign n3208 = n3174 | n3207 ;
  assign n3209 = n3148 | n3208 ;
  assign n30185 = ~x8 ;
  assign n3211 = n30185 & n3209 ;
  assign n30186 = ~n3209 ;
  assign n3210 = x8 & n30186 ;
  assign n3212 = n3210 | n3211 ;
  assign n3213 = n336 | n1049 ;
  assign n3214 = n216 | n811 ;
  assign n3215 = n2918 | n3214 ;
  assign n3216 = n3213 | n3215 ;
  assign n3217 = n1463 | n2157 ;
  assign n3218 = n2569 | n3217 ;
  assign n3219 = n3216 | n3218 ;
  assign n3220 = n214 | n319 ;
  assign n3221 = n290 | n3220 ;
  assign n3222 = n2894 | n3221 ;
  assign n3223 = n323 | n2517 ;
  assign n3224 = n293 | n1099 ;
  assign n3225 = n3223 | n3224 ;
  assign n3226 = n3222 | n3225 ;
  assign n3227 = n301 | n528 ;
  assign n3228 = n158 | n410 ;
  assign n3229 = n298 | n3228 ;
  assign n3230 = n3227 | n3229 ;
  assign n3231 = n1746 | n3230 ;
  assign n3232 = n3226 | n3231 ;
  assign n3233 = n80 | n453 ;
  assign n3234 = n460 | n3233 ;
  assign n3235 = n320 | n989 ;
  assign n3236 = n2326 | n3235 ;
  assign n3237 = n3234 | n3236 ;
  assign n3238 = n163 | n376 ;
  assign n3239 = n400 | n3238 ;
  assign n3240 = n126 | n383 ;
  assign n3241 = n1635 | n2052 ;
  assign n3242 = n3240 | n3241 ;
  assign n3243 = n3239 | n3242 ;
  assign n3244 = n3237 | n3243 ;
  assign n3245 = n3232 | n3244 ;
  assign n3246 = n3219 | n3245 ;
  assign n3247 = n174 | n568 ;
  assign n3248 = n1846 | n3247 ;
  assign n3249 = n681 | n2210 ;
  assign n3250 = n3248 | n3249 ;
  assign n3251 = n543 | n1047 ;
  assign n3252 = n157 | n159 ;
  assign n3253 = n439 | n3252 ;
  assign n3254 = n1566 | n3253 ;
  assign n3255 = n3251 | n3254 ;
  assign n3256 = n573 | n687 ;
  assign n3257 = n553 | n3256 ;
  assign n3258 = n2355 | n2711 ;
  assign n3259 = n3257 | n3258 ;
  assign n3260 = n501 | n3016 ;
  assign n3261 = n511 | n3260 ;
  assign n3262 = n3259 | n3261 ;
  assign n3263 = n3255 | n3262 ;
  assign n3264 = n3250 | n3263 ;
  assign n3265 = n358 | n379 ;
  assign n3266 = n440 | n695 ;
  assign n3267 = n3265 | n3266 ;
  assign n3268 = n327 | n452 ;
  assign n3269 = n431 | n3268 ;
  assign n3270 = n3267 | n3269 ;
  assign n3271 = n235 | n477 ;
  assign n3272 = n495 | n3271 ;
  assign n3273 = n398 | n3272 ;
  assign n3274 = n3270 | n3273 ;
  assign n3275 = n1129 | n2354 ;
  assign n3276 = n3131 | n3275 ;
  assign n3277 = n1763 | n3276 ;
  assign n3278 = n3274 | n3277 ;
  assign n3279 = n407 | n560 ;
  assign n3280 = n684 | n3279 ;
  assign n3281 = n372 | n491 ;
  assign n3282 = n698 | n3281 ;
  assign n3283 = n3280 | n3282 ;
  assign n3284 = n2133 | n3283 ;
  assign n3285 = n434 | n473 ;
  assign n3286 = n765 | n3285 ;
  assign n3287 = n296 | n399 ;
  assign n3288 = n412 | n3287 ;
  assign n3289 = n3286 | n3288 ;
  assign n3290 = n713 | n3117 ;
  assign n30187 = ~n3290 ;
  assign n3291 = n629 & n30187 ;
  assign n30188 = ~n3289 ;
  assign n3292 = n30188 & n3291 ;
  assign n30189 = ~n3284 ;
  assign n3293 = n30189 & n3292 ;
  assign n30190 = ~n3278 ;
  assign n3294 = n30190 & n3293 ;
  assign n30191 = ~n3264 ;
  assign n3295 = n30191 & n3294 ;
  assign n30192 = ~n3246 ;
  assign n3296 = n30192 & n3295 ;
  assign n3297 = n3212 | n3296 ;
  assign n30193 = ~n3211 ;
  assign n3298 = n30193 & n3297 ;
  assign n3299 = n3047 & n3298 ;
  assign n3300 = n3047 | n3298 ;
  assign n3304 = n1678 | n2828 ;
  assign n3306 = n1678 & n2828 ;
  assign n30194 = ~n3306 ;
  assign n3307 = n3304 & n30194 ;
  assign n3308 = n889 & n3307 ;
  assign n78 = x31 & n77 ;
  assign n3325 = x29 | x31 ;
  assign n30195 = ~n78 ;
  assign n3326 = n30195 & n3325 ;
  assign n3327 = x31 & n30022 ;
  assign n3328 = n29900 | n3327 ;
  assign n3329 = n3326 & n3328 ;
  assign n30196 = ~n1671 ;
  assign n3341 = n30196 & n3329 ;
  assign n30197 = ~x31 ;
  assign n3343 = n30197 & n108 ;
  assign n3355 = n1556 & n3343 ;
  assign n3357 = n3341 | n3355 ;
  assign n3311 = x31 & n29900 ;
  assign n3358 = n30105 & n3311 ;
  assign n3359 = n3357 | n3358 ;
  assign n3360 = n3308 | n3359 ;
  assign n30198 = ~n3360 ;
  assign n3361 = n3300 & n30198 ;
  assign n3362 = n3299 | n3361 ;
  assign n30199 = ~n3111 ;
  assign n3364 = n30199 & n3362 ;
  assign n3365 = n3109 | n3364 ;
  assign n3366 = n3050 | n3365 ;
  assign n3367 = n3050 & n3365 ;
  assign n30200 = ~n3367 ;
  assign n3368 = n3366 & n30200 ;
  assign n30201 = ~n1451 ;
  assign n3369 = n30201 & n2833 ;
  assign n30202 = ~n2833 ;
  assign n3370 = n1451 & n30202 ;
  assign n3371 = n3369 | n3370 ;
  assign n30203 = ~n3371 ;
  assign n3372 = n889 & n30203 ;
  assign n3322 = n1556 & n3311 ;
  assign n3339 = n1445 & n3329 ;
  assign n3375 = n3322 | n3339 ;
  assign n3376 = n30082 & n3343 ;
  assign n3377 = n3375 | n3376 ;
  assign n3378 = n3372 | n3377 ;
  assign n30204 = ~n3378 ;
  assign n3379 = n3368 & n30204 ;
  assign n30205 = ~n3368 ;
  assign n3380 = n30205 & n3378 ;
  assign n3381 = n3379 | n3380 ;
  assign n30206 = ~n3362 ;
  assign n3363 = n3111 & n30206 ;
  assign n3382 = n3363 | n3364 ;
  assign n30207 = ~n2830 ;
  assign n2831 = n1564 & n30207 ;
  assign n30208 = ~n1564 ;
  assign n3383 = n30208 & n2830 ;
  assign n3384 = n2831 | n3383 ;
  assign n30209 = ~n3384 ;
  assign n3385 = n889 & n30209 ;
  assign n3323 = n30196 & n3311 ;
  assign n3336 = n1556 & n3329 ;
  assign n3388 = n3323 | n3336 ;
  assign n3389 = n1445 & n3343 ;
  assign n3390 = n3388 | n3389 ;
  assign n3391 = n3385 | n3390 ;
  assign n3392 = n3382 | n3391 ;
  assign n30210 = ~n1226 ;
  assign n3393 = n30210 & n2839 ;
  assign n30211 = ~n2839 ;
  assign n3395 = n1226 & n30211 ;
  assign n3396 = n3393 | n3395 ;
  assign n30212 = ~n3396 ;
  assign n3397 = n895 & n30212 ;
  assign n1024 = n894 & n30074 ;
  assign n2866 = n30082 & n2861 ;
  assign n3400 = n1024 | n2866 ;
  assign n3401 = n1219 & n2849 ;
  assign n3402 = n3400 | n3401 ;
  assign n3403 = n3397 | n3402 ;
  assign n30213 = ~n3403 ;
  assign n3404 = x29 & n30213 ;
  assign n3405 = n30024 & n3403 ;
  assign n3406 = n3404 | n3405 ;
  assign n3407 = n3382 & n3391 ;
  assign n30214 = ~n3407 ;
  assign n3408 = n3392 & n30214 ;
  assign n30215 = ~n3406 ;
  assign n3409 = n30215 & n3408 ;
  assign n30216 = ~n3409 ;
  assign n3410 = n3392 & n30216 ;
  assign n30217 = ~n3381 ;
  assign n3411 = n30217 & n3410 ;
  assign n30218 = ~n3410 ;
  assign n3412 = n3381 & n30218 ;
  assign n3413 = n3411 | n3412 ;
  assign n30219 = ~n2881 ;
  assign n3414 = n30219 & n3413 ;
  assign n30220 = ~n3413 ;
  assign n3415 = n2881 & n30220 ;
  assign n3416 = n3414 | n3415 ;
  assign n30221 = ~n3408 ;
  assign n3417 = n3406 & n30221 ;
  assign n3418 = n3409 | n3417 ;
  assign n3419 = n3212 & n3296 ;
  assign n30222 = ~n3419 ;
  assign n3420 = n3297 & n30222 ;
  assign n3421 = n240 | n441 ;
  assign n3422 = n139 | n323 ;
  assign n3423 = n711 | n3422 ;
  assign n3424 = n3421 | n3423 ;
  assign n3425 = n248 | n2204 ;
  assign n3426 = n489 | n658 ;
  assign n3427 = n695 | n814 ;
  assign n3428 = n3426 | n3427 ;
  assign n3429 = n3425 | n3428 ;
  assign n3430 = n3424 | n3429 ;
  assign n3431 = n2091 | n3430 ;
  assign n3432 = n417 | n721 ;
  assign n3433 = n813 | n3432 ;
  assign n3434 = n854 | n3433 ;
  assign n3435 = n3039 | n3434 ;
  assign n3436 = n487 | n989 ;
  assign n3437 = n1100 | n1126 ;
  assign n3438 = n3436 | n3437 ;
  assign n3439 = n1426 | n3438 ;
  assign n3440 = n3435 | n3439 ;
  assign n3441 = n3431 | n3440 ;
  assign n3442 = n1230 | n1472 ;
  assign n3443 = n2324 | n3099 ;
  assign n3444 = n3442 | n3443 ;
  assign n3445 = n255 | n461 ;
  assign n3446 = n662 | n934 ;
  assign n3447 = n3445 | n3446 ;
  assign n3448 = n3444 | n3447 ;
  assign n3449 = n422 | n553 ;
  assign n3450 = n506 | n517 ;
  assign n3451 = n3449 | n3450 ;
  assign n3452 = n309 | n587 ;
  assign n3453 = n1152 | n3452 ;
  assign n3454 = n181 | n283 ;
  assign n3455 = n1271 | n3454 ;
  assign n3456 = n3453 | n3455 ;
  assign n3457 = n3451 | n3456 ;
  assign n3458 = n3448 | n3457 ;
  assign n3459 = n159 | n244 ;
  assign n3460 = n905 | n3459 ;
  assign n3461 = n235 | n249 ;
  assign n3462 = n371 | n767 ;
  assign n3463 = n3461 | n3462 ;
  assign n3464 = n103 | n220 ;
  assign n3465 = n381 | n3464 ;
  assign n3466 = n3463 | n3465 ;
  assign n3467 = n3460 | n3466 ;
  assign n3468 = n714 | n1857 ;
  assign n3469 = n2016 | n2410 ;
  assign n3470 = n3468 | n3469 ;
  assign n3471 = n3127 | n3470 ;
  assign n3472 = n3467 | n3471 ;
  assign n3473 = n3243 | n3472 ;
  assign n3474 = n2649 | n3473 ;
  assign n3475 = n3458 | n3474 ;
  assign n3476 = n3441 | n3475 ;
  assign n3478 = n3296 & n3476 ;
  assign n3477 = n3296 | n3476 ;
  assign n3479 = x2 | x5 ;
  assign n29885 = x2 & x5 ;
  assign n3480 = n399 | n480 ;
  assign n3481 = n2243 | n3051 ;
  assign n3482 = n3480 | n3481 ;
  assign n3483 = n283 | n446 ;
  assign n3484 = n996 | n3483 ;
  assign n3485 = n2317 | n3224 ;
  assign n3486 = n3484 | n3485 ;
  assign n3487 = n3482 | n3486 ;
  assign n3488 = n770 | n1010 ;
  assign n3489 = n272 | n453 ;
  assign n3490 = n540 | n3489 ;
  assign n3491 = n2186 | n3490 ;
  assign n3492 = n3488 | n3491 ;
  assign n3493 = n635 | n900 ;
  assign n3494 = n368 | n554 ;
  assign n3495 = n3493 | n3494 ;
  assign n3496 = n167 | n348 ;
  assign n3497 = n1928 | n2558 ;
  assign n3498 = n3496 | n3497 ;
  assign n3499 = n3495 | n3498 ;
  assign n3500 = n3492 | n3499 ;
  assign n3501 = n116 | n677 ;
  assign n3502 = n2767 | n3501 ;
  assign n3503 = n410 | n417 ;
  assign n3504 = n187 | n687 ;
  assign n3505 = n870 | n3504 ;
  assign n3506 = n3503 | n3505 ;
  assign n3507 = n300 | n309 ;
  assign n3508 = n369 | n591 ;
  assign n3509 = n3507 | n3508 ;
  assign n3510 = n158 | n174 ;
  assign n3511 = n780 | n3510 ;
  assign n3512 = n3509 | n3511 ;
  assign n3513 = n3506 | n3512 ;
  assign n3514 = n3502 | n3513 ;
  assign n3515 = n3500 | n3514 ;
  assign n3516 = n3487 | n3515 ;
  assign n3517 = n376 | n630 ;
  assign n3518 = n978 | n3517 ;
  assign n3519 = n232 | n244 ;
  assign n3520 = n781 | n3519 ;
  assign n3521 = n3518 | n3520 ;
  assign n3522 = n107 | n302 ;
  assign n3523 = n905 | n3522 ;
  assign n3524 = n464 | n679 ;
  assign n3525 = n814 | n3524 ;
  assign n3526 = n3523 | n3525 ;
  assign n3527 = n3521 | n3526 ;
  assign n3528 = n90 | n314 ;
  assign n3529 = n290 | n3528 ;
  assign n3530 = n452 | n529 ;
  assign n3531 = n676 | n3530 ;
  assign n3532 = n535 | n1200 ;
  assign n3533 = n3531 | n3532 ;
  assign n3534 = n3529 | n3533 ;
  assign n3535 = n130 | n276 ;
  assign n3536 = n1787 | n3535 ;
  assign n3537 = n439 | n865 ;
  assign n3538 = n313 | n793 ;
  assign n3539 = n3537 | n3538 ;
  assign n3540 = n3536 | n3539 ;
  assign n3541 = n1496 | n1717 ;
  assign n3542 = n1820 | n3201 ;
  assign n3543 = n3541 | n3542 ;
  assign n3544 = n3540 | n3543 ;
  assign n3545 = n3534 | n3544 ;
  assign n3546 = n3527 | n3545 ;
  assign n3547 = n176 | n765 ;
  assign n3548 = n186 | n989 ;
  assign n3549 = n3547 | n3548 ;
  assign n3550 = n451 | n517 ;
  assign n3551 = n542 | n795 ;
  assign n3552 = n3550 | n3551 ;
  assign n3553 = n355 | n396 ;
  assign n3554 = n273 | n319 ;
  assign n3555 = n3553 | n3554 ;
  assign n3556 = n3552 | n3555 ;
  assign n3557 = n759 | n3556 ;
  assign n3558 = n3549 | n3557 ;
  assign n3559 = n159 | n334 ;
  assign n3560 = n1766 | n3559 ;
  assign n3561 = n2517 | n3560 ;
  assign n3562 = n611 | n751 ;
  assign n3563 = n1129 | n3562 ;
  assign n3564 = n2601 | n3563 ;
  assign n3565 = n3561 | n3564 ;
  assign n3566 = n312 | n405 ;
  assign n3567 = n621 | n3566 ;
  assign n3568 = n80 | n401 ;
  assign n3569 = n1371 | n3568 ;
  assign n3570 = n3567 | n3569 ;
  assign n3571 = n299 | n3570 ;
  assign n3572 = n474 | n532 ;
  assign n3573 = n811 | n3572 ;
  assign n3574 = n203 | n258 ;
  assign n3575 = n301 | n430 ;
  assign n3576 = n3574 | n3575 ;
  assign n3577 = n3573 | n3576 ;
  assign n3578 = n622 | n666 ;
  assign n3579 = n150 | n433 ;
  assign n3580 = n3578 | n3579 ;
  assign n3581 = n3577 | n3580 ;
  assign n3582 = n3571 | n3581 ;
  assign n3583 = n3565 | n3582 ;
  assign n3584 = n3558 | n3583 ;
  assign n3585 = n3546 | n3584 ;
  assign n3586 = n3516 | n3585 ;
  assign n30223 = ~n29885 ;
  assign n3587 = n30223 & n3586 ;
  assign n30224 = ~n3587 ;
  assign n3588 = n3479 & n30224 ;
  assign n30225 = ~n3296 ;
  assign n3590 = n30225 & n3588 ;
  assign n30226 = ~n3588 ;
  assign n3589 = n3296 & n30226 ;
  assign n2819 = n1891 | n2818 ;
  assign n3591 = n1891 & n2818 ;
  assign n30227 = ~n3591 ;
  assign n3592 = n2819 & n30227 ;
  assign n3593 = n889 & n3592 ;
  assign n3321 = n30114 & n3311 ;
  assign n3337 = n30108 & n3329 ;
  assign n3596 = n3321 | n3337 ;
  assign n3597 = n1812 & n3343 ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n3593 | n3598 ;
  assign n3600 = n3589 | n3599 ;
  assign n30228 = ~n3590 ;
  assign n3601 = n30228 & n3600 ;
  assign n3602 = n3477 & n3601 ;
  assign n3603 = n3478 | n3602 ;
  assign n3605 = n3420 & n3603 ;
  assign n30229 = ~n3603 ;
  assign n3604 = n3420 & n30229 ;
  assign n30230 = ~n3420 ;
  assign n3606 = n30230 & n3603 ;
  assign n3607 = n3604 | n3606 ;
  assign n30231 = ~n2824 ;
  assign n2825 = n1757 & n30231 ;
  assign n30232 = ~n1757 ;
  assign n3608 = n30232 & n2824 ;
  assign n3609 = n2825 | n3608 ;
  assign n30233 = ~n3609 ;
  assign n3610 = n889 & n30233 ;
  assign n3316 = n1812 & n3311 ;
  assign n3354 = n30196 & n3343 ;
  assign n3613 = n3316 | n3354 ;
  assign n3614 = n30105 & n3329 ;
  assign n3615 = n3613 | n3614 ;
  assign n3616 = n3610 | n3615 ;
  assign n3618 = n3607 & n3616 ;
  assign n3619 = n3605 | n3618 ;
  assign n30234 = ~n3299 ;
  assign n3620 = n30234 & n3300 ;
  assign n3621 = n30198 & n3620 ;
  assign n30235 = ~n3620 ;
  assign n3622 = n3360 & n30235 ;
  assign n3623 = n3621 | n3622 ;
  assign n3625 = n3619 & n3623 ;
  assign n30236 = ~n1343 ;
  assign n2836 = n30236 & n2835 ;
  assign n30237 = ~n2835 ;
  assign n3626 = n1343 & n30237 ;
  assign n3627 = n2836 | n3626 ;
  assign n30238 = ~n3627 ;
  assign n3628 = n895 & n30238 ;
  assign n1222 = n894 & n1219 ;
  assign n2871 = n1445 & n2861 ;
  assign n3631 = n1222 | n2871 ;
  assign n3632 = n30082 & n2849 ;
  assign n3633 = n3631 | n3632 ;
  assign n3634 = n3628 | n3633 ;
  assign n3635 = x29 | n3634 ;
  assign n3636 = x29 & n3634 ;
  assign n30239 = ~n3636 ;
  assign n3637 = n3635 & n30239 ;
  assign n3624 = n3619 | n3623 ;
  assign n30240 = ~n3625 ;
  assign n3638 = n3624 & n30240 ;
  assign n3639 = n3637 & n3638 ;
  assign n3640 = n3625 | n3639 ;
  assign n3642 = n3418 & n3640 ;
  assign n3643 = n202 | n808 ;
  assign n3644 = n1573 | n3643 ;
  assign n3645 = n1092 | n1726 ;
  assign n3646 = n2360 | n3197 ;
  assign n3647 = n3645 | n3646 ;
  assign n3648 = n2760 | n3647 ;
  assign n3649 = n3644 | n3648 ;
  assign n3650 = n273 | n698 ;
  assign n3651 = n116 | n3650 ;
  assign n3652 = n318 | n1687 ;
  assign n3653 = n2923 | n3652 ;
  assign n3654 = n2185 | n3653 ;
  assign n3655 = n3651 | n3654 ;
  assign n3656 = n412 | n1243 ;
  assign n3657 = n2389 | n3247 ;
  assign n3658 = n3656 | n3657 ;
  assign n3659 = n232 | n381 ;
  assign n3660 = n853 | n3659 ;
  assign n3661 = n3658 | n3660 ;
  assign n3662 = n2747 | n3661 ;
  assign n3663 = n3655 | n3662 ;
  assign n3664 = n3649 | n3663 ;
  assign n3665 = n642 | n3129 ;
  assign n3666 = n324 | n405 ;
  assign n3667 = n636 | n3666 ;
  assign n3668 = n290 | n1859 ;
  assign n3669 = n3496 | n3668 ;
  assign n3670 = n3667 | n3669 ;
  assign n3671 = n960 | n3670 ;
  assign n3672 = n3665 | n3671 ;
  assign n3673 = n171 | n383 ;
  assign n3674 = n543 | n679 ;
  assign n3675 = n3673 | n3674 ;
  assign n3676 = n1597 | n3675 ;
  assign n3677 = n715 | n1996 ;
  assign n3678 = n112 | n1099 ;
  assign n3679 = n3090 | n3678 ;
  assign n3680 = n3677 | n3679 ;
  assign n3681 = n3676 | n3680 ;
  assign n3682 = n195 | n1199 ;
  assign n3683 = n205 | n240 ;
  assign n3684 = n1483 | n2051 ;
  assign n3685 = n3683 | n3684 ;
  assign n3686 = n3682 | n3685 ;
  assign n3687 = n464 | n839 ;
  assign n3688 = n921 | n3687 ;
  assign n3689 = n1129 | n3688 ;
  assign n3690 = n399 | n418 ;
  assign n3691 = n506 | n647 ;
  assign n3692 = n3690 | n3691 ;
  assign n3693 = n323 | n376 ;
  assign n3694 = n1495 | n3693 ;
  assign n3695 = n3692 | n3694 ;
  assign n3696 = n3689 | n3695 ;
  assign n3697 = n3686 | n3696 ;
  assign n3698 = n3681 | n3697 ;
  assign n3699 = n3672 | n3698 ;
  assign n3700 = n3664 | n3699 ;
  assign n3710 = n661 | n920 ;
  assign n3711 = n1114 | n3710 ;
  assign n3712 = n512 | n564 ;
  assign n3713 = n568 | n3712 ;
  assign n3714 = n365 | n508 ;
  assign n3715 = n141 | n3714 ;
  assign n3716 = n3713 | n3715 ;
  assign n3717 = n771 | n1853 ;
  assign n3718 = n3716 | n3717 ;
  assign n3719 = n3711 | n3718 ;
  assign n3720 = n293 | n358 ;
  assign n3721 = n687 | n3720 ;
  assign n3722 = n223 | n257 ;
  assign n3723 = n1688 | n3722 ;
  assign n3724 = n3721 | n3723 ;
  assign n3725 = n1006 | n3724 ;
  assign n3726 = n2763 | n3425 ;
  assign n3727 = n202 | n349 ;
  assign n3728 = n764 | n3727 ;
  assign n3729 = n573 | n698 ;
  assign n3730 = n3728 | n3729 ;
  assign n3731 = n3726 | n3730 ;
  assign n3732 = n3725 | n3731 ;
  assign n3733 = n3719 | n3732 ;
  assign n3734 = n290 | n395 ;
  assign n3735 = n982 | n3734 ;
  assign n3736 = n258 | n327 ;
  assign n3737 = n711 | n3736 ;
  assign n3738 = n130 | n1423 ;
  assign n3739 = n3737 | n3738 ;
  assign n3740 = n3735 | n3739 ;
  assign n3741 = n381 | n433 ;
  assign n3742 = n1731 | n2938 ;
  assign n3743 = n3741 | n3742 ;
  assign n3744 = n662 | n2746 ;
  assign n3745 = n3132 | n3744 ;
  assign n3746 = n3743 | n3745 ;
  assign n3747 = n3740 | n3746 ;
  assign n3748 = n126 | n167 ;
  assign n3749 = n334 | n3748 ;
  assign n3750 = n353 | n469 ;
  assign n3751 = n797 | n3750 ;
  assign n3752 = n3749 | n3751 ;
  assign n3753 = n319 | n666 ;
  assign n3754 = n270 | n677 ;
  assign n3755 = n3753 | n3754 ;
  assign n3756 = n3752 | n3755 ;
  assign n3757 = n232 | n668 ;
  assign n3758 = n602 | n3757 ;
  assign n3759 = n1918 | n3758 ;
  assign n3760 = n1411 | n3759 ;
  assign n3761 = n3756 | n3760 ;
  assign n3762 = n3747 | n3761 ;
  assign n3763 = n1780 | n3762 ;
  assign n3764 = n3733 | n3763 ;
  assign n3765 = n3700 | n3764 ;
  assign n3774 = n3700 & n3764 ;
  assign n30241 = ~n3774 ;
  assign n3775 = n3765 & n30241 ;
  assign n3776 = n1074 | n3764 ;
  assign n30242 = ~n3764 ;
  assign n3773 = n1074 & n30242 ;
  assign n30243 = ~n1074 ;
  assign n3777 = n30243 & n3764 ;
  assign n3778 = n3773 | n3777 ;
  assign n3779 = n1023 & n30243 ;
  assign n3780 = n1082 | n2841 ;
  assign n30244 = ~n3779 ;
  assign n3781 = n30244 & n3780 ;
  assign n30245 = ~n3781 ;
  assign n3783 = n3778 & n30245 ;
  assign n30246 = ~n3783 ;
  assign n3784 = n3776 & n30246 ;
  assign n30247 = ~n3784 ;
  assign n3785 = n3775 & n30247 ;
  assign n30248 = ~n3775 ;
  assign n3786 = n30248 & n3784 ;
  assign n3787 = n3785 | n3786 ;
  assign n30249 = ~n37283 ;
  assign n2444 = n30249 & n2443 ;
  assign n3791 = n260 & n2444 ;
  assign n3798 = n3787 & n3791 ;
  assign n1080 = n209 & n1074 ;
  assign n30250 = ~n2444 ;
  assign n3818 = n260 & n30250 ;
  assign n3830 = n3700 & n3818 ;
  assign n3835 = n1080 | n3830 ;
  assign n30251 = ~n29910 ;
  assign n121 = n30251 & n73 ;
  assign n30252 = ~n260 ;
  assign n3802 = n121 & n30252 ;
  assign n3836 = n3764 & n3802 ;
  assign n3837 = n3835 | n3836 ;
  assign n3838 = n3798 | n3837 ;
  assign n30253 = ~n3838 ;
  assign n3839 = x26 & n30253 ;
  assign n3840 = n30019 & n3838 ;
  assign n3841 = n3839 | n3840 ;
  assign n3641 = n3418 | n3640 ;
  assign n30254 = ~n3642 ;
  assign n3842 = n3641 & n30254 ;
  assign n3844 = n3841 & n3842 ;
  assign n3845 = n3642 | n3844 ;
  assign n3846 = n3416 | n3845 ;
  assign n3847 = n3416 & n3845 ;
  assign n30255 = ~n3847 ;
  assign n3848 = n3846 & n30255 ;
  assign n3849 = n116 | n797 ;
  assign n3850 = n1821 | n3166 ;
  assign n3851 = n3849 | n3850 ;
  assign n3852 = n313 | n470 ;
  assign n3853 = n186 | n301 ;
  assign n3854 = n795 | n857 ;
  assign n3855 = n3853 | n3854 ;
  assign n3856 = n3852 | n3855 ;
  assign n3857 = n3851 | n3856 ;
  assign n3858 = n1266 | n3857 ;
  assign n3859 = n3644 | n3858 ;
  assign n30256 = ~n986 ;
  assign n3860 = n909 & n30256 ;
  assign n30257 = ~n3859 ;
  assign n3861 = n30257 & n3860 ;
  assign n3862 = n30151 & n3861 ;
  assign n30258 = ~n3074 ;
  assign n3863 = n30258 & n3862 ;
  assign n3866 = n3700 & n3863 ;
  assign n3867 = n3700 | n3863 ;
  assign n30259 = ~n3866 ;
  assign n3868 = n30259 & n3867 ;
  assign n30260 = ~n3785 ;
  assign n3869 = n3765 & n30260 ;
  assign n30261 = ~n3868 ;
  assign n3870 = n30261 & n3869 ;
  assign n30262 = ~n3869 ;
  assign n3871 = n3868 & n30262 ;
  assign n3872 = n3870 | n3871 ;
  assign n30263 = ~n3872 ;
  assign n3873 = n3791 & n30263 ;
  assign n3768 = n209 & n3764 ;
  assign n3808 = n3700 & n3802 ;
  assign n3877 = n3768 | n3808 ;
  assign n30264 = ~n3863 ;
  assign n3878 = n3818 & n30264 ;
  assign n3879 = n3877 | n3878 ;
  assign n3880 = n3873 | n3879 ;
  assign n30265 = ~n3880 ;
  assign n3881 = x26 & n30265 ;
  assign n3882 = n30019 & n3880 ;
  assign n3883 = n3881 | n3882 ;
  assign n30266 = ~n3883 ;
  assign n3884 = n3848 & n30266 ;
  assign n30267 = ~n3848 ;
  assign n3885 = n30267 & n3883 ;
  assign n3886 = n3884 | n3885 ;
  assign n3887 = n666 | n750 ;
  assign n3888 = n225 | n696 ;
  assign n3889 = n2600 | n3888 ;
  assign n3890 = n3887 | n3889 ;
  assign n3891 = n978 | n2016 ;
  assign n30268 = ~n337 ;
  assign n3892 = n145 & n30268 ;
  assign n30269 = ~n3201 ;
  assign n3893 = n30269 & n3892 ;
  assign n30270 = ~n3891 ;
  assign n3894 = n30270 & n3893 ;
  assign n3895 = n773 | n2200 ;
  assign n30271 = ~n3895 ;
  assign n3896 = n3894 & n30271 ;
  assign n3897 = n509 | n520 ;
  assign n3898 = n844 | n3897 ;
  assign n3899 = n2139 | n2389 ;
  assign n3900 = n3898 | n3899 ;
  assign n3901 = n2350 | n3900 ;
  assign n30272 = ~n3901 ;
  assign n3902 = n3896 & n30272 ;
  assign n30273 = ~n3890 ;
  assign n3903 = n30273 & n3902 ;
  assign n30274 = ~n2736 ;
  assign n3904 = n30274 & n3903 ;
  assign n3905 = n124 | n591 ;
  assign n3906 = n276 | n412 ;
  assign n3907 = n1141 | n3906 ;
  assign n3908 = n3905 | n3907 ;
  assign n3909 = n920 | n1346 ;
  assign n3910 = n2231 | n3909 ;
  assign n3911 = n474 | n1199 ;
  assign n3912 = n535 | n3911 ;
  assign n3913 = n722 | n846 ;
  assign n3914 = n3912 | n3913 ;
  assign n3915 = n385 | n955 ;
  assign n3916 = n3914 | n3915 ;
  assign n3917 = n3910 | n3916 ;
  assign n3918 = n3908 | n3917 ;
  assign n3919 = n771 | n2248 ;
  assign n3920 = n3493 | n3919 ;
  assign n3921 = n270 | n335 ;
  assign n3922 = n159 | n432 ;
  assign n3923 = n2748 | n3922 ;
  assign n3924 = n3921 | n3923 ;
  assign n3925 = n1147 | n1423 ;
  assign n3926 = n1435 | n1892 ;
  assign n3927 = n3925 | n3926 ;
  assign n3928 = n441 | n489 ;
  assign n3929 = n793 | n3928 ;
  assign n3930 = n83 | n369 ;
  assign n3931 = n237 | n3930 ;
  assign n3932 = n3929 | n3931 ;
  assign n3933 = n3927 | n3932 ;
  assign n3934 = n3924 | n3933 ;
  assign n3935 = n3920 | n3934 ;
  assign n3936 = n1839 | n3935 ;
  assign n3937 = n3918 | n3936 ;
  assign n30275 = ~n3937 ;
  assign n3938 = n3904 & n30275 ;
  assign n3948 = n107 | n445 ;
  assign n3949 = n214 | n1058 ;
  assign n3950 = n3948 | n3949 ;
  assign n3951 = n174 | n480 ;
  assign n3952 = n925 | n3951 ;
  assign n3953 = n780 | n1856 ;
  assign n3954 = n2282 | n2525 ;
  assign n3955 = n3953 | n3954 ;
  assign n3956 = n3952 | n3955 ;
  assign n3957 = n3950 | n3956 ;
  assign n3958 = n2653 | n3684 ;
  assign n3959 = n235 | n430 ;
  assign n3960 = n460 | n543 ;
  assign n3961 = n3959 | n3960 ;
  assign n3962 = n186 | n446 ;
  assign n3963 = n689 | n3962 ;
  assign n3964 = n3961 | n3963 ;
  assign n3965 = n3958 | n3964 ;
  assign n3966 = n159 | n957 ;
  assign n3967 = n248 | n682 ;
  assign n3968 = n80 | n313 ;
  assign n3969 = n3967 | n3968 ;
  assign n3970 = n3966 | n3969 ;
  assign n2496 = n378 | n384 ;
  assign n3971 = n533 | n572 ;
  assign n3972 = n2496 | n3971 ;
  assign n3973 = n319 | n366 ;
  assign n3974 = n1853 | n3973 ;
  assign n3975 = n3972 | n3974 ;
  assign n3976 = n3970 | n3975 ;
  assign n3977 = n3965 | n3976 ;
  assign n3978 = n3957 | n3977 ;
  assign n3979 = n217 | n453 ;
  assign n3980 = n477 | n845 ;
  assign n3981 = n3979 | n3980 ;
  assign n3982 = n853 | n3981 ;
  assign n3983 = n1846 | n1912 ;
  assign n3984 = n3982 | n3983 ;
  assign n3985 = n221 | n332 ;
  assign n3986 = n3197 | n3985 ;
  assign n3987 = n621 | n794 ;
  assign n3988 = n2016 | n3987 ;
  assign n3989 = n3986 | n3988 ;
  assign n3990 = n3984 | n3989 ;
  assign n3991 = n97 | n401 ;
  assign n3992 = n1688 | n3991 ;
  assign n3993 = n335 | n611 ;
  assign n3994 = n1683 | n3993 ;
  assign n3995 = n3992 | n3994 ;
  assign n3996 = n1948 | n2154 ;
  assign n3997 = n302 | n722 ;
  assign n3998 = n2163 | n3997 ;
  assign n3999 = n3996 | n3998 ;
  assign n4000 = n3995 | n3999 ;
  assign n4001 = n3990 | n4000 ;
  assign n4002 = n1028 | n2941 ;
  assign n4003 = n3422 | n4002 ;
  assign n4004 = n976 | n990 ;
  assign n4005 = n695 | n770 ;
  assign n4006 = n1776 | n4005 ;
  assign n4007 = n4004 | n4006 ;
  assign n4008 = n4003 | n4007 ;
  assign n4009 = n418 | n1689 ;
  assign n4010 = n314 | n622 ;
  assign n4011 = n432 | n630 ;
  assign n4012 = n4010 | n4011 ;
  assign n4013 = n539 | n4012 ;
  assign n4014 = n4009 | n4013 ;
  assign n4015 = n501 | n1049 ;
  assign n4016 = n381 | n4015 ;
  assign n4017 = n1681 | n4016 ;
  assign n4018 = n396 | n534 ;
  assign n4019 = n1531 | n4018 ;
  assign n4020 = n245 | n797 ;
  assign n4021 = n4019 | n4020 ;
  assign n4022 = n4017 | n4021 ;
  assign n4023 = n554 | n591 ;
  assign n4024 = n827 | n4023 ;
  assign n4025 = n479 | n548 ;
  assign n4026 = n195 | n4025 ;
  assign n4027 = n4024 | n4026 ;
  assign n4028 = n2523 | n4027 ;
  assign n4029 = n4022 | n4028 ;
  assign n4030 = n4014 | n4029 ;
  assign n4031 = n4008 | n4030 ;
  assign n4032 = n4001 | n4031 ;
  assign n4033 = n3978 | n4032 ;
  assign n4037 = n222 | n1249 ;
  assign n4038 = n1596 | n4037 ;
  assign n4039 = n290 | n360 ;
  assign n4040 = n83 | n338 ;
  assign n4041 = n422 | n4040 ;
  assign n4042 = n2502 | n4041 ;
  assign n4043 = n4039 | n4042 ;
  assign n4044 = n4038 | n4043 ;
  assign n4045 = n224 | n554 ;
  assign n4046 = n2113 | n4045 ;
  assign n4047 = n130 | n365 ;
  assign n4048 = n3131 | n4047 ;
  assign n4049 = n4046 | n4048 ;
  assign n4050 = n1642 | n2601 ;
  assign n4051 = n4049 | n4050 ;
  assign n4052 = n417 | n1422 ;
  assign n4053 = n1487 | n2732 ;
  assign n4054 = n4052 | n4053 ;
  assign n4055 = n368 | n587 ;
  assign n4056 = n272 | n564 ;
  assign n4057 = n989 | n4056 ;
  assign n4058 = n4055 | n4057 ;
  assign n4059 = n189 | n294 ;
  assign n4060 = n4058 | n4059 ;
  assign n4061 = n4054 | n4060 ;
  assign n4062 = n4051 | n4061 ;
  assign n4063 = n4044 | n4062 ;
  assign n4064 = n349 | n418 ;
  assign n4065 = n501 | n1091 ;
  assign n4066 = n4064 | n4065 ;
  assign n4067 = n204 | n722 ;
  assign n4068 = n4066 | n4067 ;
  assign n4069 = n273 | n344 ;
  assign n4070 = n3223 | n4069 ;
  assign n4071 = n4068 | n4070 ;
  assign n4072 = n452 | n982 ;
  assign n4073 = n217 | n573 ;
  assign n4074 = n326 | n410 ;
  assign n4075 = n2288 | n4074 ;
  assign n4076 = n4073 | n4075 ;
  assign n4077 = n4072 | n4076 ;
  assign n4078 = n4071 | n4077 ;
  assign n4079 = n1434 | n4078 ;
  assign n4080 = n163 | n318 ;
  assign n4081 = n310 | n4080 ;
  assign n4082 = n510 | n533 ;
  assign n4083 = n4081 | n4082 ;
  assign n4084 = n3251 | n4083 ;
  assign n4085 = n931 | n1050 ;
  assign n4086 = n451 | n560 ;
  assign n4087 = n3214 | n4086 ;
  assign n4088 = n4085 | n4087 ;
  assign n4089 = n2086 | n4088 ;
  assign n4090 = n2903 | n4089 ;
  assign n4091 = n4084 | n4090 ;
  assign n4092 = n4079 | n4091 ;
  assign n4093 = n4063 | n4092 ;
  assign n30276 = ~n4093 ;
  assign n4107 = n3863 & n30276 ;
  assign n30277 = ~n3700 ;
  assign n4108 = n30277 & n3863 ;
  assign n4109 = n3868 | n3869 ;
  assign n30278 = ~n4108 ;
  assign n4110 = n30278 & n4109 ;
  assign n4100 = n3863 & n4093 ;
  assign n4111 = n3863 | n4093 ;
  assign n30279 = ~n4100 ;
  assign n4112 = n30279 & n4111 ;
  assign n4113 = n4110 | n4112 ;
  assign n30280 = ~n4107 ;
  assign n4114 = n30280 & n4113 ;
  assign n4115 = n4093 & n4114 ;
  assign n4117 = n4033 | n4115 ;
  assign n4118 = n4093 | n4114 ;
  assign n4119 = n4033 & n4118 ;
  assign n30281 = ~n4119 ;
  assign n4121 = n4117 & n30281 ;
  assign n30282 = ~n3938 ;
  assign n4122 = n30282 & n4121 ;
  assign n30283 = ~n4121 ;
  assign n4123 = n3938 & n30283 ;
  assign n4124 = n4122 | n4123 ;
  assign n29890 = x20 & x21 ;
  assign n4129 = x20 | x21 ;
  assign n30284 = ~n29890 ;
  assign n4132 = n30284 & n4129 ;
  assign n37286 = x22 & x23 ;
  assign n4133 = x22 | x23 ;
  assign n30285 = ~n37286 ;
  assign n4134 = n30285 & n4133 ;
  assign n4135 = n4132 & n4134 ;
  assign n30286 = ~n4124 ;
  assign n4142 = n30286 & n4135 ;
  assign n30287 = ~n4134 ;
  assign n4165 = n4132 & n30287 ;
  assign n4176 = n30282 & n4165 ;
  assign n30288 = ~n4129 ;
  assign n4130 = x22 & n30288 ;
  assign n30289 = ~x22 ;
  assign n4147 = n30289 & n29890 ;
  assign n4148 = n4130 | n4147 ;
  assign n4183 = n4132 | n4148 ;
  assign n30290 = ~n4183 ;
  assign n4185 = n4134 & n30290 ;
  assign n4200 = n4093 & n4185 ;
  assign n4204 = n4176 | n4200 ;
  assign n4205 = n4033 & n4148 ;
  assign n4206 = n4204 | n4205 ;
  assign n4207 = n4142 | n4206 ;
  assign n4208 = x23 | n4207 ;
  assign n4209 = x23 & n4207 ;
  assign n30291 = ~n4209 ;
  assign n4210 = n4208 & n30291 ;
  assign n30292 = ~n3886 ;
  assign n4211 = n30292 & n4210 ;
  assign n30293 = ~n4210 ;
  assign n4212 = n3886 & n30293 ;
  assign n4213 = n4211 | n4212 ;
  assign n30294 = ~n3841 ;
  assign n3843 = n30294 & n3842 ;
  assign n30295 = ~n3842 ;
  assign n4214 = n3841 & n30295 ;
  assign n4215 = n3843 | n4214 ;
  assign n4216 = n3637 | n3638 ;
  assign n30296 = ~n3639 ;
  assign n4217 = n30296 & n4216 ;
  assign n3373 = n895 & n30203 ;
  assign n1339 = n894 & n30082 ;
  assign n2869 = n1556 & n2861 ;
  assign n4218 = n1339 | n2869 ;
  assign n4219 = n1445 & n2849 ;
  assign n4220 = n4218 | n4219 ;
  assign n4221 = n3373 | n4220 ;
  assign n4222 = x29 | n4221 ;
  assign n4223 = x29 & n4221 ;
  assign n30297 = ~n4223 ;
  assign n4224 = n4222 & n30297 ;
  assign n30298 = ~n3478 ;
  assign n4225 = n3477 & n30298 ;
  assign n4226 = n3601 & n4225 ;
  assign n4227 = n3601 | n4225 ;
  assign n30299 = ~n4226 ;
  assign n4228 = n30299 & n4227 ;
  assign n3303 = n1819 | n2822 ;
  assign n4229 = n1819 & n2822 ;
  assign n30300 = ~n4229 ;
  assign n4230 = n3303 & n30300 ;
  assign n4231 = n889 & n4230 ;
  assign n3333 = n1812 & n3329 ;
  assign n3353 = n30105 & n3343 ;
  assign n4236 = n3333 | n3353 ;
  assign n4237 = n30108 & n3311 ;
  assign n4238 = n4236 | n4237 ;
  assign n4239 = n4231 | n4238 ;
  assign n4240 = n4228 | n4239 ;
  assign n4241 = n492 | n569 ;
  assign n4242 = n1928 | n2584 ;
  assign n4243 = n4241 | n4242 ;
  assign n4244 = n185 | n445 ;
  assign n4245 = n460 | n500 ;
  assign n4246 = n767 | n4245 ;
  assign n4247 = n4244 | n4246 ;
  assign n4248 = n4243 | n4247 ;
  assign n4249 = n220 | n245 ;
  assign n4250 = n1091 | n2423 ;
  assign n4251 = n4249 | n4250 ;
  assign n4252 = n2156 | n4251 ;
  assign n4253 = n4248 | n4252 ;
  assign n4254 = n204 | n666 ;
  assign n4255 = n139 | n190 ;
  assign n4256 = n3522 | n4255 ;
  assign n4257 = n4254 | n4256 ;
  assign n4258 = n317 | n4257 ;
  assign n4259 = n159 | n452 ;
  assign n4260 = n554 | n4259 ;
  assign n4261 = n407 | n839 ;
  assign n4262 = n1982 | n4261 ;
  assign n4263 = n4260 | n4262 ;
  assign n4264 = n2884 | n4263 ;
  assign n4265 = n4258 | n4264 ;
  assign n4266 = n489 | n594 ;
  assign n4267 = n1582 | n2427 ;
  assign n4268 = n4266 | n4267 ;
  assign n4269 = n811 | n2685 ;
  assign n4270 = n2524 | n4269 ;
  assign n4271 = n4268 | n4270 ;
  assign n4272 = n1758 | n3087 ;
  assign n4273 = n195 | n610 ;
  assign n4274 = n233 | n516 ;
  assign n4275 = n4273 | n4274 ;
  assign n4276 = n4272 | n4275 ;
  assign n4277 = n4271 | n4276 ;
  assign n4278 = n4265 | n4277 ;
  assign n4279 = n4253 | n4278 ;
  assign n4280 = n30119 & n2331 ;
  assign n30301 = ~n4279 ;
  assign n4281 = n30301 & n4280 ;
  assign n30302 = ~n4281 ;
  assign n4282 = x2 & n30302 ;
  assign n4283 = n30049 & n4281 ;
  assign n4284 = n195 | n1528 ;
  assign n4285 = n257 | n323 ;
  assign n4286 = n331 | n925 ;
  assign n4287 = n4285 | n4286 ;
  assign n4288 = n4284 | n4287 ;
  assign n4289 = n187 | n767 ;
  assign n4290 = n816 | n4289 ;
  assign n4291 = n2532 | n4290 ;
  assign n4292 = n2653 | n4291 ;
  assign n4293 = n4288 | n4292 ;
  assign n4294 = n116 | n232 ;
  assign n4295 = n1483 | n4294 ;
  assign n4296 = n3042 | n4295 ;
  assign n4297 = n204 | n849 ;
  assign n4298 = n4056 | n4297 ;
  assign n4299 = n957 | n1100 ;
  assign n4300 = n4298 | n4299 ;
  assign n4301 = n4296 | n4300 ;
  assign n4302 = n354 | n434 ;
  assign n4303 = n550 | n651 ;
  assign n4304 = n3948 | n4303 ;
  assign n4305 = n4302 | n4304 ;
  assign n4306 = n3905 | n4305 ;
  assign n4307 = n269 | n469 ;
  assign n4308 = n532 | n684 ;
  assign n4309 = n4307 | n4308 ;
  assign n4310 = n258 | n349 ;
  assign n4311 = n1249 | n4310 ;
  assign n4312 = n4309 | n4311 ;
  assign n4313 = n1267 | n1831 ;
  assign n4314 = n4312 | n4313 ;
  assign n4315 = n4306 | n4314 ;
  assign n4316 = n4301 | n4315 ;
  assign n4317 = n4293 | n4316 ;
  assign n4318 = n3935 | n4317 ;
  assign n4319 = n2599 | n4318 ;
  assign n4320 = x2 & n4319 ;
  assign n4321 = x2 | n4319 ;
  assign n4322 = n331 | n534 ;
  assign n4323 = n651 | n1199 ;
  assign n4324 = n4322 | n4323 ;
  assign n4325 = n2570 | n4324 ;
  assign n4326 = n3082 | n3966 ;
  assign n4327 = n4325 | n4326 ;
  assign n4328 = n141 | n242 ;
  assign n4329 = n1468 | n3538 ;
  assign n4330 = n4328 | n4329 ;
  assign n4331 = n1759 | n4330 ;
  assign n4332 = n4327 | n4331 ;
  assign n4333 = n3237 | n4332 ;
  assign n4334 = n910 | n3488 ;
  assign n4335 = n768 | n2558 ;
  assign n4336 = n4255 | n4302 ;
  assign n4337 = n4335 | n4336 ;
  assign n4338 = n861 | n4337 ;
  assign n4339 = n4334 | n4338 ;
  assign n4340 = n428 | n684 ;
  assign n4341 = n158 | n797 ;
  assign n4342 = n2732 | n4341 ;
  assign n4343 = n4340 | n4342 ;
  assign n4344 = n288 | n4343 ;
  assign n4345 = n4339 | n4344 ;
  assign n4346 = n2485 | n4345 ;
  assign n4347 = n4333 | n4346 ;
  assign n4348 = n1173 | n4347 ;
  assign n4349 = x2 & n4348 ;
  assign n4350 = x2 | n4348 ;
  assign n3349 = n2102 & n3343 ;
  assign n4357 = n2295 & n3311 ;
  assign n4358 = n2216 & n3329 ;
  assign n4359 = n4357 | n4358 ;
  assign n4360 = n3349 | n4359 ;
  assign n2809 = n2223 & n2808 ;
  assign n4351 = n2223 | n2808 ;
  assign n30303 = ~n2809 ;
  assign n4352 = n30303 & n4351 ;
  assign n4361 = n889 & n4352 ;
  assign n4362 = n4360 | n4361 ;
  assign n4363 = n4350 & n4362 ;
  assign n4364 = n4349 | n4363 ;
  assign n4365 = n4321 & n4364 ;
  assign n4366 = n4320 | n4365 ;
  assign n30304 = ~n4283 ;
  assign n4367 = n30304 & n4366 ;
  assign n4368 = n4282 | n4367 ;
  assign n4369 = n30223 & n3479 ;
  assign n30305 = ~n3586 ;
  assign n4370 = n30305 & n4369 ;
  assign n30306 = ~n4369 ;
  assign n4371 = n3586 & n30306 ;
  assign n4372 = n4370 | n4371 ;
  assign n4374 = n4368 & n4372 ;
  assign n4373 = n4368 | n4372 ;
  assign n30307 = ~n4374 ;
  assign n4375 = n4373 & n30307 ;
  assign n30308 = ~n2816 ;
  assign n3302 = n1966 & n30308 ;
  assign n30309 = ~n1966 ;
  assign n4376 = n30309 & n2816 ;
  assign n4377 = n3302 | n4376 ;
  assign n30310 = ~n4377 ;
  assign n4378 = n889 & n30310 ;
  assign n3319 = n30123 & n3311 ;
  assign n3340 = n30114 & n3329 ;
  assign n4383 = n3319 | n3340 ;
  assign n4384 = n30108 & n3343 ;
  assign n4385 = n4383 | n4384 ;
  assign n4386 = n4378 | n4385 ;
  assign n4388 = n4375 & n4386 ;
  assign n4389 = n4374 | n4388 ;
  assign n4390 = n3589 | n3590 ;
  assign n4391 = n3599 | n4390 ;
  assign n4392 = n3599 & n4390 ;
  assign n30311 = ~n4392 ;
  assign n4393 = n4391 & n30311 ;
  assign n30312 = ~n4389 ;
  assign n4394 = n30312 & n4393 ;
  assign n3309 = n895 & n3307 ;
  assign n1558 = n894 & n1556 ;
  assign n2870 = n30105 & n2861 ;
  assign n4395 = n1558 | n2870 ;
  assign n4396 = n30196 & n2849 ;
  assign n4397 = n4395 | n4396 ;
  assign n4398 = n3309 | n4397 ;
  assign n30313 = ~n4398 ;
  assign n4399 = x29 & n30313 ;
  assign n4400 = n30024 & n4398 ;
  assign n4401 = n4399 | n4400 ;
  assign n30314 = ~n4393 ;
  assign n4402 = n4389 & n30314 ;
  assign n4403 = n4394 | n4402 ;
  assign n4404 = n4401 | n4403 ;
  assign n30315 = ~n4394 ;
  assign n4405 = n30315 & n4404 ;
  assign n4406 = n4228 & n4239 ;
  assign n30316 = ~n4406 ;
  assign n4407 = n4240 & n30316 ;
  assign n30317 = ~n4405 ;
  assign n4408 = n30317 & n4407 ;
  assign n30318 = ~n4408 ;
  assign n4409 = n4240 & n30318 ;
  assign n4411 = n4224 | n4409 ;
  assign n30319 = ~n3616 ;
  assign n3617 = n3607 & n30319 ;
  assign n30320 = ~n3607 ;
  assign n4412 = n30320 & n3616 ;
  assign n4413 = n3617 | n4412 ;
  assign n4410 = n4224 & n4409 ;
  assign n30321 = ~n4410 ;
  assign n4414 = n30321 & n4411 ;
  assign n30322 = ~n4413 ;
  assign n4415 = n30322 & n4414 ;
  assign n30323 = ~n4415 ;
  assign n4416 = n4411 & n30323 ;
  assign n4418 = n4217 | n4416 ;
  assign n3782 = n3778 & n3781 ;
  assign n4419 = n3778 | n3781 ;
  assign n30324 = ~n3782 ;
  assign n4420 = n30324 & n4419 ;
  assign n4421 = n3791 & n4420 ;
  assign n3813 = n1074 & n3802 ;
  assign n3831 = n3764 & n3818 ;
  assign n4426 = n3813 | n3831 ;
  assign n4427 = n209 & n30074 ;
  assign n4428 = n4426 | n4427 ;
  assign n4429 = n4421 | n4428 ;
  assign n30325 = ~n4429 ;
  assign n4430 = x26 & n30325 ;
  assign n4431 = n30019 & n4429 ;
  assign n4432 = n4430 | n4431 ;
  assign n4417 = n4217 & n4416 ;
  assign n30326 = ~n4417 ;
  assign n4433 = n30326 & n4418 ;
  assign n30327 = ~n4432 ;
  assign n4434 = n30327 & n4433 ;
  assign n30328 = ~n4434 ;
  assign n4435 = n4418 & n30328 ;
  assign n4437 = n4215 | n4435 ;
  assign n30329 = ~n4033 ;
  assign n4116 = n30329 & n4114 ;
  assign n30330 = ~n4114 ;
  assign n4438 = n4033 & n30330 ;
  assign n4439 = n4116 | n4438 ;
  assign n4440 = n4093 & n4439 ;
  assign n4441 = n4093 | n4439 ;
  assign n30331 = ~n4440 ;
  assign n4442 = n30331 & n4441 ;
  assign n4443 = n4135 & n4442 ;
  assign n4158 = n4093 & n4148 ;
  assign n4179 = n4033 & n4165 ;
  assign n4448 = n4158 | n4179 ;
  assign n4449 = n30264 & n4185 ;
  assign n4450 = n4448 | n4449 ;
  assign n4451 = n4443 | n4450 ;
  assign n30332 = ~n4451 ;
  assign n4452 = x23 & n30332 ;
  assign n4453 = n30030 & n4451 ;
  assign n4454 = n4452 | n4453 ;
  assign n4436 = n4215 & n4435 ;
  assign n30333 = ~n4436 ;
  assign n4455 = n30333 & n4437 ;
  assign n30334 = ~n4454 ;
  assign n4456 = n30334 & n4455 ;
  assign n30335 = ~n4456 ;
  assign n4457 = n4437 & n30335 ;
  assign n4458 = n4213 & n4457 ;
  assign n4459 = n4213 | n4457 ;
  assign n30336 = ~n4458 ;
  assign n4460 = n30336 & n4459 ;
  assign n30337 = ~n4455 ;
  assign n4461 = n4454 & n30337 ;
  assign n4462 = n4456 | n4461 ;
  assign n30338 = ~n4433 ;
  assign n4463 = n4432 & n30338 ;
  assign n4464 = n4434 | n4463 ;
  assign n30339 = ~n4414 ;
  assign n4465 = n4413 & n30339 ;
  assign n4466 = n4415 | n4465 ;
  assign n3797 = n30173 & n3791 ;
  assign n1221 = n209 & n1219 ;
  assign n3825 = n1074 & n3818 ;
  assign n4467 = n1221 | n3825 ;
  assign n4468 = n30074 & n3802 ;
  assign n4469 = n4467 | n4468 ;
  assign n4470 = n3797 | n4469 ;
  assign n4471 = x26 | n4470 ;
  assign n4472 = x26 & n4470 ;
  assign n30340 = ~n4472 ;
  assign n4473 = n4471 & n30340 ;
  assign n4475 = n4466 & n4473 ;
  assign n30341 = ~n4466 ;
  assign n4474 = n30341 & n4473 ;
  assign n30342 = ~n4473 ;
  assign n4476 = n4466 & n30342 ;
  assign n4477 = n4474 | n4476 ;
  assign n30343 = ~n4407 ;
  assign n4478 = n4405 & n30343 ;
  assign n4479 = n4408 | n4478 ;
  assign n3386 = n895 & n30209 ;
  assign n1449 = n894 & n1445 ;
  assign n2858 = n1556 & n2849 ;
  assign n4480 = n1449 | n2858 ;
  assign n4481 = n30196 & n2861 ;
  assign n4482 = n4480 | n4481 ;
  assign n4483 = n3386 | n4482 ;
  assign n4484 = x29 | n4483 ;
  assign n4485 = x29 & n4483 ;
  assign n30344 = ~n4485 ;
  assign n4486 = n4484 & n30344 ;
  assign n4488 = n4479 & n4486 ;
  assign n3793 = n30212 & n3791 ;
  assign n3811 = n1219 & n3802 ;
  assign n3827 = n30074 & n3818 ;
  assign n4489 = n3811 | n3827 ;
  assign n4490 = n209 & n30082 ;
  assign n4491 = n4489 | n4490 ;
  assign n4492 = n3793 | n4491 ;
  assign n30345 = ~n4492 ;
  assign n4493 = x26 & n30345 ;
  assign n4494 = n30019 & n4492 ;
  assign n4495 = n4493 | n4494 ;
  assign n30346 = ~n4479 ;
  assign n4487 = n30346 & n4486 ;
  assign n30347 = ~n4486 ;
  assign n4496 = n4479 & n30347 ;
  assign n4497 = n4487 | n4496 ;
  assign n4499 = n4495 & n4497 ;
  assign n4500 = n4488 | n4499 ;
  assign n4502 = n4477 & n4500 ;
  assign n4503 = n4475 | n4502 ;
  assign n4504 = n4464 | n4503 ;
  assign n4505 = n4110 & n4112 ;
  assign n30348 = ~n4505 ;
  assign n4506 = n4113 & n30348 ;
  assign n30349 = ~n4506 ;
  assign n4508 = n4135 & n30349 ;
  assign n4170 = n4093 & n4165 ;
  assign n4197 = n3700 & n4185 ;
  assign n4512 = n4170 | n4197 ;
  assign n4513 = n30264 & n4148 ;
  assign n4514 = n4512 | n4513 ;
  assign n4515 = n4508 | n4514 ;
  assign n30350 = ~n4515 ;
  assign n4516 = x23 & n30350 ;
  assign n4517 = n30030 & n4515 ;
  assign n4518 = n4516 | n4517 ;
  assign n4519 = n4464 & n4503 ;
  assign n30351 = ~n4519 ;
  assign n4520 = n4504 & n30351 ;
  assign n30352 = ~n4518 ;
  assign n4521 = n30352 & n4520 ;
  assign n30353 = ~n4521 ;
  assign n4522 = n4504 & n30353 ;
  assign n4524 = n4462 | n4522 ;
  assign n4525 = n150 | n203 ;
  assign n4526 = n279 | n1010 ;
  assign n30354 = ~n235 ;
  assign n4527 = n145 & n30354 ;
  assign n30355 = ~n4526 ;
  assign n4528 = n30355 & n4527 ;
  assign n4529 = n94 & n2447 ;
  assign n30356 = ~n4529 ;
  assign n4530 = n4528 & n30356 ;
  assign n30357 = ~n4525 ;
  assign n4531 = n30357 & n4530 ;
  assign n30358 = ~n2362 ;
  assign n4532 = n30358 & n4531 ;
  assign n4533 = n568 | n839 ;
  assign n4534 = n572 | n4533 ;
  assign n4535 = n699 | n1141 ;
  assign n4536 = n4534 | n4535 ;
  assign n4537 = n815 | n858 ;
  assign n4538 = n337 | n608 ;
  assign n4539 = n2014 | n4538 ;
  assign n4540 = n4537 | n4539 ;
  assign n4541 = n130 | n220 ;
  assign n4542 = n461 | n4541 ;
  assign n4543 = n523 | n4542 ;
  assign n4544 = n4540 | n4543 ;
  assign n4545 = n1741 | n3561 ;
  assign n4546 = n4544 | n4545 ;
  assign n4547 = n4536 | n4546 ;
  assign n30359 = ~n4547 ;
  assign n4548 = n4532 & n30359 ;
  assign n4549 = n139 | n348 ;
  assign n4550 = n486 | n573 ;
  assign n4551 = n4549 | n4550 ;
  assign n4552 = n478 | n637 ;
  assign n4553 = n4551 | n4552 ;
  assign n4554 = n2147 | n2763 ;
  assign n4555 = n4553 | n4554 ;
  assign n4556 = n349 | n721 ;
  assign n4557 = n380 | n1415 ;
  assign n4558 = n4556 | n4557 ;
  assign n4559 = n1294 | n2451 ;
  assign n4560 = n3921 | n4559 ;
  assign n4561 = n4558 | n4560 ;
  assign n4562 = n4555 | n4561 ;
  assign n4563 = n3558 | n4562 ;
  assign n4564 = n3045 | n4563 ;
  assign n30360 = ~n4564 ;
  assign n4565 = n4548 & n30360 ;
  assign n4581 = n3938 & n4565 ;
  assign n30361 = ~n4565 ;
  assign n4570 = n3938 & n30361 ;
  assign n4582 = n30282 & n4565 ;
  assign n4583 = n4570 | n4582 ;
  assign n4120 = n3938 & n30281 ;
  assign n30362 = ~n4120 ;
  assign n4584 = n4117 & n30362 ;
  assign n30363 = ~n4584 ;
  assign n4586 = n4583 & n30363 ;
  assign n4587 = n4581 | n4586 ;
  assign n4588 = n139 | n277 ;
  assign n4589 = n359 | n448 ;
  assign n4590 = n4588 | n4589 ;
  assign n4591 = n176 | n323 ;
  assign n4592 = n1917 | n2014 ;
  assign n4593 = n4591 | n4592 ;
  assign n4594 = n4590 | n4593 ;
  assign n4595 = n2110 | n2624 ;
  assign n4596 = n318 | n1199 ;
  assign n4597 = n377 | n501 ;
  assign n4598 = n4596 | n4597 ;
  assign n4599 = n4595 | n4598 ;
  assign n4600 = n823 | n1132 ;
  assign n4601 = n1940 | n4600 ;
  assign n4602 = n1922 | n3922 ;
  assign n4603 = n3683 | n4602 ;
  assign n4604 = n4601 | n4603 ;
  assign n4605 = n4599 | n4604 ;
  assign n4606 = n4594 | n4605 ;
  assign n4607 = n4044 | n4606 ;
  assign n4608 = n3753 | n4286 ;
  assign n4609 = n433 | n491 ;
  assign n4610 = n845 | n4609 ;
  assign n4611 = n203 | n216 ;
  assign n4612 = n1943 | n4611 ;
  assign n4613 = n4610 | n4612 ;
  assign n4614 = n519 | n4613 ;
  assign n4615 = n4608 | n4614 ;
  assign n4616 = n4607 | n4615 ;
  assign n4617 = n1468 | n2282 ;
  assign n4618 = n327 | n512 ;
  assign n4619 = n3131 | n4618 ;
  assign n4620 = n4617 | n4619 ;
  assign n4621 = n488 | n827 ;
  assign n4622 = n2974 | n4621 ;
  assign n4623 = n4620 | n4622 ;
  assign n4624 = n133 | n446 ;
  assign n4625 = n1853 | n4624 ;
  assign n4626 = n2937 | n4625 ;
  assign n4627 = n4623 | n4626 ;
  assign n4628 = n416 | n528 ;
  assign n4629 = n972 | n1129 ;
  assign n4630 = n309 | n687 ;
  assign n4631 = n2030 | n4630 ;
  assign n4632 = n4629 | n4631 ;
  assign n4633 = n4628 | n4632 ;
  assign n4634 = n3062 | n4269 ;
  assign n4635 = n258 | n381 ;
  assign n4636 = n233 | n241 ;
  assign n4637 = n4635 | n4636 ;
  assign n4638 = n4634 | n4637 ;
  assign n4639 = n4633 | n4638 ;
  assign n4640 = n4627 | n4639 ;
  assign n4641 = n138 | n257 ;
  assign n4642 = n587 | n4641 ;
  assign n4643 = n1513 | n3568 ;
  assign n4644 = n4642 | n4643 ;
  assign n4645 = n302 | n337 ;
  assign n4646 = n383 | n4645 ;
  assign n4647 = n809 | n4646 ;
  assign n4648 = n4644 | n4647 ;
  assign n4649 = n1759 | n4648 ;
  assign n4650 = n283 | n470 ;
  assign n4651 = n116 | n185 ;
  assign n4652 = n224 | n369 ;
  assign n4653 = n384 | n4652 ;
  assign n4654 = n4651 | n4653 ;
  assign n4655 = n4650 | n4654 ;
  assign n4656 = n1389 | n3153 ;
  assign n4657 = n520 | n568 ;
  assign n4658 = n1099 | n4657 ;
  assign n4659 = n3961 | n4658 ;
  assign n4660 = n4656 | n4659 ;
  assign n4661 = n4655 | n4660 ;
  assign n4662 = n4649 | n4661 ;
  assign n4663 = n4640 | n4662 ;
  assign n4664 = n4616 | n4663 ;
  assign n4669 = n4565 | n4664 ;
  assign n4670 = n4565 & n4664 ;
  assign n30364 = ~n4670 ;
  assign n4671 = n4669 & n30364 ;
  assign n30365 = ~n4671 ;
  assign n4672 = n4587 & n30365 ;
  assign n30366 = ~n4587 ;
  assign n4673 = n30366 & n4671 ;
  assign n4674 = n4672 | n4673 ;
  assign n29892 = x17 & x18 ;
  assign n4680 = x17 | x18 ;
  assign n30367 = ~n29892 ;
  assign n4683 = n30367 & n4680 ;
  assign n37287 = x19 & x20 ;
  assign n4684 = x19 | x20 ;
  assign n30368 = ~n37287 ;
  assign n4685 = n30368 & n4684 ;
  assign n4686 = n4683 & n4685 ;
  assign n4688 = n4674 & n4686 ;
  assign n30369 = ~n4680 ;
  assign n4681 = x19 & n30369 ;
  assign n30370 = ~x19 ;
  assign n4705 = n30370 & n29892 ;
  assign n4706 = n4681 | n4705 ;
  assign n4715 = n30361 & n4706 ;
  assign n30371 = ~n4685 ;
  assign n4748 = n4683 & n30371 ;
  assign n4758 = n4664 & n4748 ;
  assign n4767 = n4715 | n4758 ;
  assign n4724 = n4683 | n4706 ;
  assign n30372 = ~n4724 ;
  assign n4726 = n4685 & n30372 ;
  assign n4768 = n30282 & n4726 ;
  assign n4769 = n4767 | n4768 ;
  assign n4770 = n4688 | n4769 ;
  assign n30373 = ~n4770 ;
  assign n4771 = x20 & n30373 ;
  assign n30374 = ~x20 ;
  assign n4772 = n30374 & n4770 ;
  assign n4773 = n4771 | n4772 ;
  assign n30375 = ~n4462 ;
  assign n4523 = n30375 & n4522 ;
  assign n30376 = ~n4522 ;
  assign n4774 = n4462 & n30376 ;
  assign n4775 = n4523 | n4774 ;
  assign n30377 = ~n4773 ;
  assign n4776 = n30377 & n4775 ;
  assign n30378 = ~n4776 ;
  assign n4777 = n4524 & n30378 ;
  assign n30379 = ~n4460 ;
  assign n4778 = n30379 & n4777 ;
  assign n30380 = ~n4777 ;
  assign n4779 = n4460 & n30380 ;
  assign n4780 = n4778 | n4779 ;
  assign n4781 = n326 | n1101 ;
  assign n4782 = n2176 | n4781 ;
  assign n4783 = n623 | n4782 ;
  assign n4784 = n703 | n1587 ;
  assign n4785 = n4783 | n4784 ;
  assign n4786 = n296 | n417 ;
  assign n4787 = n477 | n4786 ;
  assign n4788 = n653 | n4787 ;
  assign n4789 = n1902 | n4788 ;
  assign n4790 = n168 | n795 ;
  assign n4791 = n564 | n978 ;
  assign n4792 = n200 | n279 ;
  assign n4793 = n4791 | n4792 ;
  assign n4794 = n4790 | n4793 ;
  assign n4795 = n3451 | n4794 ;
  assign n4796 = n4789 | n4795 ;
  assign n4797 = n4253 | n4796 ;
  assign n4798 = n4785 | n4797 ;
  assign n4799 = n103 | n138 ;
  assign n4800 = n572 | n4799 ;
  assign n4801 = n234 | n4800 ;
  assign n4802 = n1361 | n1843 ;
  assign n4803 = n4801 | n4802 ;
  assign n4804 = n534 | n676 ;
  assign n4805 = n1129 | n1469 ;
  assign n4806 = n4804 | n4805 ;
  assign n4807 = n792 | n4806 ;
  assign n4808 = n1925 | n4807 ;
  assign n4809 = n4803 | n4808 ;
  assign n4810 = n1839 | n4809 ;
  assign n4811 = n4798 | n4810 ;
  assign n30381 = ~n4664 ;
  assign n4823 = n30381 & n4811 ;
  assign n30382 = ~n4811 ;
  assign n4831 = n4664 & n30382 ;
  assign n4832 = n4823 | n4831 ;
  assign n4833 = n4565 & n30381 ;
  assign n4834 = n4672 | n4833 ;
  assign n30383 = ~n4834 ;
  assign n4835 = n4832 & n30383 ;
  assign n30384 = ~n4832 ;
  assign n4836 = n30384 & n4834 ;
  assign n4837 = n4835 | n4836 ;
  assign n30385 = ~n4837 ;
  assign n4838 = n4686 & n30385 ;
  assign n4741 = n30361 & n4726 ;
  assign n4824 = n4748 & n4811 ;
  assign n4844 = n4741 | n4824 ;
  assign n4845 = n4664 & n4706 ;
  assign n4846 = n4844 | n4845 ;
  assign n4847 = n4838 | n4846 ;
  assign n30386 = ~n4847 ;
  assign n4848 = x20 & n30386 ;
  assign n4849 = n30374 & n4847 ;
  assign n4850 = n4848 | n4849 ;
  assign n30387 = ~n4850 ;
  assign n4851 = n4780 & n30387 ;
  assign n30388 = ~n4780 ;
  assign n4852 = n30388 & n4850 ;
  assign n4853 = n4851 | n4852 ;
  assign n4854 = n614 | n2951 ;
  assign n4855 = n1238 | n1361 ;
  assign n4856 = n4854 | n4855 ;
  assign n4857 = n433 | n451 ;
  assign n4858 = n2410 | n4857 ;
  assign n4859 = n636 | n676 ;
  assign n4860 = n338 | n660 ;
  assign n4861 = n4859 | n4860 ;
  assign n4862 = n4858 | n4861 ;
  assign n4863 = n272 | n277 ;
  assign n4864 = n418 | n4863 ;
  assign n4865 = n216 | n221 ;
  assign n4866 = n711 | n4865 ;
  assign n4867 = n4864 | n4866 ;
  assign n4868 = n4862 | n4867 ;
  assign n4869 = n4856 | n4868 ;
  assign n4870 = n585 | n3421 ;
  assign n4871 = n133 | n841 ;
  assign n4872 = n202 | n245 ;
  assign n4873 = n4871 | n4872 ;
  assign n4874 = n4870 | n4873 ;
  assign n4875 = n186 | n684 ;
  assign n4876 = n925 | n4875 ;
  assign n4877 = n3992 | n4876 ;
  assign n4878 = n4874 | n4877 ;
  assign n4879 = n924 | n3729 ;
  assign n4880 = n1633 | n4879 ;
  assign n4881 = n4878 | n4880 ;
  assign n4882 = n179 | n296 ;
  assign n4883 = n326 | n446 ;
  assign n4884 = n4882 | n4883 ;
  assign n4885 = n239 | n913 ;
  assign n4886 = n4884 | n4885 ;
  assign n4887 = n355 | n906 ;
  assign n4888 = n4886 | n4887 ;
  assign n4889 = n554 | n677 ;
  assign n4890 = n695 | n788 ;
  assign n4891 = n217 | n4890 ;
  assign n4892 = n4889 | n4891 ;
  assign n4893 = n4888 | n4892 ;
  assign n4894 = n4881 | n4893 ;
  assign n4895 = n4869 | n4894 ;
  assign n4896 = n630 | n2500 ;
  assign n4897 = n811 | n4896 ;
  assign n4898 = n469 | n487 ;
  assign n4899 = n795 | n4898 ;
  assign n4900 = n2046 | n4899 ;
  assign n4901 = n2175 | n2458 ;
  assign n4902 = n4900 | n4901 ;
  assign n4903 = n4897 | n4902 ;
  assign n4904 = n256 | n270 ;
  assign n3812 = x26 | n3802 ;
  assign n4905 = n86 & n3812 ;
  assign n4906 = n566 | n4905 ;
  assign n4907 = n4904 | n4906 ;
  assign n4908 = n513 | n611 ;
  assign n4909 = n930 | n1129 ;
  assign n4910 = n4908 | n4909 ;
  assign n4911 = n185 | n235 ;
  assign n4912 = n495 | n568 ;
  assign n4913 = n687 | n4912 ;
  assign n4914 = n4911 | n4913 ;
  assign n4915 = n4910 | n4914 ;
  assign n4916 = n532 | n1370 ;
  assign n30389 = ~n4916 ;
  assign n4917 = n145 & n30389 ;
  assign n4918 = n320 | n345 ;
  assign n4919 = n2477 | n3736 ;
  assign n4920 = n4918 | n4919 ;
  assign n30390 = ~n4920 ;
  assign n4921 = n4917 & n30390 ;
  assign n30391 = ~n4915 ;
  assign n4922 = n30391 & n4921 ;
  assign n30392 = ~n4907 ;
  assign n4923 = n30392 & n4922 ;
  assign n30393 = ~n4903 ;
  assign n4924 = n30393 & n4923 ;
  assign n30394 = ~n4895 ;
  assign n4925 = n30394 & n4924 ;
  assign n4943 = n509 | n622 ;
  assign n4944 = n434 | n4073 ;
  assign n4945 = n4943 | n4944 ;
  assign n4946 = n3655 | n4945 ;
  assign n4947 = n396 | n1129 ;
  assign n4948 = n601 | n4947 ;
  assign n4949 = n199 | n651 ;
  assign n4950 = n1572 | n4949 ;
  assign n4951 = n4948 | n4950 ;
  assign n4952 = n255 | n513 ;
  assign n4953 = n1311 | n1688 ;
  assign n4954 = n4952 | n4953 ;
  assign n4955 = n205 | n1787 ;
  assign n4956 = n365 | n489 ;
  assign n4957 = n925 | n1179 ;
  assign n4958 = n4956 | n4957 ;
  assign n4959 = n4955 | n4958 ;
  assign n4960 = n4954 | n4959 ;
  assign n4961 = n200 | n314 ;
  assign n4962 = n371 | n4961 ;
  assign n4963 = n245 | n349 ;
  assign n4964 = n453 | n1049 ;
  assign n4965 = n4963 | n4964 ;
  assign n4966 = n4962 | n4965 ;
  assign n4967 = n280 | n568 ;
  assign n4968 = n2584 | n3422 ;
  assign n4969 = n4967 | n4968 ;
  assign n4970 = n4966 | n4969 ;
  assign n4971 = n4960 | n4970 ;
  assign n4972 = n4951 | n4971 ;
  assign n4973 = n4946 | n4972 ;
  assign n4974 = n232 | n369 ;
  assign n4975 = n445 | n554 ;
  assign n4976 = n636 | n4975 ;
  assign n4977 = n4974 | n4976 ;
  assign n4978 = n270 | n290 ;
  assign n4979 = n1713 | n4978 ;
  assign n4980 = n4977 | n4979 ;
  assign n1484 = n283 | n310 ;
  assign n4981 = n379 | n1484 ;
  assign n4982 = n924 | n4981 ;
  assign n4983 = n3129 | n4982 ;
  assign n4984 = n4980 | n4983 ;
  assign n4985 = n704 | n3753 ;
  assign n4986 = n223 | n857 ;
  assign n4987 = n163 | n474 ;
  assign n4988 = n4986 | n4987 ;
  assign n4989 = n1286 | n4988 ;
  assign n4990 = n4985 | n4989 ;
  assign n4991 = n2721 | n4990 ;
  assign n4992 = n4984 | n4991 ;
  assign n4993 = n4973 | n4992 ;
  assign n4994 = n529 | n594 ;
  assign n4995 = n833 | n4994 ;
  assign n4996 = n921 | n1193 ;
  assign n4997 = n80 | n497 ;
  assign n4998 = n2477 | n4997 ;
  assign n4999 = n4996 | n4998 ;
  assign n5000 = n770 | n1662 ;
  assign n5001 = n460 | n659 ;
  assign n5002 = n5000 | n5001 ;
  assign n5003 = n4999 | n5002 ;
  assign n5004 = n4995 | n5003 ;
  assign n5005 = n500 | n1497 ;
  assign n30395 = ~n2441 ;
  assign n5006 = n82 & n30395 ;
  assign n5007 = n2456 | n5006 ;
  assign n5008 = n5005 | n5007 ;
  assign n5009 = n1279 | n5008 ;
  assign n5010 = n97 | n133 ;
  assign n5011 = n452 | n5010 ;
  assign n5012 = n4860 | n5011 ;
  assign n5013 = n196 | n3093 ;
  assign n5014 = n5012 | n5013 ;
  assign n5015 = n5009 | n5014 ;
  assign n5016 = n5004 | n5015 ;
  assign n5017 = n4993 | n5016 ;
  assign n5025 = n4925 | n5017 ;
  assign n5026 = n4925 & n5017 ;
  assign n30396 = ~n5026 ;
  assign n5027 = n5025 & n30396 ;
  assign n5028 = n344 | n549 ;
  assign n5029 = n921 | n5028 ;
  assign n5030 = n410 | n816 ;
  assign n5031 = n239 | n5030 ;
  assign n5032 = n2717 | n5031 ;
  assign n5033 = n319 | n324 ;
  assign n5034 = n313 | n477 ;
  assign n5035 = n5033 | n5034 ;
  assign n5036 = n1051 | n3922 ;
  assign n5037 = n5035 | n5036 ;
  assign n5038 = n5032 | n5037 ;
  assign n5039 = n5029 | n5038 ;
  assign n5040 = n300 | n4244 ;
  assign n5041 = n564 | n608 ;
  assign n5042 = n767 | n1787 ;
  assign n5043 = n5041 | n5042 ;
  assign n5044 = n1532 | n5043 ;
  assign n5045 = n5040 | n5044 ;
  assign n30397 = ~n174 ;
  assign n5046 = n145 & n30397 ;
  assign n30398 = ~n401 ;
  assign n5047 = n30398 & n5046 ;
  assign n5048 = n1286 | n1618 ;
  assign n30399 = ~n5048 ;
  assign n5049 = n5047 & n30399 ;
  assign n30400 = ~n5045 ;
  assign n5050 = n30400 & n5049 ;
  assign n30401 = ~n5039 ;
  assign n5051 = n30401 & n5050 ;
  assign n5052 = n167 | n566 ;
  assign n5053 = n355 | n470 ;
  assign n5054 = n602 | n833 ;
  assign n5055 = n2748 | n5054 ;
  assign n5056 = n5053 | n5055 ;
  assign n5057 = n5052 | n5056 ;
  assign n5058 = n513 | n865 ;
  assign n5059 = n3738 | n5058 ;
  assign n5060 = n696 | n1688 ;
  assign n5061 = n369 | n439 ;
  assign n5062 = n689 | n5061 ;
  assign n5063 = n5060 | n5062 ;
  assign n5064 = n5059 | n5063 ;
  assign n5065 = n150 | n1495 ;
  assign n5066 = n809 | n5065 ;
  assign n5067 = n916 | n962 ;
  assign n5068 = n5066 | n5067 ;
  assign n5069 = n223 | n1967 ;
  assign n5070 = n4949 | n5069 ;
  assign n5071 = n289 | n418 ;
  assign n5072 = n279 | n534 ;
  assign n5073 = n176 | n520 ;
  assign n5074 = n5072 | n5073 ;
  assign n5075 = n5071 | n5074 ;
  assign n5076 = n5070 | n5075 ;
  assign n5077 = n5068 | n5076 ;
  assign n5078 = n5064 | n5077 ;
  assign n5079 = n5057 | n5078 ;
  assign n30402 = ~n5079 ;
  assign n5080 = n5051 & n30402 ;
  assign n5081 = n1879 | n3729 ;
  assign n5082 = n248 | n2954 ;
  assign n5083 = n4020 | n5082 ;
  assign n5084 = n5081 | n5083 ;
  assign n5085 = n151 | n380 ;
  assign n5086 = n2477 | n3128 ;
  assign n5087 = n5085 | n5086 ;
  assign n5088 = n240 | n460 ;
  assign n5089 = n487 | n610 ;
  assign n5090 = n5088 | n5089 ;
  assign n5091 = n113 | n846 ;
  assign n5092 = n5090 | n5091 ;
  assign n5093 = n5087 | n5092 ;
  assign n5094 = n186 | n214 ;
  assign n5095 = n2681 | n5094 ;
  assign n5096 = n448 | n676 ;
  assign n5097 = n4086 | n5096 ;
  assign n5098 = n5095 | n5097 ;
  assign n5099 = n312 | n946 ;
  assign n5100 = n4261 | n5099 ;
  assign n5101 = n5098 | n5100 ;
  assign n5102 = n5093 | n5101 ;
  assign n5103 = n5084 | n5102 ;
  assign n5104 = n3487 | n5103 ;
  assign n30403 = ~n5104 ;
  assign n5105 = n5080 & n30403 ;
  assign n30404 = ~n5017 ;
  assign n5120 = n30404 & n5105 ;
  assign n30405 = ~n5105 ;
  assign n5122 = n5017 & n30405 ;
  assign n5123 = n5120 | n5122 ;
  assign n5121 = n30382 & n5105 ;
  assign n5124 = n4811 & n30405 ;
  assign n5125 = n5121 | n5124 ;
  assign n5126 = n4664 | n4811 ;
  assign n5127 = n4832 & n4834 ;
  assign n30406 = ~n5127 ;
  assign n5128 = n5126 & n30406 ;
  assign n5129 = n5125 | n5128 ;
  assign n30407 = ~n5121 ;
  assign n5130 = n30407 & n5129 ;
  assign n5132 = n5123 | n5130 ;
  assign n30408 = ~n5120 ;
  assign n5133 = n30408 & n5132 ;
  assign n5134 = n5027 | n5133 ;
  assign n5135 = n5027 & n5133 ;
  assign n30409 = ~n5135 ;
  assign n5136 = n5134 & n30409 ;
  assign n30410 = ~n5136 ;
  assign n5137 = n37300 & n30410 ;
  assign n30411 = ~n37294 ;
  assign n37295 = x16 & n30411 ;
  assign n30412 = ~x16 ;
  assign n5143 = n30412 & n29877 ;
  assign n5144 = n37295 | n5143 ;
  assign n5164 = n37297 | n5144 ;
  assign n30413 = ~n5164 ;
  assign n5166 = n37299 & n30413 ;
  assign n5179 = n30405 & n5166 ;
  assign n30414 = ~n37299 ;
  assign n5191 = n37297 & n30414 ;
  assign n30415 = ~n4925 ;
  assign n5204 = n30415 & n5191 ;
  assign n5213 = n5179 | n5204 ;
  assign n5214 = n5017 & n5144 ;
  assign n5215 = n5213 | n5214 ;
  assign n5216 = n5137 | n5215 ;
  assign n5217 = x17 | n5216 ;
  assign n5218 = x17 & n5216 ;
  assign n30416 = ~n5218 ;
  assign n5219 = n5217 & n30416 ;
  assign n30417 = ~n4853 ;
  assign n5220 = n30417 & n5219 ;
  assign n30418 = ~n5219 ;
  assign n5221 = n4853 & n30418 ;
  assign n5222 = n5220 | n5221 ;
  assign n30419 = ~n4775 ;
  assign n5223 = n4773 & n30419 ;
  assign n5224 = n4776 | n5223 ;
  assign n30420 = ~n4520 ;
  assign n5225 = n4518 & n30420 ;
  assign n5226 = n4521 | n5225 ;
  assign n30421 = ~n4500 ;
  assign n4501 = n4477 & n30421 ;
  assign n30422 = ~n4477 ;
  assign n5227 = n30422 & n4500 ;
  assign n5228 = n4501 | n5227 ;
  assign n4137 = n30263 & n4135 ;
  assign n4153 = n3700 & n4148 ;
  assign n4186 = n3764 & n4185 ;
  assign n5229 = n4153 | n4186 ;
  assign n5230 = n30264 & n4165 ;
  assign n5231 = n5229 | n5230 ;
  assign n5232 = n4137 | n5231 ;
  assign n5233 = x23 | n5232 ;
  assign n5234 = x23 & n5232 ;
  assign n30423 = ~n5234 ;
  assign n5235 = n5233 & n30423 ;
  assign n5237 = n5228 | n5235 ;
  assign n30424 = ~n5228 ;
  assign n5236 = n30424 & n5235 ;
  assign n30425 = ~n5235 ;
  assign n5238 = n5228 & n30425 ;
  assign n5239 = n5236 | n5238 ;
  assign n30426 = ~n4495 ;
  assign n4498 = n30426 & n4497 ;
  assign n30427 = ~n4497 ;
  assign n5240 = n4495 & n30427 ;
  assign n5241 = n4498 | n5240 ;
  assign n5242 = n4401 & n4403 ;
  assign n30428 = ~n5242 ;
  assign n5243 = n4404 & n30428 ;
  assign n30429 = ~n4386 ;
  assign n4387 = n4375 & n30429 ;
  assign n30430 = ~n4375 ;
  assign n5244 = n30430 & n4386 ;
  assign n5245 = n4387 | n5244 ;
  assign n5246 = n4282 | n4283 ;
  assign n30431 = ~n5246 ;
  assign n5247 = n4366 & n30431 ;
  assign n30432 = ~n4366 ;
  assign n5248 = n30432 & n5246 ;
  assign n5249 = n5247 | n5248 ;
  assign n2814 = n2065 & n2813 ;
  assign n5250 = n2065 | n2813 ;
  assign n30433 = ~n2814 ;
  assign n5251 = n30433 & n5250 ;
  assign n5252 = n889 & n5251 ;
  assign n3332 = n30123 & n3329 ;
  assign n3351 = n30114 & n3343 ;
  assign n5258 = n3332 | n3351 ;
  assign n5259 = n2102 & n3311 ;
  assign n5260 = n5258 | n5259 ;
  assign n5261 = n5252 | n5260 ;
  assign n30434 = ~n5249 ;
  assign n5263 = n30434 & n5261 ;
  assign n30435 = ~n4320 ;
  assign n5264 = n30435 & n4321 ;
  assign n30436 = ~n4364 ;
  assign n5265 = n30436 & n5264 ;
  assign n30437 = ~n5264 ;
  assign n5266 = n4364 & n30437 ;
  assign n5267 = n5265 | n5266 ;
  assign n30438 = ~n2109 ;
  assign n3301 = n30438 & n2811 ;
  assign n30439 = ~n2811 ;
  assign n5268 = n2109 & n30439 ;
  assign n5269 = n3301 | n5268 ;
  assign n30440 = ~n5269 ;
  assign n5271 = n889 & n30440 ;
  assign n3317 = n2216 & n3311 ;
  assign n3335 = n2102 & n3329 ;
  assign n5276 = n3317 | n3335 ;
  assign n5277 = n30123 & n3343 ;
  assign n5278 = n5276 | n5277 ;
  assign n5279 = n5271 | n5278 ;
  assign n5281 = n5267 & n5279 ;
  assign n5280 = n5267 | n5279 ;
  assign n30441 = ~n5281 ;
  assign n5282 = n5280 & n30441 ;
  assign n5283 = n112 | n658 ;
  assign n5284 = n239 | n5283 ;
  assign n5285 = n384 | n521 ;
  assign n5286 = n5284 | n5285 ;
  assign n5287 = n256 | n4294 ;
  assign n5288 = n5286 | n5287 ;
  assign n5289 = n216 | n289 ;
  assign n5290 = n318 | n961 ;
  assign n5291 = n5289 | n5290 ;
  assign n5292 = n3754 | n5291 ;
  assign n5293 = n642 | n683 ;
  assign n5294 = n202 | n469 ;
  assign n5295 = n696 | n5294 ;
  assign n5296 = n5293 | n5295 ;
  assign n5297 = n2583 | n5296 ;
  assign n5298 = n5292 | n5297 ;
  assign n5299 = n5288 | n5298 ;
  assign n5300 = n1723 | n5299 ;
  assign n5301 = n429 | n858 ;
  assign n5302 = n162 | n249 ;
  assign n5303 = n973 | n5302 ;
  assign n5304 = n1101 | n3118 ;
  assign n5305 = n5303 | n5304 ;
  assign n5306 = n425 | n5305 ;
  assign n5307 = n5301 | n5306 ;
  assign n5308 = n273 | n407 ;
  assign n5309 = n568 | n1787 ;
  assign n5310 = n5308 | n5309 ;
  assign n5311 = n2974 | n5310 ;
  assign n1353 = n199 | n360 ;
  assign n5312 = n1353 | n3729 ;
  assign n5313 = n5311 | n5312 ;
  assign n5314 = n3172 | n5313 ;
  assign n5315 = n5307 | n5314 ;
  assign n5316 = n713 | n3227 ;
  assign n5317 = n3547 | n5316 ;
  assign n5318 = n1366 | n4299 ;
  assign n5319 = n5317 | n5318 ;
  assign n5320 = n377 | n509 ;
  assign n5321 = n2650 | n5320 ;
  assign n5322 = n2677 | n3523 ;
  assign n5323 = n5321 | n5322 ;
  assign n5324 = n130 | n332 ;
  assign n5325 = n660 | n5324 ;
  assign n5326 = n3568 | n5325 ;
  assign n5327 = n294 | n1609 ;
  assign n5328 = n5326 | n5327 ;
  assign n5329 = n5323 | n5328 ;
  assign n5330 = n5319 | n5329 ;
  assign n5331 = n3500 | n5330 ;
  assign n5332 = n5315 | n5331 ;
  assign n5333 = n5300 | n5332 ;
  assign n30442 = ~n2805 ;
  assign n2806 = n2302 & n30442 ;
  assign n30443 = ~n2302 ;
  assign n5334 = n30443 & n2805 ;
  assign n5335 = n2806 | n5334 ;
  assign n30444 = ~n5335 ;
  assign n5336 = n889 & n30444 ;
  assign n3331 = n2295 & n3329 ;
  assign n3346 = n2216 & n3343 ;
  assign n5342 = n3331 | n3346 ;
  assign n30445 = ~n2376 ;
  assign n5343 = n30445 & n3311 ;
  assign n5344 = n5342 | n5343 ;
  assign n5345 = n5336 | n5344 ;
  assign n5346 = n5333 | n5345 ;
  assign n5347 = n5333 & n5345 ;
  assign n30446 = ~n5347 ;
  assign n5348 = n5346 & n30446 ;
  assign n5349 = n224 | n480 ;
  assign n5350 = n215 | n5349 ;
  assign n5351 = n1609 | n5350 ;
  assign n5352 = n3488 | n5060 ;
  assign n5353 = n5351 | n5352 ;
  assign n5354 = n90 | n793 ;
  assign n5355 = n2110 | n2611 ;
  assign n5356 = n5354 | n5355 ;
  assign n5357 = n533 | n609 ;
  assign n5358 = n1662 | n1859 ;
  assign n5359 = n5357 | n5358 ;
  assign n5360 = n5356 | n5359 ;
  assign n5361 = n232 | n300 ;
  assign n5362 = n333 | n5361 ;
  assign n5363 = n2458 | n5362 ;
  assign n5364 = n236 | n430 ;
  assign n5365 = n678 | n5364 ;
  assign n5366 = n5363 | n5365 ;
  assign n5367 = n5360 | n5366 ;
  assign n5368 = n5353 | n5367 ;
  assign n5369 = n2892 | n5368 ;
  assign n5370 = n553 | n841 ;
  assign n5371 = n900 | n5370 ;
  assign n5372 = n428 | n1513 ;
  assign n5373 = n3201 | n5372 ;
  assign n5374 = n314 | n344 ;
  assign n5375 = n1714 | n5374 ;
  assign n5376 = n5373 | n5375 ;
  assign n5377 = n5371 | n5376 ;
  assign n5378 = n241 | n978 ;
  assign n5379 = n687 | n865 ;
  assign n5380 = n788 | n5379 ;
  assign n5381 = n5378 | n5380 ;
  assign n5382 = n357 | n5381 ;
  assign n5383 = n2394 | n3023 ;
  assign n5384 = n277 | n666 ;
  assign n5385 = n1353 | n5384 ;
  assign n5386 = n5383 | n5385 ;
  assign n5387 = n5382 | n5386 ;
  assign n5388 = n5377 | n5387 ;
  assign n5389 = n3918 | n5388 ;
  assign n5390 = n5369 | n5389 ;
  assign n2803 = n2381 | n2802 ;
  assign n5391 = n2381 & n2802 ;
  assign n30447 = ~n5391 ;
  assign n5392 = n2803 & n30447 ;
  assign n5393 = n889 & n5392 ;
  assign n3318 = n30157 & n3311 ;
  assign n3348 = n2295 & n3343 ;
  assign n5399 = n3318 | n3348 ;
  assign n5400 = n30445 & n3329 ;
  assign n5401 = n5399 | n5400 ;
  assign n5402 = n5393 | n5401 ;
  assign n5403 = n5390 | n5402 ;
  assign n5404 = n5390 & n5402 ;
  assign n30448 = ~n5404 ;
  assign n5405 = n5403 & n30448 ;
  assign n5406 = n466 | n594 ;
  assign n5407 = n159 | n258 ;
  assign n5408 = n3201 | n5407 ;
  assign n5409 = n5406 | n5408 ;
  assign n5410 = n255 | n451 ;
  assign n5411 = n1996 | n5410 ;
  assign n5412 = n3493 | n5411 ;
  assign n5413 = n5409 | n5412 ;
  assign n5414 = n190 | n808 ;
  assign n5415 = n248 | n764 ;
  assign n5416 = n5414 | n5415 ;
  assign n5417 = n1371 | n4611 ;
  assign n5418 = n5416 | n5417 ;
  assign n5419 = n1183 | n5418 ;
  assign n5420 = n2247 | n5419 ;
  assign n5421 = n293 | n989 ;
  assign n5422 = n421 | n5421 ;
  assign n5423 = n4990 | n5422 ;
  assign n5424 = n5420 | n5423 ;
  assign n5425 = n5413 | n5424 ;
  assign n5426 = n1509 | n1880 ;
  assign n5427 = n5058 | n5426 ;
  assign n5428 = n756 | n1230 ;
  assign n5429 = n1323 | n2517 ;
  assign n5430 = n5428 | n5429 ;
  assign n5431 = n83 | n103 ;
  assign n5432 = n658 | n679 ;
  assign n5433 = n5431 | n5432 ;
  assign n5434 = n470 | n553 ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = n5430 | n5435 ;
  assign n5437 = n614 | n797 ;
  assign n5438 = n2687 | n5437 ;
  assign n5439 = n3096 | n5438 ;
  assign n5440 = n5436 | n5439 ;
  assign n5441 = n5427 | n5440 ;
  assign n30449 = ~n5441 ;
  assign n5442 = n3294 & n30449 ;
  assign n30450 = ~n5425 ;
  assign n5443 = n30450 & n5442 ;
  assign n5444 = n2376 | n2800 ;
  assign n30451 = ~n2801 ;
  assign n5445 = n30451 & n5444 ;
  assign n30452 = ~n5445 ;
  assign n5446 = n889 & n30452 ;
  assign n3334 = n30157 & n3329 ;
  assign n3350 = n30445 & n3343 ;
  assign n5452 = n3334 | n3350 ;
  assign n30453 = ~n2701 ;
  assign n5453 = n30453 & n3311 ;
  assign n5454 = n5452 | n5453 ;
  assign n5455 = n5446 | n5454 ;
  assign n30454 = ~n5455 ;
  assign n5456 = n5443 & n30454 ;
  assign n30455 = ~n5443 ;
  assign n5457 = n30455 & n5455 ;
  assign n5458 = n5456 | n5457 ;
  assign n5459 = n338 | n509 ;
  assign n5460 = n550 | n5459 ;
  assign n5461 = n107 | n174 ;
  assign n5462 = n4804 | n5461 ;
  assign n5463 = n5460 | n5462 ;
  assign n5464 = n566 | n1391 ;
  assign n5465 = n179 | n473 ;
  assign n5466 = n540 | n5465 ;
  assign n5467 = n2733 | n5466 ;
  assign n5468 = n5464 | n5467 ;
  assign n5469 = n5463 | n5468 ;
  assign n5470 = n1129 | n2659 ;
  assign n5471 = n4302 | n5470 ;
  assign n5472 = n245 | n380 ;
  assign n5473 = n448 | n512 ;
  assign n5474 = n5472 | n5473 ;
  assign n5475 = n126 | n808 ;
  assign n5476 = n946 | n5475 ;
  assign n5477 = n5474 | n5476 ;
  assign n5478 = n1041 | n1501 ;
  assign n5479 = n5477 | n5478 ;
  assign n5480 = n5471 | n5479 ;
  assign n5481 = n2628 | n3729 ;
  assign n5482 = n97 | n474 ;
  assign n5483 = n168 | n334 ;
  assign n5484 = n5482 | n5483 ;
  assign n5485 = n200 | n401 ;
  assign n5486 = n1249 | n5485 ;
  assign n5487 = n5484 | n5486 ;
  assign n5488 = n5481 | n5487 ;
  assign n5489 = n878 | n5488 ;
  assign n5490 = n5480 | n5489 ;
  assign n5491 = n5469 | n5490 ;
  assign n5492 = n2153 | n5491 ;
  assign n30456 = ~n2798 ;
  assign n5493 = n2702 & n30456 ;
  assign n5494 = n30157 & n5493 ;
  assign n30457 = ~n5493 ;
  assign n5495 = n2779 & n30457 ;
  assign n5496 = n5494 | n5495 ;
  assign n30458 = ~n5496 ;
  assign n5497 = n889 & n30458 ;
  assign n3314 = n2639 & n3311 ;
  assign n3347 = n30157 & n3343 ;
  assign n5503 = n3314 | n3347 ;
  assign n5504 = n30453 & n3329 ;
  assign n5505 = n5503 | n5504 ;
  assign n5506 = n5497 | n5505 ;
  assign n5507 = n5492 | n5506 ;
  assign n5508 = n5492 & n5506 ;
  assign n30459 = ~n5508 ;
  assign n5509 = n5507 & n30459 ;
  assign n5510 = n2204 | n2351 ;
  assign n5511 = n5407 | n5510 ;
  assign n5512 = n113 | n384 ;
  assign n5513 = n1513 | n1574 ;
  assign n5514 = n5512 | n5513 ;
  assign n5515 = n190 | n296 ;
  assign n5516 = n814 | n5515 ;
  assign n5517 = n1177 | n5516 ;
  assign n5518 = n5514 | n5517 ;
  assign n5519 = n5511 | n5518 ;
  assign n5520 = n150 | n2426 ;
  assign n5521 = n2748 | n5520 ;
  assign n5522 = n337 | n647 ;
  assign n5523 = n767 | n5522 ;
  assign n5524 = n127 & n209 ;
  assign n5525 = n5523 | n5524 ;
  assign n5526 = n5521 | n5525 ;
  assign n5527 = n1091 | n1179 ;
  assign n5528 = n5096 | n5527 ;
  assign n5529 = n3032 | n3682 ;
  assign n5530 = n5528 | n5529 ;
  assign n5531 = n5526 | n5530 ;
  assign n5532 = n5519 | n5531 ;
  assign n30460 = ~n5532 ;
  assign n5533 = n2035 & n30460 ;
  assign n5534 = n3529 | n4889 ;
  assign n5535 = n151 | n1967 ;
  assign n5536 = n5484 | n5535 ;
  assign n5537 = n5534 | n5536 ;
  assign n5538 = n901 | n2500 ;
  assign n5539 = n2653 | n3290 ;
  assign n5540 = n5538 | n5539 ;
  assign n5541 = n310 | n407 ;
  assign n5542 = n614 | n5541 ;
  assign n5543 = n1495 | n5542 ;
  assign n5544 = n1925 | n5543 ;
  assign n5545 = n5540 | n5544 ;
  assign n5546 = n5537 | n5545 ;
  assign n5547 = n1970 | n2352 ;
  assign n5548 = n3165 | n5547 ;
  assign n5549 = n552 | n5548 ;
  assign n5550 = n630 | n766 ;
  assign n5551 = n683 | n1047 ;
  assign n5552 = n5550 | n5551 ;
  assign n5553 = n1149 | n5552 ;
  assign n5554 = n5549 | n5553 ;
  assign n5555 = n162 | n245 ;
  assign n5556 = n440 | n608 ;
  assign n5557 = n5555 | n5556 ;
  assign n5558 = n215 | n946 ;
  assign n5559 = n5557 | n5558 ;
  assign n5560 = n1902 | n3738 ;
  assign n5561 = n5559 | n5560 ;
  assign n5562 = n5382 | n5561 ;
  assign n5563 = n5554 | n5562 ;
  assign n5564 = n5546 | n5563 ;
  assign n30461 = ~n5564 ;
  assign n5565 = n5533 & n30461 ;
  assign n2788 = n30155 & n2567 ;
  assign n2795 = n2639 & n2788 ;
  assign n5566 = n2639 | n2788 ;
  assign n30462 = ~n2795 ;
  assign n5567 = n30462 & n5566 ;
  assign n5568 = n889 & n5567 ;
  assign n3330 = n30155 & n3329 ;
  assign n3345 = n2639 & n3343 ;
  assign n5574 = n3330 | n3345 ;
  assign n30463 = ~n2567 ;
  assign n5575 = n30463 & n3311 ;
  assign n5576 = n5574 | n5575 ;
  assign n5577 = n5568 | n5576 ;
  assign n30464 = ~n5565 ;
  assign n5579 = n30464 & n5577 ;
  assign n30465 = ~n372 ;
  assign n5580 = n145 & n30465 ;
  assign n5581 = n516 | n1179 ;
  assign n30466 = ~n5581 ;
  assign n5582 = n5580 & n30466 ;
  assign n5583 = n2410 | n2951 ;
  assign n30467 = ~n5583 ;
  assign n5584 = n5582 & n30467 ;
  assign n5585 = n809 | n1546 ;
  assign n30468 = ~n5585 ;
  assign n5586 = n5584 & n30468 ;
  assign n5587 = n402 | n586 ;
  assign n5588 = n613 | n1050 ;
  assign n5589 = n5587 | n5588 ;
  assign n5590 = n158 | n500 ;
  assign n5591 = n3450 | n5590 ;
  assign n5592 = n212 | n257 ;
  assign n5593 = n865 | n5592 ;
  assign n5594 = n5591 | n5593 ;
  assign n5595 = n5589 | n5594 ;
  assign n5596 = n396 | n2025 ;
  assign n5597 = n2326 | n3247 ;
  assign n5598 = n248 | n448 ;
  assign n5599 = n4871 | n5598 ;
  assign n5600 = n5597 | n5599 ;
  assign n5601 = n5596 | n5600 ;
  assign n5602 = n5595 | n5601 ;
  assign n30469 = ~n5602 ;
  assign n5603 = n5586 & n30469 ;
  assign n5604 = n529 | n2746 ;
  assign n5605 = n233 | n5604 ;
  assign n5606 = n917 | n1099 ;
  assign n5607 = n263 | n348 ;
  assign n5608 = n698 | n5607 ;
  assign n5609 = n2017 | n2748 ;
  assign n5610 = n5608 | n5609 ;
  assign n5611 = n5606 | n5610 ;
  assign n5612 = n5605 | n5611 ;
  assign n5613 = n313 | n711 ;
  assign n5614 = n998 | n2403 ;
  assign n5615 = n5613 | n5614 ;
  assign n5616 = n82 & n2447 ;
  assign n5617 = n152 | n5616 ;
  assign n5618 = n1530 | n5617 ;
  assign n5619 = n5615 | n5618 ;
  assign n5620 = n5612 | n5619 ;
  assign n5621 = n2610 | n5620 ;
  assign n30470 = ~n5621 ;
  assign n5622 = n5603 & n30470 ;
  assign n30471 = ~n1259 ;
  assign n5623 = n30471 & n5622 ;
  assign n30472 = ~n5623 ;
  assign n5625 = n5579 & n30472 ;
  assign n5624 = n5579 & n5623 ;
  assign n5626 = n5579 | n5623 ;
  assign n30473 = ~n5624 ;
  assign n5627 = n30473 & n5626 ;
  assign n5628 = n2641 | n2794 ;
  assign n30474 = ~n5628 ;
  assign n5629 = n2701 & n30474 ;
  assign n5630 = n30453 & n5628 ;
  assign n5631 = n5629 | n5630 ;
  assign n5632 = n889 & n5631 ;
  assign n3315 = n30155 & n3311 ;
  assign n3344 = n30453 & n3343 ;
  assign n5638 = n3315 | n3344 ;
  assign n5639 = n2639 & n3329 ;
  assign n5640 = n5638 | n5639 ;
  assign n5641 = n5632 | n5640 ;
  assign n30475 = ~n5627 ;
  assign n5643 = n30475 & n5641 ;
  assign n5644 = n5625 | n5643 ;
  assign n30476 = ~n5644 ;
  assign n5646 = n5509 & n30476 ;
  assign n30477 = ~n5646 ;
  assign n5647 = n5507 & n30477 ;
  assign n5649 = n5458 | n5647 ;
  assign n30478 = ~n5456 ;
  assign n5650 = n30478 & n5649 ;
  assign n30479 = ~n5650 ;
  assign n5652 = n5405 & n30479 ;
  assign n30480 = ~n5652 ;
  assign n5653 = n5403 & n30480 ;
  assign n30481 = ~n5653 ;
  assign n5655 = n5348 & n30481 ;
  assign n30482 = ~n5655 ;
  assign n5656 = n5346 & n30482 ;
  assign n30483 = ~n4349 ;
  assign n5657 = n30483 & n4350 ;
  assign n5658 = n4362 & n5657 ;
  assign n5659 = n4362 | n5657 ;
  assign n30484 = ~n5658 ;
  assign n5660 = n30484 & n5659 ;
  assign n5662 = n5656 | n5660 ;
  assign n4379 = n895 & n30310 ;
  assign n2851 = n30114 & n2849 ;
  assign n2867 = n30123 & n2861 ;
  assign n5663 = n2851 | n2867 ;
  assign n5664 = n894 & n30108 ;
  assign n5665 = n5663 | n5664 ;
  assign n5666 = n4379 | n5665 ;
  assign n30485 = ~n5666 ;
  assign n5667 = x29 & n30485 ;
  assign n5668 = n30024 & n5666 ;
  assign n5669 = n5667 | n5668 ;
  assign n5661 = n5656 & n5660 ;
  assign n30486 = ~n5661 ;
  assign n5670 = n30486 & n5662 ;
  assign n30487 = ~n5669 ;
  assign n5671 = n30487 & n5670 ;
  assign n30488 = ~n5671 ;
  assign n5672 = n5662 & n30488 ;
  assign n5673 = n5282 & n5672 ;
  assign n5674 = n5281 | n5673 ;
  assign n5262 = n5249 | n5261 ;
  assign n5675 = n5249 & n5261 ;
  assign n30489 = ~n5675 ;
  assign n5676 = n5262 & n30489 ;
  assign n30490 = ~n5676 ;
  assign n5678 = n5674 & n30490 ;
  assign n5679 = n5263 | n5678 ;
  assign n5680 = n5245 | n5679 ;
  assign n3611 = n895 & n30233 ;
  assign n1673 = n894 & n30196 ;
  assign n2859 = n30105 & n2849 ;
  assign n5681 = n1673 | n2859 ;
  assign n5682 = n1812 & n2861 ;
  assign n5683 = n5681 | n5682 ;
  assign n5684 = n3611 | n5683 ;
  assign n30491 = ~n5684 ;
  assign n5685 = x29 & n30491 ;
  assign n5686 = n30024 & n5684 ;
  assign n5687 = n5685 | n5686 ;
  assign n5688 = n5245 & n5679 ;
  assign n30492 = ~n5688 ;
  assign n5689 = n5680 & n30492 ;
  assign n30493 = ~n5687 ;
  assign n5690 = n30493 & n5689 ;
  assign n30494 = ~n5690 ;
  assign n5691 = n5680 & n30494 ;
  assign n30495 = ~n5691 ;
  assign n5693 = n5243 & n30495 ;
  assign n3800 = n30238 & n3791 ;
  assign n1448 = n209 & n1445 ;
  assign n3817 = n30082 & n3802 ;
  assign n5694 = n1448 | n3817 ;
  assign n5695 = n1219 & n3818 ;
  assign n5696 = n5694 | n5695 ;
  assign n5697 = n3800 | n5696 ;
  assign n30496 = ~n5697 ;
  assign n5698 = x26 & n30496 ;
  assign n5699 = n30019 & n5697 ;
  assign n5700 = n5698 | n5699 ;
  assign n5692 = n5243 & n5691 ;
  assign n5701 = n5243 | n5691 ;
  assign n30497 = ~n5692 ;
  assign n5702 = n30497 & n5701 ;
  assign n5703 = n5700 | n5702 ;
  assign n30498 = ~n5693 ;
  assign n5704 = n30498 & n5703 ;
  assign n5706 = n5241 | n5704 ;
  assign n4143 = n3787 & n4135 ;
  assign n4149 = n3764 & n4148 ;
  assign n4193 = n1074 & n4185 ;
  assign n5707 = n4149 | n4193 ;
  assign n5708 = n3700 & n4165 ;
  assign n5709 = n5707 | n5708 ;
  assign n5710 = n4143 | n5709 ;
  assign n30499 = ~n5710 ;
  assign n5711 = x23 & n30499 ;
  assign n5712 = n30030 & n5710 ;
  assign n5713 = n5711 | n5712 ;
  assign n5705 = n5241 & n5704 ;
  assign n30500 = ~n5705 ;
  assign n5714 = n30500 & n5706 ;
  assign n30501 = ~n5713 ;
  assign n5715 = n30501 & n5714 ;
  assign n30502 = ~n5715 ;
  assign n5716 = n5706 & n30502 ;
  assign n30503 = ~n5716 ;
  assign n5718 = n5239 & n30503 ;
  assign n30504 = ~n5718 ;
  assign n5719 = n5237 & n30504 ;
  assign n5721 = n5226 | n5719 ;
  assign n4585 = n4583 & n4584 ;
  assign n5722 = n4583 | n4584 ;
  assign n30505 = ~n4585 ;
  assign n5723 = n30505 & n5722 ;
  assign n5724 = n4686 & n5723 ;
  assign n4740 = n4033 & n4726 ;
  assign n4757 = n30361 & n4748 ;
  assign n5730 = n4740 | n4757 ;
  assign n5731 = n30282 & n4706 ;
  assign n5732 = n5730 | n5731 ;
  assign n5733 = n5724 | n5732 ;
  assign n30506 = ~n5733 ;
  assign n5734 = x20 & n30506 ;
  assign n5735 = n30374 & n5733 ;
  assign n5736 = n5734 | n5735 ;
  assign n30507 = ~n5226 ;
  assign n5720 = n30507 & n5719 ;
  assign n30508 = ~n5719 ;
  assign n5737 = n5226 & n30508 ;
  assign n5738 = n5720 | n5737 ;
  assign n30509 = ~n5736 ;
  assign n5739 = n30509 & n5738 ;
  assign n30510 = ~n5739 ;
  assign n5740 = n5721 & n30510 ;
  assign n5742 = n5224 | n5740 ;
  assign n5131 = n5123 & n5130 ;
  assign n30511 = ~n5131 ;
  assign n5743 = n30511 & n5132 ;
  assign n30512 = ~n5743 ;
  assign n5744 = n37300 & n30512 ;
  assign n5153 = n30405 & n5144 ;
  assign n5190 = n4811 & n5166 ;
  assign n5750 = n5153 | n5190 ;
  assign n5751 = n5017 & n5191 ;
  assign n5752 = n5750 | n5751 ;
  assign n5753 = n5744 | n5752 ;
  assign n5754 = x17 | n5753 ;
  assign n5755 = x17 & n5753 ;
  assign n30513 = ~n5755 ;
  assign n5756 = n5754 & n30513 ;
  assign n5741 = n5224 & n5740 ;
  assign n30514 = ~n5741 ;
  assign n5757 = n30514 & n5742 ;
  assign n30515 = ~n5756 ;
  assign n5759 = n30515 & n5757 ;
  assign n30516 = ~n5759 ;
  assign n5760 = n5742 & n30516 ;
  assign n5761 = n5222 & n5760 ;
  assign n5762 = n5222 | n5760 ;
  assign n30517 = ~n5761 ;
  assign n5763 = n30517 & n5762 ;
  assign n5764 = n80 | n473 ;
  assign n30518 = ~n257 ;
  assign n5765 = n142 & n30518 ;
  assign n30519 = ~n5085 ;
  assign n5766 = n30519 & n5765 ;
  assign n30520 = ~n5764 ;
  assign n5767 = n30520 & n5766 ;
  assign n5768 = n358 | n529 ;
  assign n5769 = n688 | n5768 ;
  assign n5770 = n788 | n1249 ;
  assign n5771 = n5769 | n5770 ;
  assign n5772 = n542 | n554 ;
  assign n5773 = n865 | n5772 ;
  assign n5774 = n1352 | n5773 ;
  assign n5775 = n1714 | n5774 ;
  assign n5776 = n5771 | n5775 ;
  assign n2445 = x24 & n2444 ;
  assign n5777 = n102 | n2445 ;
  assign n5778 = n209 | n5777 ;
  assign n5779 = n192 & n5778 ;
  assign n5780 = n2224 | n2952 ;
  assign n5781 = n3736 | n5780 ;
  assign n5782 = n335 | n1311 ;
  assign n5783 = n1662 | n2139 ;
  assign n5784 = n5782 | n5783 ;
  assign n5785 = n5781 | n5784 ;
  assign n5786 = n5779 | n5785 ;
  assign n5787 = n5776 | n5786 ;
  assign n5788 = n249 | n5787 ;
  assign n30521 = ~n129 ;
  assign n2446 = n30521 & n2444 ;
  assign n30522 = ~n95 ;
  assign n5789 = n79 & n30522 ;
  assign n5790 = n2446 & n5789 ;
  assign n5791 = n309 | n5790 ;
  assign n5792 = n5788 | n5791 ;
  assign n30523 = ~n5792 ;
  assign n5793 = n5767 & n30523 ;
  assign n5800 = n164 | n280 ;
  assign n5801 = n431 | n722 ;
  assign n5802 = n1320 | n5072 ;
  assign n5803 = n5801 | n5802 ;
  assign n5804 = n5800 | n5803 ;
  assign n5805 = n205 | n289 ;
  assign n5806 = n232 | n432 ;
  assign n5807 = n5805 | n5806 ;
  assign n5808 = n354 | n553 ;
  assign n5809 = n1211 | n5808 ;
  assign n5810 = n5807 | n5809 ;
  assign n5811 = n659 | n2718 ;
  assign n30524 = ~n5811 ;
  assign n5812 = n4527 & n30524 ;
  assign n30525 = ~n5810 ;
  assign n5813 = n30525 & n5812 ;
  assign n30526 = ~n5804 ;
  assign n5814 = n30526 & n5813 ;
  assign n5815 = n395 | n1166 ;
  assign n5816 = n138 | n996 ;
  assign n5817 = n2052 | n5816 ;
  assign n5818 = n5815 | n5817 ;
  assign n5819 = n2694 | n5818 ;
  assign n5820 = n2450 | n5819 ;
  assign n5821 = n793 | n816 ;
  assign n5822 = n521 | n5821 ;
  assign n5823 = n497 | n1712 ;
  assign n5824 = n572 | n5823 ;
  assign n5825 = n5822 | n5824 ;
  assign n5826 = n5070 | n5825 ;
  assign n5827 = n5820 | n5826 ;
  assign n30527 = ~n5827 ;
  assign n5828 = n5814 & n30527 ;
  assign n5829 = n244 | n276 ;
  assign n5830 = n516 | n1010 ;
  assign n5831 = n713 | n5830 ;
  assign n5832 = n5829 | n5831 ;
  assign n5833 = n2676 | n5832 ;
  assign n5834 = n1366 | n5833 ;
  assign n5835 = n764 | n5834 ;
  assign n5836 = n721 | n5835 ;
  assign n5837 = n2050 | n3480 ;
  assign n5838 = n4918 | n5837 ;
  assign n5839 = n204 | n433 ;
  assign n5840 = n272 | n460 ;
  assign n5841 = n509 | n695 ;
  assign n5842 = n5840 | n5841 ;
  assign n5843 = n5839 | n5842 ;
  assign n5844 = n5838 | n5843 ;
  assign n5845 = n4888 | n5844 ;
  assign n5846 = n4897 | n4907 ;
  assign n5847 = n5845 | n5846 ;
  assign n5848 = n5836 | n5847 ;
  assign n30528 = ~n5848 ;
  assign n5849 = n5828 & n30528 ;
  assign n5850 = n224 | n797 ;
  assign n5851 = n2389 | n5850 ;
  assign n5852 = n2628 | n5851 ;
  assign n5853 = n2179 | n5852 ;
  assign n5854 = n376 | n3736 ;
  assign n5855 = n282 | n991 ;
  assign n5856 = n2335 | n5855 ;
  assign n5857 = n5854 | n5856 ;
  assign n5858 = n5009 | n5857 ;
  assign n5859 = n5853 | n5858 ;
  assign n5860 = n332 | n491 ;
  assign n5861 = n359 | n1091 ;
  assign n5862 = n269 | n5861 ;
  assign n5863 = n5860 | n5862 ;
  assign n5864 = n2761 | n3852 ;
  assign n5865 = n5863 | n5864 ;
  assign n5866 = n368 | n689 ;
  assign n5867 = n5790 | n5866 ;
  assign n5868 = n5865 | n5867 ;
  assign n5869 = n5859 | n5868 ;
  assign n30529 = ~n5869 ;
  assign n5870 = n5849 & n30529 ;
  assign n5877 = n30415 & n5870 ;
  assign n30530 = ~n5870 ;
  assign n5878 = n4925 & n30530 ;
  assign n5879 = n5877 | n5878 ;
  assign n5880 = n4925 & n30404 ;
  assign n30531 = ~n5880 ;
  assign n5881 = n5134 & n30531 ;
  assign n30532 = ~n5881 ;
  assign n5883 = n5879 & n30532 ;
  assign n5884 = n4925 & n5870 ;
  assign n5885 = n5883 | n5884 ;
  assign n5886 = n429 | n689 ;
  assign n5887 = n401 | n476 ;
  assign n5888 = n635 | n676 ;
  assign n5889 = n5887 | n5888 ;
  assign n5890 = n269 | n346 ;
  assign n5891 = n1035 | n5890 ;
  assign n5892 = n1500 | n5891 ;
  assign n5893 = n5889 | n5892 ;
  assign n5894 = n5886 | n5893 ;
  assign n5895 = n379 | n978 ;
  assign n5896 = n5853 | n5895 ;
  assign n5897 = n5894 | n5896 ;
  assign n5898 = n2168 | n5897 ;
  assign n5901 = n99 | n1047 ;
  assign n3801 = n121 | n260 ;
  assign n5902 = x26 & n213 ;
  assign n5903 = n3801 & n5902 ;
  assign n5904 = n5901 | n5903 ;
  assign n5905 = n445 | n2584 ;
  assign n5906 = n3753 | n5905 ;
  assign n5907 = n4916 | n5906 ;
  assign n5908 = n5904 | n5907 ;
  assign n5909 = n5898 | n5908 ;
  assign n5910 = n309 | n679 ;
  assign n30533 = ~n5910 ;
  assign n5911 = n5767 & n30533 ;
  assign n30534 = ~n5909 ;
  assign n5912 = n30534 & n5911 ;
  assign n30535 = ~n5912 ;
  assign n5918 = n5870 & n30535 ;
  assign n5919 = n5885 & n5918 ;
  assign n5920 = n30530 & n5912 ;
  assign n30536 = ~n5883 ;
  assign n5921 = n30536 & n5920 ;
  assign n5922 = n5919 | n5921 ;
  assign n5923 = n5793 | n5922 ;
  assign n5924 = n5793 & n5922 ;
  assign n30537 = ~n5924 ;
  assign n5925 = n5923 & n30537 ;
  assign n29896 = x11 & x12 ;
  assign n5932 = x11 | x12 ;
  assign n30538 = ~n29896 ;
  assign n5934 = n30538 & n5932 ;
  assign n37288 = x13 & x14 ;
  assign n5935 = x13 | x14 ;
  assign n30539 = ~n37288 ;
  assign n5936 = n30539 & n5935 ;
  assign n5937 = n5934 & n5936 ;
  assign n30540 = ~n5925 ;
  assign n5948 = n30540 & n5937 ;
  assign n30541 = ~n5932 ;
  assign n5933 = x13 & n30541 ;
  assign n30542 = ~x13 ;
  assign n5969 = n30542 & n29896 ;
  assign n5970 = n5933 | n5969 ;
  assign n5992 = n5934 | n5970 ;
  assign n30543 = ~n5992 ;
  assign n5994 = n5936 & n30543 ;
  assign n6007 = n30530 & n5994 ;
  assign n30544 = ~n5936 ;
  assign n6018 = n5934 & n30544 ;
  assign n30545 = ~n5793 ;
  assign n6031 = n30545 & n6018 ;
  assign n6043 = n6007 | n6031 ;
  assign n6044 = n30535 & n5970 ;
  assign n6045 = n6043 | n6044 ;
  assign n6046 = n5948 | n6045 ;
  assign n30546 = ~n6046 ;
  assign n6047 = x14 & n30546 ;
  assign n30547 = ~x14 ;
  assign n6048 = n30547 & n6046 ;
  assign n6049 = n6047 | n6048 ;
  assign n6050 = n5763 | n6049 ;
  assign n6051 = n5763 & n6049 ;
  assign n30548 = ~n6051 ;
  assign n6052 = n6050 & n30548 ;
  assign n5758 = n5756 & n5757 ;
  assign n6053 = n5756 | n5757 ;
  assign n30549 = ~n5758 ;
  assign n6054 = n30549 & n6053 ;
  assign n30550 = ~n5738 ;
  assign n6055 = n5736 & n30550 ;
  assign n6056 = n5739 | n6055 ;
  assign n5717 = n5239 & n5716 ;
  assign n6057 = n5239 | n5716 ;
  assign n30551 = ~n5717 ;
  assign n6058 = n30551 & n6057 ;
  assign n30552 = ~n5714 ;
  assign n6059 = n5713 & n30552 ;
  assign n6060 = n5715 | n6059 ;
  assign n6061 = n5700 & n5702 ;
  assign n30553 = ~n6061 ;
  assign n6062 = n5703 & n30553 ;
  assign n3792 = n30203 & n3791 ;
  assign n1560 = n209 & n1556 ;
  assign n3809 = n1445 & n3802 ;
  assign n6063 = n1560 | n3809 ;
  assign n6064 = n30082 & n3818 ;
  assign n6065 = n6063 | n6064 ;
  assign n6066 = n3792 | n6065 ;
  assign n6067 = x26 | n6066 ;
  assign n6068 = x26 & n6066 ;
  assign n30554 = ~n6068 ;
  assign n6069 = n6067 & n30554 ;
  assign n5677 = n5674 | n5676 ;
  assign n6070 = n5674 & n5676 ;
  assign n30555 = ~n6070 ;
  assign n6071 = n5677 & n30555 ;
  assign n4232 = n895 & n4230 ;
  assign n1755 = n894 & n30105 ;
  assign n2854 = n1812 & n2849 ;
  assign n6072 = n1755 | n2854 ;
  assign n6073 = n30108 & n2861 ;
  assign n6074 = n6072 | n6073 ;
  assign n6075 = n4232 | n6074 ;
  assign n6076 = x29 | n6075 ;
  assign n6077 = x29 & n6075 ;
  assign n30556 = ~n6077 ;
  assign n6078 = n6076 & n30556 ;
  assign n30557 = ~n6078 ;
  assign n6080 = n6071 & n30557 ;
  assign n3794 = n30209 & n3791 ;
  assign n1672 = n209 & n30196 ;
  assign n3815 = n1556 & n3802 ;
  assign n6081 = n1672 | n3815 ;
  assign n6082 = n1445 & n3818 ;
  assign n6083 = n6081 | n6082 ;
  assign n6084 = n3794 | n6083 ;
  assign n30558 = ~n6084 ;
  assign n6085 = x26 & n30558 ;
  assign n6086 = n30019 & n6084 ;
  assign n6087 = n6085 | n6086 ;
  assign n30559 = ~n6071 ;
  assign n6079 = n30559 & n6078 ;
  assign n6088 = n6079 | n6080 ;
  assign n6089 = n6087 | n6088 ;
  assign n30560 = ~n6080 ;
  assign n6090 = n30560 & n6089 ;
  assign n6091 = n6069 & n6090 ;
  assign n30561 = ~n5689 ;
  assign n6092 = n5687 & n30561 ;
  assign n6093 = n5690 | n6092 ;
  assign n6094 = n6069 | n6090 ;
  assign n30562 = ~n6091 ;
  assign n6095 = n30562 & n6094 ;
  assign n6097 = n6093 & n6095 ;
  assign n6098 = n6091 | n6097 ;
  assign n30563 = ~n6098 ;
  assign n6099 = n6062 & n30563 ;
  assign n4423 = n4135 & n4420 ;
  assign n4152 = n1074 & n4148 ;
  assign n4174 = n3764 & n4165 ;
  assign n6100 = n4152 | n4174 ;
  assign n6101 = n30074 & n4185 ;
  assign n6102 = n6100 | n6101 ;
  assign n6103 = n4423 | n6102 ;
  assign n30564 = ~n6103 ;
  assign n6104 = x23 & n30564 ;
  assign n6105 = n30030 & n6103 ;
  assign n6106 = n6104 | n6105 ;
  assign n30565 = ~n6062 ;
  assign n6107 = n30565 & n6098 ;
  assign n6108 = n6099 | n6107 ;
  assign n6109 = n6106 | n6108 ;
  assign n30566 = ~n6099 ;
  assign n6110 = n30566 & n6109 ;
  assign n6112 = n6060 | n6110 ;
  assign n4693 = n4442 & n4686 ;
  assign n4710 = n4093 & n4706 ;
  assign n4727 = n30264 & n4726 ;
  assign n6113 = n4710 | n4727 ;
  assign n6114 = n4033 & n4748 ;
  assign n6115 = n6113 | n6114 ;
  assign n6116 = n4693 | n6115 ;
  assign n30567 = ~n6116 ;
  assign n6117 = x20 & n30567 ;
  assign n6118 = n30374 & n6116 ;
  assign n6119 = n6117 | n6118 ;
  assign n30568 = ~n6060 ;
  assign n6111 = n30568 & n6110 ;
  assign n30569 = ~n6110 ;
  assign n6120 = n6060 & n30569 ;
  assign n6121 = n6111 | n6120 ;
  assign n30570 = ~n6119 ;
  assign n6122 = n30570 & n6121 ;
  assign n30571 = ~n6122 ;
  assign n6123 = n6112 & n30571 ;
  assign n6125 = n6058 | n6123 ;
  assign n4690 = n30286 & n4686 ;
  assign n4739 = n4093 & n4726 ;
  assign n4755 = n30282 & n4748 ;
  assign n6126 = n4739 | n4755 ;
  assign n6127 = n4033 & n4706 ;
  assign n6128 = n6126 | n6127 ;
  assign n6129 = n4690 | n6128 ;
  assign n30572 = ~n6129 ;
  assign n6130 = x20 & n30572 ;
  assign n6131 = n30374 & n6129 ;
  assign n6132 = n6130 | n6131 ;
  assign n30573 = ~n6058 ;
  assign n6124 = n30573 & n6123 ;
  assign n30574 = ~n6123 ;
  assign n6133 = n6058 & n30574 ;
  assign n6134 = n6124 | n6133 ;
  assign n30575 = ~n6132 ;
  assign n6135 = n30575 & n6134 ;
  assign n30576 = ~n6135 ;
  assign n6136 = n6125 & n30576 ;
  assign n6138 = n6056 | n6136 ;
  assign n6139 = n5125 & n5128 ;
  assign n30577 = ~n6139 ;
  assign n6140 = n5129 & n30577 ;
  assign n30578 = ~n6140 ;
  assign n6141 = n37300 & n30578 ;
  assign n5146 = n4811 & n5144 ;
  assign n5176 = n4664 & n5166 ;
  assign n6148 = n5146 | n5176 ;
  assign n6149 = n30405 & n5191 ;
  assign n6150 = n6148 | n6149 ;
  assign n6151 = n6141 | n6150 ;
  assign n30579 = ~n6151 ;
  assign n6152 = x17 & n30579 ;
  assign n30580 = ~x17 ;
  assign n6153 = n30580 & n6151 ;
  assign n6154 = n6152 | n6153 ;
  assign n30581 = ~n6056 ;
  assign n6137 = n30581 & n6136 ;
  assign n30582 = ~n6136 ;
  assign n6155 = n6056 & n30582 ;
  assign n6156 = n6137 | n6155 ;
  assign n30583 = ~n6154 ;
  assign n6157 = n30583 & n6156 ;
  assign n30584 = ~n6157 ;
  assign n6158 = n6138 & n30584 ;
  assign n6159 = n6054 & n6158 ;
  assign n6160 = n5918 | n5920 ;
  assign n30585 = ~n6160 ;
  assign n6161 = n5885 & n30585 ;
  assign n30586 = ~n5885 ;
  assign n6162 = n30586 & n6160 ;
  assign n6163 = n6161 | n6162 ;
  assign n30587 = ~n6163 ;
  assign n6164 = n5937 & n30587 ;
  assign n5983 = n30530 & n5970 ;
  assign n6009 = n30415 & n5994 ;
  assign n6171 = n5983 | n6009 ;
  assign n6172 = n30535 & n6018 ;
  assign n6173 = n6171 | n6172 ;
  assign n6174 = n6164 | n6173 ;
  assign n6175 = x14 | n6174 ;
  assign n6176 = x14 & n6174 ;
  assign n30588 = ~n6176 ;
  assign n6177 = n6175 & n30588 ;
  assign n6178 = n6054 | n6158 ;
  assign n30589 = ~n6159 ;
  assign n6179 = n30589 & n6178 ;
  assign n6180 = n6177 & n6179 ;
  assign n6181 = n6159 | n6180 ;
  assign n30590 = ~n6181 ;
  assign n6182 = n6052 & n30590 ;
  assign n30591 = ~n6052 ;
  assign n6183 = n30591 & n6181 ;
  assign n6184 = n6182 | n6183 ;
  assign n29897 = x8 & x9 ;
  assign n6185 = x8 | x9 ;
  assign n30592 = ~n29897 ;
  assign n6188 = n30592 & n6185 ;
  assign n30593 = ~n6185 ;
  assign n6186 = x10 & n30593 ;
  assign n30594 = ~x10 ;
  assign n6189 = n30594 & n29897 ;
  assign n6190 = n6186 | n6189 ;
  assign n6213 = n6188 | n6190 ;
  assign n37289 = x10 & x11 ;
  assign n6215 = x10 | x11 ;
  assign n30595 = ~n37289 ;
  assign n6216 = n30595 & n6215 ;
  assign n30596 = ~n6213 ;
  assign n6244 = n30596 & n6216 ;
  assign n6265 = n5870 | n5885 ;
  assign n6266 = n5912 & n6265 ;
  assign n6272 = n6188 & n6216 ;
  assign n30597 = ~n6266 ;
  assign n6288 = n30597 & n6272 ;
  assign n6307 = n6244 | n6288 ;
  assign n6308 = n30545 & n6307 ;
  assign n6309 = x11 & n6308 ;
  assign n6310 = x11 | n6308 ;
  assign n30598 = ~n6309 ;
  assign n6311 = n30598 & n6310 ;
  assign n30599 = ~n6156 ;
  assign n6312 = n6154 & n30599 ;
  assign n6313 = n6157 | n6312 ;
  assign n4839 = n37300 & n30385 ;
  assign n5169 = n30361 & n5166 ;
  assign n5205 = n4811 & n5191 ;
  assign n6314 = n5169 | n5205 ;
  assign n6315 = n4664 & n5144 ;
  assign n6316 = n6314 | n6315 ;
  assign n6317 = n4839 | n6316 ;
  assign n6318 = x17 | n6317 ;
  assign n6319 = x17 & n6317 ;
  assign n30600 = ~n6319 ;
  assign n6320 = n6318 & n30600 ;
  assign n30601 = ~n6121 ;
  assign n6321 = n6119 & n30601 ;
  assign n6322 = n6122 | n6321 ;
  assign n6323 = n6106 & n6108 ;
  assign n30602 = ~n6323 ;
  assign n6324 = n6109 & n30602 ;
  assign n30603 = ~n6093 ;
  assign n6096 = n30603 & n6095 ;
  assign n30604 = ~n6095 ;
  assign n6325 = n6093 & n30604 ;
  assign n6326 = n6096 | n6325 ;
  assign n6327 = n6087 & n6088 ;
  assign n30605 = ~n6327 ;
  assign n6328 = n6089 & n30605 ;
  assign n6329 = n5282 | n5672 ;
  assign n30606 = ~n5673 ;
  assign n6330 = n30606 & n6329 ;
  assign n3594 = n895 & n3592 ;
  assign n1815 = n894 & n1812 ;
  assign n2862 = n30114 & n2861 ;
  assign n6331 = n1815 | n2862 ;
  assign n6332 = n30108 & n2849 ;
  assign n6333 = n6331 | n6332 ;
  assign n6334 = n3594 | n6333 ;
  assign n6335 = x29 | n6334 ;
  assign n6336 = x29 & n6334 ;
  assign n30607 = ~n6336 ;
  assign n6337 = n6335 & n30607 ;
  assign n6338 = n6330 & n6337 ;
  assign n3799 = n3307 & n3791 ;
  assign n3805 = n30196 & n3802 ;
  assign n3826 = n1556 & n3818 ;
  assign n6339 = n3805 | n3826 ;
  assign n6340 = n209 & n30105 ;
  assign n6341 = n6339 | n6340 ;
  assign n6342 = n3799 | n6341 ;
  assign n6343 = x26 | n6342 ;
  assign n6344 = x26 & n6342 ;
  assign n30608 = ~n6344 ;
  assign n6345 = n6343 & n30608 ;
  assign n6346 = n6330 | n6337 ;
  assign n30609 = ~n6338 ;
  assign n6347 = n30609 & n6346 ;
  assign n6348 = n6345 & n6347 ;
  assign n6349 = n6338 | n6348 ;
  assign n30610 = ~n6328 ;
  assign n6351 = n30610 & n6349 ;
  assign n4141 = n30212 & n4135 ;
  assign n4155 = n1219 & n4148 ;
  assign n4192 = n30082 & n4185 ;
  assign n6352 = n4155 | n4192 ;
  assign n6353 = n30074 & n4165 ;
  assign n6354 = n6352 | n6353 ;
  assign n6355 = n4141 | n6354 ;
  assign n30611 = ~n6355 ;
  assign n6356 = x23 & n30611 ;
  assign n6357 = n30030 & n6355 ;
  assign n6358 = n6356 | n6357 ;
  assign n30612 = ~n6349 ;
  assign n6350 = n6328 & n30612 ;
  assign n6359 = n6350 | n6351 ;
  assign n30613 = ~n6359 ;
  assign n6361 = n6358 & n30613 ;
  assign n6362 = n6351 | n6361 ;
  assign n6364 = n6326 | n6362 ;
  assign n30614 = ~n6362 ;
  assign n6363 = n6326 & n30614 ;
  assign n30615 = ~n6326 ;
  assign n6365 = n30615 & n6362 ;
  assign n6366 = n6363 | n6365 ;
  assign n4146 = n30173 & n4135 ;
  assign n4173 = n1074 & n4165 ;
  assign n4194 = n1219 & n4185 ;
  assign n6367 = n4173 | n4194 ;
  assign n6368 = n30074 & n4148 ;
  assign n6369 = n6367 | n6368 ;
  assign n6370 = n4146 | n6369 ;
  assign n30616 = ~n6370 ;
  assign n6371 = x23 & n30616 ;
  assign n6372 = n30030 & n6370 ;
  assign n6373 = n6371 | n6372 ;
  assign n30617 = ~n6373 ;
  assign n6374 = n6366 & n30617 ;
  assign n30618 = ~n6374 ;
  assign n6375 = n6364 & n30618 ;
  assign n30619 = ~n6324 ;
  assign n6377 = n30619 & n6375 ;
  assign n4704 = n30349 & n4686 ;
  assign n4738 = n3700 & n4726 ;
  assign n4760 = n4093 & n4748 ;
  assign n6378 = n4738 | n4760 ;
  assign n6379 = n30264 & n4706 ;
  assign n6380 = n6378 | n6379 ;
  assign n6381 = n4704 | n6380 ;
  assign n30620 = ~n6381 ;
  assign n6382 = x20 & n30620 ;
  assign n6383 = n30374 & n6381 ;
  assign n6384 = n6382 | n6383 ;
  assign n6376 = n6324 & n6375 ;
  assign n6385 = n6324 | n6375 ;
  assign n30621 = ~n6376 ;
  assign n6386 = n30621 & n6385 ;
  assign n30622 = ~n6386 ;
  assign n6388 = n6384 & n30622 ;
  assign n6389 = n6377 | n6388 ;
  assign n6390 = n6322 | n6389 ;
  assign n6391 = n6322 & n6389 ;
  assign n30623 = ~n6391 ;
  assign n6392 = n6390 & n30623 ;
  assign n4675 = n37300 & n4674 ;
  assign n5152 = n30361 & n5144 ;
  assign n5203 = n4664 & n5191 ;
  assign n6393 = n5152 | n5203 ;
  assign n6394 = n30282 & n5166 ;
  assign n6395 = n6393 | n6394 ;
  assign n6396 = n4675 | n6395 ;
  assign n30624 = ~n6396 ;
  assign n6397 = x17 & n30624 ;
  assign n6398 = n30580 & n6396 ;
  assign n6399 = n6397 | n6398 ;
  assign n30625 = ~n6399 ;
  assign n6400 = n6392 & n30625 ;
  assign n30626 = ~n6400 ;
  assign n6401 = n6390 & n30626 ;
  assign n6402 = n6320 & n6401 ;
  assign n30627 = ~n6134 ;
  assign n6403 = n6132 & n30627 ;
  assign n6404 = n6135 | n6403 ;
  assign n6405 = n6320 | n6401 ;
  assign n30628 = ~n6402 ;
  assign n6406 = n30628 & n6405 ;
  assign n6408 = n6404 & n6406 ;
  assign n6409 = n6402 | n6408 ;
  assign n6410 = n6313 | n6409 ;
  assign n30629 = ~n5879 ;
  assign n5882 = n30629 & n5881 ;
  assign n6411 = n5882 | n5883 ;
  assign n6412 = n5937 & n6411 ;
  assign n5982 = n30415 & n5970 ;
  assign n6006 = n5017 & n5994 ;
  assign n6420 = n5982 | n6006 ;
  assign n6421 = n30530 & n6018 ;
  assign n6422 = n6420 | n6421 ;
  assign n6423 = n6412 | n6422 ;
  assign n30630 = ~n6423 ;
  assign n6424 = x14 & n30630 ;
  assign n6425 = n30547 & n6423 ;
  assign n6426 = n6424 | n6425 ;
  assign n6427 = n6313 & n6409 ;
  assign n30631 = ~n6427 ;
  assign n6428 = n6410 & n30631 ;
  assign n30632 = ~n6426 ;
  assign n6429 = n30632 & n6428 ;
  assign n30633 = ~n6429 ;
  assign n6430 = n6410 & n30633 ;
  assign n6432 = n6311 | n6430 ;
  assign n6433 = n6177 | n6179 ;
  assign n30634 = ~n6180 ;
  assign n6434 = n30634 & n6433 ;
  assign n6431 = n6311 & n6430 ;
  assign n30635 = ~n6431 ;
  assign n6435 = n30635 & n6432 ;
  assign n30636 = ~n6434 ;
  assign n6436 = n30636 & n6435 ;
  assign n30637 = ~n6436 ;
  assign n6437 = n6432 & n30637 ;
  assign n30638 = ~n6184 ;
  assign n6438 = n30638 & n6437 ;
  assign n30639 = ~n6437 ;
  assign n6439 = n6184 & n30639 ;
  assign n6440 = n6438 | n6439 ;
  assign n30640 = ~n6435 ;
  assign n6441 = n6434 & n30640 ;
  assign n6442 = n6436 | n6441 ;
  assign n5917 = n30523 & n5912 ;
  assign n6443 = n142 | n5912 ;
  assign n30641 = ~n5917 ;
  assign n6444 = n30641 & n6443 ;
  assign n30642 = ~n5922 ;
  assign n6445 = n30642 & n6444 ;
  assign n6446 = n6272 & n6445 ;
  assign n6454 = n30545 & n6190 ;
  assign n6455 = n30535 & n6244 ;
  assign n6456 = n6454 | n6455 ;
  assign n6457 = n6446 | n6456 ;
  assign n6458 = x11 | n6457 ;
  assign n6459 = x11 & n6457 ;
  assign n30643 = ~n6459 ;
  assign n6460 = n6458 & n30643 ;
  assign n5964 = n30410 & n5937 ;
  assign n6013 = n30405 & n5994 ;
  assign n6030 = n30415 & n6018 ;
  assign n6461 = n6013 | n6030 ;
  assign n6462 = n5017 & n5970 ;
  assign n6463 = n6461 | n6462 ;
  assign n6464 = n5964 | n6463 ;
  assign n6465 = x14 | n6464 ;
  assign n6466 = x14 & n6464 ;
  assign n30644 = ~n6466 ;
  assign n6467 = n6465 & n30644 ;
  assign n30645 = ~n6392 ;
  assign n6468 = n30645 & n6399 ;
  assign n6469 = n6400 | n6468 ;
  assign n6387 = n6384 | n6386 ;
  assign n6470 = n6384 & n6386 ;
  assign n30646 = ~n6470 ;
  assign n6471 = n6387 & n30646 ;
  assign n30647 = ~n6366 ;
  assign n6472 = n30647 & n6373 ;
  assign n6473 = n6374 | n6472 ;
  assign n6360 = n6358 | n6359 ;
  assign n6474 = n6358 & n6359 ;
  assign n30648 = ~n6474 ;
  assign n6475 = n6360 & n30648 ;
  assign n6476 = n6345 | n6347 ;
  assign n30649 = ~n6348 ;
  assign n6477 = n30649 & n6476 ;
  assign n30650 = ~n5670 ;
  assign n6478 = n5669 & n30650 ;
  assign n6479 = n5671 | n6478 ;
  assign n5654 = n5348 & n5653 ;
  assign n6480 = n5348 | n5653 ;
  assign n30651 = ~n5654 ;
  assign n6481 = n30651 & n6480 ;
  assign n5253 = n895 & n5251 ;
  assign n1958 = n894 & n30114 ;
  assign n2855 = n30123 & n2849 ;
  assign n6482 = n1958 | n2855 ;
  assign n6483 = n2102 & n2861 ;
  assign n6484 = n6482 | n6483 ;
  assign n6485 = n5253 | n6484 ;
  assign n6486 = x29 | n6485 ;
  assign n6487 = x29 & n6485 ;
  assign n30652 = ~n6487 ;
  assign n6488 = n6486 & n30652 ;
  assign n6490 = n6481 | n6488 ;
  assign n30653 = ~n6481 ;
  assign n6489 = n30653 & n6488 ;
  assign n30654 = ~n6488 ;
  assign n6491 = n6481 & n30654 ;
  assign n6492 = n6489 | n6491 ;
  assign n5651 = n5405 & n5650 ;
  assign n6493 = n5405 | n5650 ;
  assign n30655 = ~n5651 ;
  assign n6494 = n30655 & n6493 ;
  assign n5272 = n895 & n30440 ;
  assign n2856 = n2102 & n2849 ;
  assign n2865 = n2216 & n2861 ;
  assign n6495 = n2856 | n2865 ;
  assign n6496 = n894 & n30123 ;
  assign n6497 = n6495 | n6496 ;
  assign n6498 = n5272 | n6497 ;
  assign n6499 = x29 | n6498 ;
  assign n6500 = x29 & n6498 ;
  assign n30656 = ~n6500 ;
  assign n6501 = n6499 & n30656 ;
  assign n6503 = n6494 | n6501 ;
  assign n30657 = ~n6494 ;
  assign n6502 = n30657 & n6501 ;
  assign n30658 = ~n6501 ;
  assign n6504 = n6494 & n30658 ;
  assign n6505 = n6502 | n6504 ;
  assign n30659 = ~n5458 ;
  assign n5648 = n30659 & n5647 ;
  assign n30660 = ~n5647 ;
  assign n6506 = n5458 & n30660 ;
  assign n6507 = n5648 | n6506 ;
  assign n4353 = n895 & n4352 ;
  assign n2106 = n894 & n2102 ;
  assign n2872 = n2295 & n2861 ;
  assign n6508 = n2106 | n2872 ;
  assign n6509 = n2216 & n2849 ;
  assign n6510 = n6508 | n6509 ;
  assign n6511 = n4353 | n6510 ;
  assign n6512 = x29 | n6511 ;
  assign n6513 = x29 & n6511 ;
  assign n30661 = ~n6513 ;
  assign n6514 = n6512 & n30661 ;
  assign n30662 = ~n6514 ;
  assign n6516 = n6507 & n30662 ;
  assign n30663 = ~n6507 ;
  assign n6515 = n30663 & n6514 ;
  assign n6517 = n6515 | n6516 ;
  assign n5645 = n5509 | n5644 ;
  assign n6518 = n5509 & n5644 ;
  assign n30664 = ~n6518 ;
  assign n6519 = n5645 & n30664 ;
  assign n5337 = n895 & n30444 ;
  assign n2220 = n894 & n2216 ;
  assign n2852 = n2295 & n2849 ;
  assign n6520 = n2220 | n2852 ;
  assign n6521 = n30445 & n2861 ;
  assign n6522 = n6520 | n6521 ;
  assign n6523 = n5337 | n6522 ;
  assign n6524 = x29 | n6523 ;
  assign n6525 = x29 & n6523 ;
  assign n30665 = ~n6525 ;
  assign n6526 = n6524 & n30665 ;
  assign n6528 = n6519 | n6526 ;
  assign n5642 = n5627 | n5641 ;
  assign n6529 = n5627 & n5641 ;
  assign n30666 = ~n6529 ;
  assign n6530 = n5642 & n30666 ;
  assign n5394 = n895 & n5392 ;
  assign n2298 = n894 & n2295 ;
  assign n2873 = n30157 & n2861 ;
  assign n6531 = n2298 | n2873 ;
  assign n6532 = n30445 & n2849 ;
  assign n6533 = n6531 | n6532 ;
  assign n6534 = n5394 | n6533 ;
  assign n6535 = x29 | n6534 ;
  assign n6536 = x29 & n6534 ;
  assign n30667 = ~n6536 ;
  assign n6537 = n6535 & n30667 ;
  assign n30668 = ~n6537 ;
  assign n6539 = n6530 & n30668 ;
  assign n6538 = n6530 & n6537 ;
  assign n6540 = n6530 | n6537 ;
  assign n30669 = ~n6538 ;
  assign n6541 = n30669 & n6540 ;
  assign n30670 = ~n5577 ;
  assign n5578 = n5565 & n30670 ;
  assign n6542 = n5578 | n5579 ;
  assign n5447 = n895 & n30452 ;
  assign n2377 = n894 & n30445 ;
  assign n2857 = n30157 & n2849 ;
  assign n6543 = n2377 | n2857 ;
  assign n6544 = n30453 & n2861 ;
  assign n6545 = n6543 | n6544 ;
  assign n6546 = n5447 | n6545 ;
  assign n6547 = x29 | n6546 ;
  assign n6548 = x29 & n6546 ;
  assign n30671 = ~n6548 ;
  assign n6549 = n6547 & n30671 ;
  assign n30672 = ~n6542 ;
  assign n6550 = n30672 & n6549 ;
  assign n30673 = ~n6549 ;
  assign n6551 = n6542 & n30673 ;
  assign n6552 = n6550 | n6551 ;
  assign n5498 = n895 & n30458 ;
  assign n2781 = n894 & n30157 ;
  assign n2868 = n2639 & n2861 ;
  assign n6553 = n2781 | n2868 ;
  assign n6554 = n30453 & n2849 ;
  assign n6555 = n6553 | n6554 ;
  assign n6556 = n5498 | n6555 ;
  assign n6557 = x29 | n6556 ;
  assign n6558 = x29 & n6556 ;
  assign n30674 = ~n6558 ;
  assign n6559 = n6557 & n30674 ;
  assign n2789 = n108 & n30155 ;
  assign n30675 = ~n2789 ;
  assign n6560 = n2567 & n30675 ;
  assign n6561 = x31 & n30061 ;
  assign n30676 = ~n6561 ;
  assign n6563 = n2471 & n30676 ;
  assign n6562 = n30197 & n77 ;
  assign n6564 = n2640 | n6562 ;
  assign n30677 = ~n6563 ;
  assign n6565 = n30677 & n6564 ;
  assign n6566 = n3329 | n6565 ;
  assign n30678 = ~n6560 ;
  assign n6567 = n30678 & n6566 ;
  assign n6569 = n6559 | n6567 ;
  assign n6570 = n891 & n30463 ;
  assign n6571 = x29 & n6570 ;
  assign n6572 = n2471 & n30463 ;
  assign n6573 = n2788 | n6572 ;
  assign n6574 = n895 & n6573 ;
  assign n6581 = n30463 & n2849 ;
  assign n6582 = n894 & n30155 ;
  assign n6583 = n6581 | n6582 ;
  assign n6584 = n6574 | n6583 ;
  assign n6586 = n6571 | n6584 ;
  assign n6587 = x29 & n6586 ;
  assign n5569 = n895 & n5567 ;
  assign n2793 = n894 & n2639 ;
  assign n2850 = n30155 & n2849 ;
  assign n6588 = n2793 | n2850 ;
  assign n6589 = n30463 & n2861 ;
  assign n6590 = n6588 | n6589 ;
  assign n6591 = n5569 | n6590 ;
  assign n6592 = n6587 | n6591 ;
  assign n5633 = n895 & n5631 ;
  assign n2797 = n894 & n30453 ;
  assign n2863 = n30155 & n2861 ;
  assign n6593 = n2797 | n2863 ;
  assign n6594 = n2639 & n2849 ;
  assign n6595 = n6593 | n6594 ;
  assign n6596 = n5633 | n6595 ;
  assign n6597 = n6592 | n6596 ;
  assign n6598 = n108 & n30463 ;
  assign n30679 = ~n6598 ;
  assign n6599 = n6597 & n30679 ;
  assign n6600 = n6592 & n6596 ;
  assign n6601 = x29 & n6600 ;
  assign n6602 = x29 | n6596 ;
  assign n30680 = ~n6601 ;
  assign n6603 = n30680 & n6602 ;
  assign n30681 = ~n6599 ;
  assign n6604 = n30681 & n6603 ;
  assign n6568 = n6559 & n6567 ;
  assign n30682 = ~n6568 ;
  assign n6605 = n30682 & n6569 ;
  assign n30683 = ~n6604 ;
  assign n6607 = n30683 & n6605 ;
  assign n30684 = ~n6607 ;
  assign n6608 = n6569 & n30684 ;
  assign n30685 = ~n6552 ;
  assign n6609 = n30685 & n6608 ;
  assign n6610 = n6550 | n6609 ;
  assign n6612 = n6541 | n6610 ;
  assign n30686 = ~n6539 ;
  assign n6613 = n30686 & n6612 ;
  assign n6527 = n6519 & n6526 ;
  assign n30687 = ~n6527 ;
  assign n6614 = n30687 & n6528 ;
  assign n30688 = ~n6613 ;
  assign n6616 = n30688 & n6614 ;
  assign n30689 = ~n6616 ;
  assign n6617 = n6528 & n30689 ;
  assign n6619 = n6517 | n6617 ;
  assign n30690 = ~n6516 ;
  assign n6620 = n30690 & n6619 ;
  assign n30691 = ~n6620 ;
  assign n6622 = n6505 & n30691 ;
  assign n30692 = ~n6622 ;
  assign n6623 = n6503 & n30692 ;
  assign n30693 = ~n6623 ;
  assign n6625 = n6492 & n30693 ;
  assign n30694 = ~n6625 ;
  assign n6626 = n6490 & n30694 ;
  assign n6628 = n6479 | n6626 ;
  assign n3795 = n30233 & n3791 ;
  assign n3810 = n30105 & n3802 ;
  assign n3824 = n30196 & n3818 ;
  assign n6629 = n3810 | n3824 ;
  assign n6630 = n209 & n1812 ;
  assign n6631 = n6629 | n6630 ;
  assign n6632 = n3795 | n6631 ;
  assign n30695 = ~n6632 ;
  assign n6633 = x26 & n30695 ;
  assign n6634 = n30019 & n6632 ;
  assign n6635 = n6633 | n6634 ;
  assign n30696 = ~n6479 ;
  assign n6627 = n30696 & n6626 ;
  assign n30697 = ~n6626 ;
  assign n6636 = n6479 & n30697 ;
  assign n6637 = n6627 | n6636 ;
  assign n30698 = ~n6635 ;
  assign n6638 = n30698 & n6637 ;
  assign n30699 = ~n6638 ;
  assign n6639 = n6628 & n30699 ;
  assign n6641 = n6477 | n6639 ;
  assign n4144 = n30238 & n4135 ;
  assign n4178 = n1219 & n4165 ;
  assign n4196 = n1445 & n4185 ;
  assign n6642 = n4178 | n4196 ;
  assign n6643 = n30082 & n4148 ;
  assign n6644 = n6642 | n6643 ;
  assign n6645 = n4144 | n6644 ;
  assign n30700 = ~n6645 ;
  assign n6646 = x23 & n30700 ;
  assign n6647 = n30030 & n6645 ;
  assign n6648 = n6646 | n6647 ;
  assign n6640 = n6477 & n6639 ;
  assign n30701 = ~n6640 ;
  assign n6649 = n30701 & n6641 ;
  assign n30702 = ~n6648 ;
  assign n6650 = n30702 & n6649 ;
  assign n30703 = ~n6650 ;
  assign n6651 = n6641 & n30703 ;
  assign n30704 = ~n6651 ;
  assign n6653 = n6475 & n30704 ;
  assign n4698 = n3787 & n4686 ;
  assign n4714 = n3764 & n4706 ;
  assign n4735 = n1074 & n4726 ;
  assign n6654 = n4714 | n4735 ;
  assign n6655 = n3700 & n4748 ;
  assign n6656 = n6654 | n6655 ;
  assign n6657 = n4698 | n6656 ;
  assign n30705 = ~n6657 ;
  assign n6658 = x20 & n30705 ;
  assign n6659 = n30374 & n6657 ;
  assign n6660 = n6658 | n6659 ;
  assign n30706 = ~n6475 ;
  assign n6652 = n30706 & n6651 ;
  assign n6661 = n6652 | n6653 ;
  assign n6662 = n6660 | n6661 ;
  assign n30707 = ~n6653 ;
  assign n6663 = n30707 & n6662 ;
  assign n6665 = n6473 | n6663 ;
  assign n30708 = ~n6473 ;
  assign n6664 = n30708 & n6663 ;
  assign n30709 = ~n6663 ;
  assign n6666 = n6473 & n30709 ;
  assign n6667 = n6664 | n6666 ;
  assign n4697 = n30263 & n4686 ;
  assign n4712 = n3700 & n4706 ;
  assign n4733 = n3764 & n4726 ;
  assign n6668 = n4712 | n4733 ;
  assign n6669 = n30264 & n4748 ;
  assign n6670 = n6668 | n6669 ;
  assign n6671 = n4697 | n6670 ;
  assign n30710 = ~n6671 ;
  assign n6672 = x20 & n30710 ;
  assign n6673 = n30374 & n6671 ;
  assign n6674 = n6672 | n6673 ;
  assign n30711 = ~n6674 ;
  assign n6675 = n6667 & n30711 ;
  assign n30712 = ~n6675 ;
  assign n6676 = n6665 & n30712 ;
  assign n30713 = ~n6676 ;
  assign n6678 = n6471 & n30713 ;
  assign n30714 = ~n6471 ;
  assign n6677 = n30714 & n6676 ;
  assign n6679 = n6677 | n6678 ;
  assign n5726 = n37300 & n5723 ;
  assign n5177 = n4033 & n5166 ;
  assign n5200 = n30361 & n5191 ;
  assign n6680 = n5177 | n5200 ;
  assign n6681 = n30282 & n5144 ;
  assign n6682 = n6680 | n6681 ;
  assign n6683 = n5726 | n6682 ;
  assign n30715 = ~n6683 ;
  assign n6684 = x17 & n30715 ;
  assign n6685 = n30580 & n6683 ;
  assign n6686 = n6684 | n6685 ;
  assign n6687 = n6679 | n6686 ;
  assign n30716 = ~n6678 ;
  assign n6688 = n30716 & n6687 ;
  assign n6690 = n6469 & n6688 ;
  assign n5953 = n30512 & n5937 ;
  assign n5984 = n30405 & n5970 ;
  assign n6001 = n4811 & n5994 ;
  assign n6691 = n5984 | n6001 ;
  assign n6692 = n5017 & n6018 ;
  assign n6693 = n6691 | n6692 ;
  assign n6694 = n5953 | n6693 ;
  assign n30717 = ~n6694 ;
  assign n6695 = x14 & n30717 ;
  assign n6696 = n30547 & n6694 ;
  assign n6697 = n6695 | n6696 ;
  assign n30718 = ~n6469 ;
  assign n6689 = n30718 & n6688 ;
  assign n30719 = ~n6688 ;
  assign n6698 = n6469 & n30719 ;
  assign n6699 = n6689 | n6698 ;
  assign n6701 = n6697 & n6699 ;
  assign n6702 = n6690 | n6701 ;
  assign n6704 = n6467 | n6702 ;
  assign n30720 = ~n6404 ;
  assign n6407 = n30720 & n6406 ;
  assign n30721 = ~n6406 ;
  assign n6705 = n6404 & n30721 ;
  assign n6706 = n6407 | n6705 ;
  assign n30722 = ~n6702 ;
  assign n6703 = n6467 & n30722 ;
  assign n30723 = ~n6467 ;
  assign n6707 = n30723 & n6702 ;
  assign n6708 = n6703 | n6707 ;
  assign n30724 = ~n6706 ;
  assign n6709 = n30724 & n6708 ;
  assign n30725 = ~n6709 ;
  assign n6711 = n6704 & n30725 ;
  assign n6712 = n6460 & n6711 ;
  assign n30726 = ~n6428 ;
  assign n6713 = n6426 & n30726 ;
  assign n6714 = n6429 | n6713 ;
  assign n6715 = n6460 | n6711 ;
  assign n30727 = ~n6712 ;
  assign n6716 = n30727 & n6715 ;
  assign n6718 = n6714 & n6716 ;
  assign n6719 = n6712 | n6718 ;
  assign n6720 = n6442 | n6719 ;
  assign n6721 = n6442 & n6719 ;
  assign n30728 = ~n6721 ;
  assign n6722 = n6720 & n30728 ;
  assign n30729 = ~n6714 ;
  assign n6717 = n30729 & n6716 ;
  assign n30730 = ~n6716 ;
  assign n6723 = n6714 & n30730 ;
  assign n6724 = n6717 | n6723 ;
  assign n6710 = n6706 & n6708 ;
  assign n6725 = n6706 | n6708 ;
  assign n30731 = ~n6710 ;
  assign n6726 = n30731 & n6725 ;
  assign n30732 = ~n6697 ;
  assign n6700 = n30732 & n6699 ;
  assign n30733 = ~n6699 ;
  assign n6727 = n6697 & n30733 ;
  assign n6728 = n6700 | n6727 ;
  assign n6729 = n6679 & n6686 ;
  assign n30734 = ~n6729 ;
  assign n6730 = n6687 & n30734 ;
  assign n30735 = ~n6667 ;
  assign n6731 = n30735 & n6674 ;
  assign n6732 = n6675 | n6731 ;
  assign n4125 = n37300 & n30286 ;
  assign n5181 = n4093 & n5166 ;
  assign n5201 = n30282 & n5191 ;
  assign n6733 = n5181 | n5201 ;
  assign n6734 = n4033 & n5144 ;
  assign n6735 = n6733 | n6734 ;
  assign n6736 = n4125 | n6735 ;
  assign n30736 = ~n6736 ;
  assign n6737 = x17 & n30736 ;
  assign n6738 = n30580 & n6736 ;
  assign n6739 = n6737 | n6738 ;
  assign n6740 = n6732 | n6739 ;
  assign n6741 = n6732 & n6739 ;
  assign n30737 = ~n6741 ;
  assign n6742 = n6740 & n30737 ;
  assign n6743 = n6660 & n6661 ;
  assign n30738 = ~n6743 ;
  assign n6744 = n6662 & n30738 ;
  assign n30739 = ~n6649 ;
  assign n6745 = n6648 & n30739 ;
  assign n6746 = n6650 | n6745 ;
  assign n4695 = n4420 & n4686 ;
  assign n4716 = n1074 & n4706 ;
  assign n4750 = n3764 & n4748 ;
  assign n6747 = n4716 | n4750 ;
  assign n6748 = n30074 & n4726 ;
  assign n6749 = n6747 | n6748 ;
  assign n6750 = n4695 | n6749 ;
  assign n30740 = ~n6750 ;
  assign n6751 = x20 & n30740 ;
  assign n6752 = n30374 & n6750 ;
  assign n6753 = n6751 | n6752 ;
  assign n6754 = n6746 | n6753 ;
  assign n6755 = n6746 & n6753 ;
  assign n30741 = ~n6755 ;
  assign n6756 = n6754 & n30741 ;
  assign n30742 = ~n6637 ;
  assign n6757 = n6635 & n30742 ;
  assign n6758 = n6638 | n6757 ;
  assign n4140 = n30203 & n4135 ;
  assign n4164 = n1445 & n4148 ;
  assign n4191 = n1556 & n4185 ;
  assign n6759 = n4164 | n4191 ;
  assign n6760 = n30082 & n4165 ;
  assign n6761 = n6759 | n6760 ;
  assign n6762 = n4140 | n6761 ;
  assign n30743 = ~n6762 ;
  assign n6763 = x23 & n30743 ;
  assign n6764 = n30030 & n6762 ;
  assign n6765 = n6763 | n6764 ;
  assign n6766 = n6758 | n6765 ;
  assign n6624 = n6492 & n6623 ;
  assign n6767 = n6492 | n6623 ;
  assign n30744 = ~n6624 ;
  assign n6768 = n30744 & n6767 ;
  assign n4234 = n3791 & n4230 ;
  assign n1889 = n209 & n30108 ;
  assign n3823 = n30105 & n3818 ;
  assign n6769 = n1889 | n3823 ;
  assign n6770 = n1812 & n3802 ;
  assign n6771 = n6769 | n6770 ;
  assign n6772 = n4234 | n6771 ;
  assign n6773 = x26 | n6772 ;
  assign n6774 = x26 & n6772 ;
  assign n30745 = ~n6774 ;
  assign n6775 = n6773 & n30745 ;
  assign n6777 = n6768 | n6775 ;
  assign n30746 = ~n6768 ;
  assign n6776 = n30746 & n6775 ;
  assign n30747 = ~n6775 ;
  assign n6778 = n6768 & n30747 ;
  assign n6779 = n6776 | n6778 ;
  assign n6621 = n6505 & n6620 ;
  assign n6780 = n6505 | n6620 ;
  assign n30748 = ~n6621 ;
  assign n6781 = n30748 & n6780 ;
  assign n3796 = n3592 & n3791 ;
  assign n1962 = n209 & n30114 ;
  assign n3822 = n1812 & n3818 ;
  assign n6782 = n1962 | n3822 ;
  assign n6783 = n30108 & n3802 ;
  assign n6784 = n6782 | n6783 ;
  assign n6785 = n3796 | n6784 ;
  assign n30749 = ~n6785 ;
  assign n6786 = x26 & n30749 ;
  assign n6787 = n30019 & n6785 ;
  assign n6788 = n6786 | n6787 ;
  assign n6789 = n6781 | n6788 ;
  assign n6790 = n6781 & n6788 ;
  assign n30750 = ~n6790 ;
  assign n6791 = n6789 & n30750 ;
  assign n30751 = ~n6517 ;
  assign n6618 = n30751 & n6617 ;
  assign n30752 = ~n6617 ;
  assign n6792 = n6517 & n30752 ;
  assign n6793 = n6618 | n6792 ;
  assign n4380 = n3791 & n30310 ;
  assign n3804 = n30114 & n3802 ;
  assign n3821 = n30108 & n3818 ;
  assign n6794 = n3804 | n3821 ;
  assign n6795 = n209 & n30123 ;
  assign n6796 = n6794 | n6795 ;
  assign n6797 = n4380 | n6796 ;
  assign n6798 = x26 | n6797 ;
  assign n6799 = x26 & n6797 ;
  assign n30753 = ~n6799 ;
  assign n6800 = n6798 & n30753 ;
  assign n30754 = ~n6800 ;
  assign n6802 = n6793 & n30754 ;
  assign n6801 = n6793 & n6800 ;
  assign n6803 = n6793 | n6800 ;
  assign n30755 = ~n6801 ;
  assign n6804 = n30755 & n6803 ;
  assign n6615 = n6613 & n6614 ;
  assign n6805 = n6613 | n6614 ;
  assign n30756 = ~n6615 ;
  assign n6806 = n30756 & n6805 ;
  assign n5254 = n3791 & n5251 ;
  assign n2105 = n209 & n2102 ;
  assign n3820 = n30114 & n3818 ;
  assign n6807 = n2105 | n3820 ;
  assign n6808 = n30123 & n3802 ;
  assign n6809 = n6807 | n6808 ;
  assign n6810 = n5254 | n6809 ;
  assign n6811 = x26 | n6810 ;
  assign n6812 = x26 & n6810 ;
  assign n30757 = ~n6812 ;
  assign n6813 = n6811 & n30757 ;
  assign n6815 = n6806 | n6813 ;
  assign n30758 = ~n6806 ;
  assign n6814 = n30758 & n6813 ;
  assign n30759 = ~n6813 ;
  assign n6816 = n6806 & n30759 ;
  assign n6817 = n6814 | n6816 ;
  assign n30760 = ~n6610 ;
  assign n6611 = n6541 & n30760 ;
  assign n30761 = ~n6541 ;
  assign n6818 = n30761 & n6610 ;
  assign n6819 = n6611 | n6818 ;
  assign n5273 = n3791 & n30440 ;
  assign n2219 = n209 & n2216 ;
  assign n3806 = n2102 & n3802 ;
  assign n6820 = n2219 | n3806 ;
  assign n6821 = n30123 & n3818 ;
  assign n6822 = n6820 | n6821 ;
  assign n6823 = n5273 | n6822 ;
  assign n6824 = x26 | n6823 ;
  assign n6825 = x26 & n6823 ;
  assign n30762 = ~n6825 ;
  assign n6826 = n6824 & n30762 ;
  assign n30763 = ~n6826 ;
  assign n6828 = n6819 & n30763 ;
  assign n30764 = ~n6819 ;
  assign n6827 = n30764 & n6826 ;
  assign n6829 = n6827 | n6828 ;
  assign n30765 = ~n6608 ;
  assign n6830 = n6552 & n30765 ;
  assign n6831 = n6609 | n6830 ;
  assign n4355 = n3791 & n4352 ;
  assign n2299 = n209 & n2295 ;
  assign n3814 = n2216 & n3802 ;
  assign n6832 = n2299 | n3814 ;
  assign n6833 = n2102 & n3818 ;
  assign n6834 = n6832 | n6833 ;
  assign n6835 = n4355 | n6834 ;
  assign n6836 = x26 | n6835 ;
  assign n6837 = x26 & n6835 ;
  assign n30766 = ~n6837 ;
  assign n6838 = n6836 & n30766 ;
  assign n30767 = ~n6838 ;
  assign n6840 = n6831 & n30767 ;
  assign n30768 = ~n6831 ;
  assign n6839 = n30768 & n6838 ;
  assign n6841 = n6839 | n6840 ;
  assign n5338 = n3791 & n30444 ;
  assign n3807 = n2295 & n3802 ;
  assign n3828 = n2216 & n3818 ;
  assign n6842 = n3807 | n3828 ;
  assign n6843 = n209 & n30445 ;
  assign n6844 = n6842 | n6843 ;
  assign n6845 = n5338 | n6844 ;
  assign n6846 = x26 | n6845 ;
  assign n6847 = x26 & n6845 ;
  assign n30769 = ~n6847 ;
  assign n6848 = n6846 & n30769 ;
  assign n6606 = n6604 & n6605 ;
  assign n6849 = n6604 | n6605 ;
  assign n30770 = ~n6606 ;
  assign n6850 = n30770 & n6849 ;
  assign n6852 = n6848 | n6850 ;
  assign n5395 = n3791 & n5392 ;
  assign n2782 = n209 & n30157 ;
  assign n3819 = n2295 & n3818 ;
  assign n6853 = n2782 | n3819 ;
  assign n6854 = n30445 & n3802 ;
  assign n6855 = n6853 | n6854 ;
  assign n6856 = n5395 | n6855 ;
  assign n6857 = x26 | n6856 ;
  assign n6858 = x26 & n6856 ;
  assign n30771 = ~n6858 ;
  assign n6859 = n6857 & n30771 ;
  assign n6860 = n6597 & n6603 ;
  assign n6861 = n30679 & n6860 ;
  assign n30772 = ~n6860 ;
  assign n6862 = n6598 & n30772 ;
  assign n6863 = n6861 | n6862 ;
  assign n6865 = n6859 & n6863 ;
  assign n30773 = ~n6863 ;
  assign n6864 = n6859 & n30773 ;
  assign n30774 = ~n6859 ;
  assign n6866 = n30774 & n6863 ;
  assign n6867 = n6864 | n6866 ;
  assign n6868 = n6587 & n6591 ;
  assign n30775 = ~n6868 ;
  assign n6869 = n6592 & n30775 ;
  assign n5448 = n3791 & n30452 ;
  assign n3816 = n30157 & n3802 ;
  assign n3829 = n30445 & n3818 ;
  assign n6870 = n3816 | n3829 ;
  assign n6871 = n209 & n30453 ;
  assign n6872 = n6870 | n6871 ;
  assign n6873 = n5448 | n6872 ;
  assign n6874 = x26 | n6873 ;
  assign n6875 = x26 & n6873 ;
  assign n30776 = ~n6875 ;
  assign n6876 = n6874 & n30776 ;
  assign n6877 = n6869 & n6876 ;
  assign n6878 = n6869 | n6876 ;
  assign n30777 = ~n6877 ;
  assign n6879 = n30777 & n6878 ;
  assign n30778 = ~n6584 ;
  assign n6585 = n6571 & n30778 ;
  assign n30779 = ~n6571 ;
  assign n6880 = n30779 & n6584 ;
  assign n6881 = n6585 | n6880 ;
  assign n5499 = n3791 & n30458 ;
  assign n2792 = n209 & n2639 ;
  assign n3832 = n30157 & n3818 ;
  assign n6882 = n2792 | n3832 ;
  assign n6883 = n30453 & n3802 ;
  assign n6884 = n6882 | n6883 ;
  assign n6885 = n5499 | n6884 ;
  assign n6886 = x26 | n6885 ;
  assign n6887 = x26 & n6885 ;
  assign n30780 = ~n6887 ;
  assign n6888 = n6886 & n30780 ;
  assign n6889 = n6881 & n6888 ;
  assign n6890 = n260 & n30463 ;
  assign n6891 = x26 & n6890 ;
  assign n6575 = n3791 & n6573 ;
  assign n6892 = n30463 & n3802 ;
  assign n6893 = n30155 & n3818 ;
  assign n6894 = n6892 | n6893 ;
  assign n6895 = n6575 | n6894 ;
  assign n6897 = n6891 | n6895 ;
  assign n6898 = x26 & n6897 ;
  assign n5570 = n3791 & n5567 ;
  assign n2568 = n209 & n30463 ;
  assign n3833 = n2639 & n3818 ;
  assign n6899 = n2568 | n3833 ;
  assign n6900 = n30155 & n3802 ;
  assign n6901 = n6899 | n6900 ;
  assign n6902 = n5570 | n6901 ;
  assign n6903 = n6898 | n6902 ;
  assign n30781 = ~n6903 ;
  assign n6904 = x26 & n30781 ;
  assign n6906 = n6570 | n6904 ;
  assign n5635 = n3791 & n5631 ;
  assign n3803 = n2639 & n3802 ;
  assign n3834 = n30453 & n3818 ;
  assign n6907 = n3803 | n3834 ;
  assign n6908 = n209 & n30155 ;
  assign n6909 = n6907 | n6908 ;
  assign n6910 = n5635 | n6909 ;
  assign n30782 = ~n6910 ;
  assign n6911 = x26 & n30782 ;
  assign n6912 = n30019 & n6910 ;
  assign n6913 = n6911 | n6912 ;
  assign n6914 = n6906 & n6913 ;
  assign n6915 = n6881 | n6888 ;
  assign n30783 = ~n6889 ;
  assign n6916 = n30783 & n6915 ;
  assign n6917 = n6914 & n6916 ;
  assign n6918 = n6889 | n6917 ;
  assign n6920 = n6879 & n6918 ;
  assign n6921 = n6877 | n6920 ;
  assign n6923 = n6867 & n6921 ;
  assign n6924 = n6865 | n6923 ;
  assign n30784 = ~n6850 ;
  assign n6851 = n6848 & n30784 ;
  assign n30785 = ~n6848 ;
  assign n6925 = n30785 & n6850 ;
  assign n6926 = n6851 | n6925 ;
  assign n30786 = ~n6924 ;
  assign n6927 = n30786 & n6926 ;
  assign n30787 = ~n6927 ;
  assign n6928 = n6852 & n30787 ;
  assign n6930 = n6841 | n6928 ;
  assign n30788 = ~n6840 ;
  assign n6931 = n30788 & n6930 ;
  assign n6933 = n6829 | n6931 ;
  assign n30789 = ~n6828 ;
  assign n6934 = n30789 & n6933 ;
  assign n30790 = ~n6934 ;
  assign n6936 = n6817 & n30790 ;
  assign n30791 = ~n6936 ;
  assign n6937 = n6815 & n30791 ;
  assign n6939 = n6804 | n6937 ;
  assign n30792 = ~n6802 ;
  assign n6940 = n30792 & n6939 ;
  assign n30793 = ~n6940 ;
  assign n6942 = n6791 & n30793 ;
  assign n30794 = ~n6942 ;
  assign n6943 = n6789 & n30794 ;
  assign n30795 = ~n6943 ;
  assign n6945 = n6779 & n30795 ;
  assign n30796 = ~n6945 ;
  assign n6946 = n6777 & n30796 ;
  assign n6947 = n6758 & n6765 ;
  assign n30797 = ~n6947 ;
  assign n6948 = n6766 & n30797 ;
  assign n30798 = ~n6946 ;
  assign n6950 = n30798 & n6948 ;
  assign n30799 = ~n6950 ;
  assign n6951 = n6766 & n30799 ;
  assign n30800 = ~n6951 ;
  assign n6953 = n6756 & n30800 ;
  assign n30801 = ~n6953 ;
  assign n6954 = n6754 & n30801 ;
  assign n30802 = ~n6954 ;
  assign n6956 = n6744 & n30802 ;
  assign n4444 = n37300 & n4442 ;
  assign n5156 = n4093 & n5144 ;
  assign n5198 = n4033 & n5191 ;
  assign n6957 = n5156 | n5198 ;
  assign n6958 = n30264 & n5166 ;
  assign n6959 = n6957 | n6958 ;
  assign n6960 = n4444 | n6959 ;
  assign n30803 = ~n6960 ;
  assign n6961 = x17 & n30803 ;
  assign n6962 = n30580 & n6960 ;
  assign n6963 = n6961 | n6962 ;
  assign n30804 = ~n6744 ;
  assign n6955 = n30804 & n6954 ;
  assign n6964 = n6955 | n6956 ;
  assign n6965 = n6963 | n6964 ;
  assign n30805 = ~n6956 ;
  assign n6966 = n30805 & n6965 ;
  assign n30806 = ~n6966 ;
  assign n6968 = n6742 & n30806 ;
  assign n30807 = ~n6968 ;
  assign n6969 = n6740 & n30807 ;
  assign n30808 = ~n6969 ;
  assign n6971 = n6730 & n30808 ;
  assign n6142 = n5937 & n30578 ;
  assign n5981 = n4811 & n5970 ;
  assign n6005 = n4664 & n5994 ;
  assign n6972 = n5981 | n6005 ;
  assign n6973 = n30405 & n6018 ;
  assign n6974 = n6972 | n6973 ;
  assign n6975 = n6142 | n6974 ;
  assign n30809 = ~n6975 ;
  assign n6976 = x14 & n30809 ;
  assign n6977 = n30547 & n6975 ;
  assign n6978 = n6976 | n6977 ;
  assign n6970 = n6730 & n6969 ;
  assign n6979 = n6730 | n6969 ;
  assign n30810 = ~n6970 ;
  assign n6980 = n30810 & n6979 ;
  assign n6981 = n6978 | n6980 ;
  assign n30811 = ~n6971 ;
  assign n6982 = n30811 & n6981 ;
  assign n6984 = n6728 | n6982 ;
  assign n6302 = n30587 & n6272 ;
  assign n30812 = ~n6216 ;
  assign n6217 = n6188 & n30812 ;
  assign n6233 = n30535 & n6217 ;
  assign n6257 = n30415 & n6244 ;
  assign n6985 = n6233 | n6257 ;
  assign n6986 = n30530 & n6190 ;
  assign n6987 = n6985 | n6986 ;
  assign n6988 = n6302 | n6987 ;
  assign n6989 = x11 | n6988 ;
  assign n6990 = x11 & n6988 ;
  assign n30813 = ~n6990 ;
  assign n6991 = n6989 & n30813 ;
  assign n6983 = n6728 & n6982 ;
  assign n30814 = ~n6983 ;
  assign n6992 = n30814 & n6984 ;
  assign n30815 = ~n6991 ;
  assign n6994 = n30815 & n6992 ;
  assign n30816 = ~n6994 ;
  assign n6995 = n6984 & n30816 ;
  assign n6997 = n6726 & n6995 ;
  assign n6292 = n30540 & n6272 ;
  assign n6212 = n30535 & n6190 ;
  assign n6240 = n30545 & n6217 ;
  assign n6998 = n6212 | n6240 ;
  assign n6999 = n30530 & n6244 ;
  assign n7000 = n6998 | n6999 ;
  assign n7001 = n6292 | n7000 ;
  assign n7002 = x11 | n7001 ;
  assign n7003 = x11 & n7001 ;
  assign n30817 = ~n7003 ;
  assign n7004 = n7002 & n30817 ;
  assign n30818 = ~n6726 ;
  assign n6996 = n30818 & n6995 ;
  assign n30819 = ~n6995 ;
  assign n7005 = n6726 & n30819 ;
  assign n7006 = n6996 | n7005 ;
  assign n7007 = n7004 & n7006 ;
  assign n7008 = n6997 | n7007 ;
  assign n7010 = n6724 | n7008 ;
  assign n30820 = ~n7008 ;
  assign n7009 = n6724 & n30820 ;
  assign n30821 = ~n6724 ;
  assign n7011 = n30821 & n7008 ;
  assign n7012 = n7009 | n7011 ;
  assign n7013 = n7004 | n7006 ;
  assign n30822 = ~n7007 ;
  assign n7014 = n30822 & n7013 ;
  assign n37290 = x7 & x8 ;
  assign n7015 = x7 | x8 ;
  assign n30823 = ~n37290 ;
  assign n7016 = n30823 & n7015 ;
  assign n30824 = ~n70 ;
  assign n7041 = n30824 & n7016 ;
  assign n7068 = n67 & n7016 ;
  assign n7086 = n30597 & n7068 ;
  assign n7106 = n7041 | n7086 ;
  assign n7107 = n30545 & n7106 ;
  assign n7108 = x8 & n7107 ;
  assign n7109 = x8 | n7107 ;
  assign n30825 = ~n7108 ;
  assign n7110 = n30825 & n7109 ;
  assign n7111 = n6978 & n6980 ;
  assign n30826 = ~n7111 ;
  assign n7112 = n6981 & n30826 ;
  assign n30827 = ~n6742 ;
  assign n6967 = n30827 & n6966 ;
  assign n7113 = n6967 | n6968 ;
  assign n5940 = n4674 & n5937 ;
  assign n5980 = n30361 & n5970 ;
  assign n6002 = n30282 & n5994 ;
  assign n7114 = n5980 | n6002 ;
  assign n7115 = n4664 & n6018 ;
  assign n7116 = n7114 | n7115 ;
  assign n7117 = n5940 | n7116 ;
  assign n30828 = ~n7117 ;
  assign n7118 = x14 & n30828 ;
  assign n7119 = n30547 & n7117 ;
  assign n7120 = n7118 | n7119 ;
  assign n7121 = n6963 & n6964 ;
  assign n30829 = ~n7121 ;
  assign n7122 = n6965 & n30829 ;
  assign n30830 = ~n7122 ;
  assign n7124 = n7120 & n30830 ;
  assign n30831 = ~n7120 ;
  assign n7123 = n30831 & n7122 ;
  assign n7125 = n7123 | n7124 ;
  assign n6952 = n6756 & n6951 ;
  assign n7126 = n6756 | n6951 ;
  assign n30832 = ~n6952 ;
  assign n7127 = n30832 & n7126 ;
  assign n4511 = n37300 & n30349 ;
  assign n5175 = n3700 & n5166 ;
  assign n5202 = n4093 & n5191 ;
  assign n7128 = n5175 | n5202 ;
  assign n7129 = n30264 & n5144 ;
  assign n7130 = n7128 | n7129 ;
  assign n7131 = n4511 | n7130 ;
  assign n7132 = x17 | n7131 ;
  assign n7133 = x17 & n7131 ;
  assign n30833 = ~n7133 ;
  assign n7134 = n7132 & n30833 ;
  assign n7136 = n7127 | n7134 ;
  assign n6949 = n6946 & n6948 ;
  assign n7137 = n6946 | n6948 ;
  assign n30834 = ~n6949 ;
  assign n7138 = n30834 & n7137 ;
  assign n4694 = n30173 & n4686 ;
  assign n4732 = n1219 & n4726 ;
  assign n4754 = n1074 & n4748 ;
  assign n7139 = n4732 | n4754 ;
  assign n7140 = n30074 & n4706 ;
  assign n7141 = n7139 | n7140 ;
  assign n7142 = n4694 | n7141 ;
  assign n7143 = x20 | n7142 ;
  assign n7144 = x20 & n7142 ;
  assign n30835 = ~n7144 ;
  assign n7145 = n7143 & n30835 ;
  assign n7147 = n7138 | n7145 ;
  assign n30836 = ~n7138 ;
  assign n7146 = n30836 & n7145 ;
  assign n30837 = ~n7145 ;
  assign n7148 = n7138 & n30837 ;
  assign n7149 = n7146 | n7148 ;
  assign n4139 = n30209 & n4135 ;
  assign n4156 = n1556 & n4148 ;
  assign n4171 = n1445 & n4165 ;
  assign n7150 = n4156 | n4171 ;
  assign n7151 = n30196 & n4185 ;
  assign n7152 = n7150 | n7151 ;
  assign n7153 = n4139 | n7152 ;
  assign n30838 = ~n7153 ;
  assign n7154 = x23 & n30838 ;
  assign n7155 = n30030 & n7153 ;
  assign n7156 = n7154 | n7155 ;
  assign n6941 = n6791 & n6940 ;
  assign n7157 = n6791 | n6940 ;
  assign n30839 = ~n6941 ;
  assign n7158 = n30839 & n7157 ;
  assign n4138 = n3307 & n4135 ;
  assign n4175 = n1556 & n4165 ;
  assign n4187 = n30105 & n4185 ;
  assign n7159 = n4175 | n4187 ;
  assign n7160 = n30196 & n4148 ;
  assign n7161 = n7159 | n7160 ;
  assign n7162 = n4138 | n7161 ;
  assign n30840 = ~n7162 ;
  assign n7163 = x23 & n30840 ;
  assign n7164 = n30030 & n7162 ;
  assign n7165 = n7163 | n7164 ;
  assign n7167 = n7158 & n7165 ;
  assign n30841 = ~n7165 ;
  assign n7166 = n7158 & n30841 ;
  assign n30842 = ~n7158 ;
  assign n7168 = n30842 & n7165 ;
  assign n7169 = n7166 | n7168 ;
  assign n6938 = n6804 & n6937 ;
  assign n30843 = ~n6938 ;
  assign n7170 = n30843 & n6939 ;
  assign n4145 = n30233 & n4135 ;
  assign n4157 = n30105 & n4148 ;
  assign n4189 = n1812 & n4185 ;
  assign n7171 = n4157 | n4189 ;
  assign n7172 = n30196 & n4165 ;
  assign n7173 = n7171 | n7172 ;
  assign n7174 = n4145 | n7173 ;
  assign n30844 = ~n7174 ;
  assign n7175 = x23 & n30844 ;
  assign n7176 = n30030 & n7174 ;
  assign n7177 = n7175 | n7176 ;
  assign n30845 = ~n7177 ;
  assign n7178 = n7170 & n30845 ;
  assign n6935 = n6817 & n6934 ;
  assign n7179 = n6817 | n6934 ;
  assign n30846 = ~n6935 ;
  assign n7180 = n30846 & n7179 ;
  assign n4233 = n4135 & n4230 ;
  assign n4163 = n1812 & n4148 ;
  assign n4168 = n30105 & n4165 ;
  assign n7181 = n4163 | n4168 ;
  assign n7182 = n30108 & n4185 ;
  assign n7183 = n7181 | n7182 ;
  assign n7184 = n4233 | n7183 ;
  assign n7185 = x23 | n7184 ;
  assign n7186 = x23 & n7184 ;
  assign n30847 = ~n7186 ;
  assign n7187 = n7185 & n30847 ;
  assign n7189 = n7180 | n7187 ;
  assign n30848 = ~n7180 ;
  assign n7188 = n30848 & n7187 ;
  assign n30849 = ~n7187 ;
  assign n7190 = n7180 & n30849 ;
  assign n7191 = n7188 | n7190 ;
  assign n30850 = ~n6829 ;
  assign n6932 = n30850 & n6931 ;
  assign n30851 = ~n6931 ;
  assign n7192 = n6829 & n30851 ;
  assign n7193 = n6932 | n7192 ;
  assign n4136 = n3592 & n4135 ;
  assign n4167 = n1812 & n4165 ;
  assign n4199 = n30114 & n4185 ;
  assign n7194 = n4167 | n4199 ;
  assign n7195 = n30108 & n4148 ;
  assign n7196 = n7194 | n7195 ;
  assign n7197 = n4136 | n7196 ;
  assign n30852 = ~n7197 ;
  assign n7198 = x23 & n30852 ;
  assign n7199 = n30030 & n7197 ;
  assign n7200 = n7198 | n7199 ;
  assign n30853 = ~n7200 ;
  assign n7202 = n7193 & n30853 ;
  assign n7201 = n7193 | n7200 ;
  assign n7203 = n7193 & n7200 ;
  assign n30854 = ~n7203 ;
  assign n7204 = n7201 & n30854 ;
  assign n30855 = ~n6841 ;
  assign n6929 = n30855 & n6928 ;
  assign n30856 = ~n6928 ;
  assign n7205 = n6841 & n30856 ;
  assign n7206 = n6929 | n7205 ;
  assign n4381 = n4135 & n30310 ;
  assign n4150 = n30114 & n4148 ;
  assign n4198 = n30123 & n4185 ;
  assign n7207 = n4150 | n4198 ;
  assign n7208 = n30108 & n4165 ;
  assign n7209 = n7207 | n7208 ;
  assign n7210 = n4381 | n7209 ;
  assign n30857 = ~n7210 ;
  assign n7211 = x23 & n30857 ;
  assign n7212 = n30030 & n7210 ;
  assign n7213 = n7211 | n7212 ;
  assign n30858 = ~n7213 ;
  assign n7214 = n7206 & n30858 ;
  assign n30859 = ~n7206 ;
  assign n7215 = n30859 & n7213 ;
  assign n7216 = n7214 | n7215 ;
  assign n30860 = ~n6926 ;
  assign n7217 = n6924 & n30860 ;
  assign n7218 = n6927 | n7217 ;
  assign n5255 = n4135 & n5251 ;
  assign n4160 = n30123 & n4148 ;
  assign n4166 = n30114 & n4165 ;
  assign n7219 = n4160 | n4166 ;
  assign n7220 = n2102 & n4185 ;
  assign n7221 = n7219 | n7220 ;
  assign n7222 = n5255 | n7221 ;
  assign n30861 = ~n7222 ;
  assign n7223 = x23 & n30861 ;
  assign n7224 = n30030 & n7222 ;
  assign n7225 = n7223 | n7224 ;
  assign n7226 = n7218 | n7225 ;
  assign n7227 = n7218 & n7225 ;
  assign n30862 = ~n7227 ;
  assign n7228 = n7226 & n30862 ;
  assign n5274 = n4135 & n30440 ;
  assign n4151 = n2102 & n4148 ;
  assign n4190 = n2216 & n4185 ;
  assign n7229 = n4151 | n4190 ;
  assign n7230 = n30123 & n4165 ;
  assign n7231 = n7229 | n7230 ;
  assign n7232 = n5274 | n7231 ;
  assign n7233 = x23 | n7232 ;
  assign n7234 = x23 & n7232 ;
  assign n30863 = ~n7234 ;
  assign n7235 = n7233 & n30863 ;
  assign n30864 = ~n6918 ;
  assign n6919 = n6879 & n30864 ;
  assign n30865 = ~n6879 ;
  assign n7236 = n30865 & n6918 ;
  assign n7237 = n6919 | n7236 ;
  assign n4356 = n4135 & n4352 ;
  assign n4159 = n2216 & n4148 ;
  assign n4201 = n2295 & n4185 ;
  assign n7238 = n4159 | n4201 ;
  assign n7239 = n2102 & n4165 ;
  assign n7240 = n7238 | n7239 ;
  assign n7241 = n4356 | n7240 ;
  assign n7242 = x23 | n7241 ;
  assign n7243 = x23 & n7241 ;
  assign n30866 = ~n7243 ;
  assign n7244 = n7242 & n30866 ;
  assign n7246 = n7237 | n7244 ;
  assign n30867 = ~n7237 ;
  assign n7245 = n30867 & n7244 ;
  assign n30868 = ~n7244 ;
  assign n7247 = n7237 & n30868 ;
  assign n7248 = n7245 | n7247 ;
  assign n7249 = n6914 | n6916 ;
  assign n30869 = ~n6917 ;
  assign n7250 = n30869 & n7249 ;
  assign n5339 = n4135 & n30444 ;
  assign n4161 = n2295 & n4148 ;
  assign n4169 = n2216 & n4165 ;
  assign n7251 = n4161 | n4169 ;
  assign n7252 = n30445 & n4185 ;
  assign n7253 = n7251 | n7252 ;
  assign n7254 = n5339 | n7253 ;
  assign n7255 = x23 | n7254 ;
  assign n7256 = x23 & n7254 ;
  assign n30870 = ~n7256 ;
  assign n7257 = n7255 & n30870 ;
  assign n7259 = n7250 | n7257 ;
  assign n7258 = n7250 & n7257 ;
  assign n30871 = ~n7258 ;
  assign n7260 = n30871 & n7259 ;
  assign n30872 = ~n6570 ;
  assign n6905 = n30872 & n6904 ;
  assign n30873 = ~n6904 ;
  assign n7261 = n6570 & n30873 ;
  assign n7262 = n6905 | n7261 ;
  assign n30874 = ~n6913 ;
  assign n7263 = n30874 & n7262 ;
  assign n30875 = ~n7262 ;
  assign n7264 = n6913 & n30875 ;
  assign n7265 = n7263 | n7264 ;
  assign n5396 = n4135 & n5392 ;
  assign n4172 = n2295 & n4165 ;
  assign n4202 = n30157 & n4185 ;
  assign n7266 = n4172 | n4202 ;
  assign n7267 = n30445 & n4148 ;
  assign n7268 = n7266 | n7267 ;
  assign n7269 = n5396 | n7268 ;
  assign n7270 = x23 | n7269 ;
  assign n7271 = x23 & n7269 ;
  assign n30876 = ~n7271 ;
  assign n7272 = n7270 & n30876 ;
  assign n7273 = n7265 & n7272 ;
  assign n7274 = n6898 & n6902 ;
  assign n30877 = ~n7274 ;
  assign n7275 = n6903 & n30877 ;
  assign n5450 = n4135 & n30452 ;
  assign n4162 = n30157 & n4148 ;
  assign n4181 = n30445 & n4165 ;
  assign n7276 = n4162 | n4181 ;
  assign n7277 = n30453 & n4185 ;
  assign n7278 = n7276 | n7277 ;
  assign n7279 = n5450 | n7278 ;
  assign n30878 = ~n7279 ;
  assign n7280 = x23 & n30878 ;
  assign n7281 = n30030 & n7279 ;
  assign n7282 = n7280 | n7281 ;
  assign n7284 = n7275 | n7282 ;
  assign n30879 = ~n7282 ;
  assign n7283 = n7275 & n30879 ;
  assign n30880 = ~n7275 ;
  assign n7285 = n30880 & n7282 ;
  assign n7286 = n7283 | n7285 ;
  assign n7287 = n30463 & n4132 ;
  assign n7288 = x23 & n7287 ;
  assign n6576 = n4135 & n6573 ;
  assign n7289 = n30463 & n4148 ;
  assign n7290 = n30155 & n4165 ;
  assign n7291 = n7289 | n7290 ;
  assign n7292 = n6576 | n7291 ;
  assign n7294 = n7288 | n7292 ;
  assign n7295 = x23 & n7294 ;
  assign n5571 = n4135 & n5567 ;
  assign n4154 = n30155 & n4148 ;
  assign n4180 = n2639 & n4165 ;
  assign n7296 = n4154 | n4180 ;
  assign n7297 = n30463 & n4185 ;
  assign n7298 = n7296 | n7297 ;
  assign n7299 = n5571 | n7298 ;
  assign n7300 = n7295 | n7299 ;
  assign n30881 = ~n7300 ;
  assign n7301 = x23 & n30881 ;
  assign n7303 = n6890 | n7301 ;
  assign n5636 = n4135 & n5631 ;
  assign n4182 = n30453 & n4165 ;
  assign n4188 = n30155 & n4185 ;
  assign n7304 = n4182 | n4188 ;
  assign n7305 = n2639 & n4148 ;
  assign n7306 = n7304 | n7305 ;
  assign n7307 = n5636 | n7306 ;
  assign n30882 = ~n7307 ;
  assign n7308 = x23 & n30882 ;
  assign n7309 = n30030 & n7307 ;
  assign n7310 = n7308 | n7309 ;
  assign n7311 = n7303 & n7310 ;
  assign n30883 = ~n6895 ;
  assign n6896 = n6891 & n30883 ;
  assign n30884 = ~n6891 ;
  assign n7312 = n30884 & n6895 ;
  assign n7313 = n6896 | n7312 ;
  assign n7314 = n7311 & n7313 ;
  assign n5500 = n4135 & n30458 ;
  assign n4177 = n30157 & n4165 ;
  assign n4203 = n2639 & n4185 ;
  assign n7315 = n4177 | n4203 ;
  assign n7316 = n30453 & n4148 ;
  assign n7317 = n7315 | n7316 ;
  assign n7318 = n5500 | n7317 ;
  assign n30885 = ~n7318 ;
  assign n7319 = x23 & n30885 ;
  assign n7320 = n30030 & n7318 ;
  assign n7321 = n7319 | n7320 ;
  assign n7322 = n7311 | n7313 ;
  assign n30886 = ~n7314 ;
  assign n7323 = n30886 & n7322 ;
  assign n7325 = n7321 & n7323 ;
  assign n7326 = n7314 | n7325 ;
  assign n30887 = ~n7326 ;
  assign n7327 = n7286 & n30887 ;
  assign n30888 = ~n7327 ;
  assign n7329 = n7284 & n30888 ;
  assign n7330 = n7265 | n7272 ;
  assign n30889 = ~n7273 ;
  assign n7331 = n30889 & n7330 ;
  assign n7332 = n7329 & n7331 ;
  assign n7333 = n7273 | n7332 ;
  assign n30890 = ~n7333 ;
  assign n7334 = n7260 & n30890 ;
  assign n30891 = ~n7334 ;
  assign n7336 = n7259 & n30891 ;
  assign n30892 = ~n7336 ;
  assign n7338 = n7248 & n30892 ;
  assign n30893 = ~n7338 ;
  assign n7339 = n7246 & n30893 ;
  assign n7341 = n7235 | n7339 ;
  assign n30894 = ~n6921 ;
  assign n6922 = n6867 & n30894 ;
  assign n30895 = ~n6867 ;
  assign n7342 = n30895 & n6921 ;
  assign n7343 = n6922 | n7342 ;
  assign n7340 = n7235 & n7339 ;
  assign n30896 = ~n7340 ;
  assign n7344 = n30896 & n7341 ;
  assign n30897 = ~n7343 ;
  assign n7345 = n30897 & n7344 ;
  assign n30898 = ~n7345 ;
  assign n7346 = n7341 & n30898 ;
  assign n30899 = ~n7346 ;
  assign n7348 = n7228 & n30899 ;
  assign n30900 = ~n7348 ;
  assign n7349 = n7226 & n30900 ;
  assign n7351 = n7216 | n7349 ;
  assign n30901 = ~n7214 ;
  assign n7352 = n30901 & n7351 ;
  assign n7354 = n7204 | n7352 ;
  assign n30902 = ~n7202 ;
  assign n7355 = n30902 & n7354 ;
  assign n30903 = ~n7355 ;
  assign n7357 = n7191 & n30903 ;
  assign n30904 = ~n7357 ;
  assign n7358 = n7189 & n30904 ;
  assign n30905 = ~n7170 ;
  assign n7359 = n30905 & n7177 ;
  assign n7360 = n7178 | n7359 ;
  assign n7361 = n7358 | n7360 ;
  assign n30906 = ~n7178 ;
  assign n7362 = n30906 & n7361 ;
  assign n7363 = n7169 & n7362 ;
  assign n7364 = n7167 | n7363 ;
  assign n7366 = n7156 & n7364 ;
  assign n6944 = n6779 & n6943 ;
  assign n7367 = n6779 | n6943 ;
  assign n30907 = ~n6944 ;
  assign n7368 = n30907 & n7367 ;
  assign n7365 = n7156 | n7364 ;
  assign n30908 = ~n7366 ;
  assign n7369 = n7365 & n30908 ;
  assign n7370 = n7368 & n7369 ;
  assign n7371 = n7366 | n7370 ;
  assign n30909 = ~n7371 ;
  assign n7372 = n7149 & n30909 ;
  assign n30910 = ~n7372 ;
  assign n7373 = n7147 & n30910 ;
  assign n7135 = n7127 & n7134 ;
  assign n30911 = ~n7135 ;
  assign n7374 = n30911 & n7136 ;
  assign n30912 = ~n7373 ;
  assign n7376 = n30912 & n7374 ;
  assign n30913 = ~n7376 ;
  assign n7377 = n7136 & n30913 ;
  assign n30914 = ~n7125 ;
  assign n7378 = n30914 & n7377 ;
  assign n7379 = n7124 | n7378 ;
  assign n7380 = n7113 | n7379 ;
  assign n5949 = n30385 & n5937 ;
  assign n5999 = n30361 & n5994 ;
  assign n6036 = n4811 & n6018 ;
  assign n7381 = n5999 | n6036 ;
  assign n7382 = n4664 & n5970 ;
  assign n7383 = n7381 | n7382 ;
  assign n7384 = n5949 | n7383 ;
  assign n30915 = ~n7384 ;
  assign n7385 = x14 & n30915 ;
  assign n7386 = n30547 & n7384 ;
  assign n7387 = n7385 | n7386 ;
  assign n7388 = n7113 & n7379 ;
  assign n30916 = ~n7388 ;
  assign n7389 = n7380 & n30916 ;
  assign n30917 = ~n7387 ;
  assign n7390 = n30917 & n7389 ;
  assign n30918 = ~n7390 ;
  assign n7391 = n7380 & n30918 ;
  assign n30919 = ~n7391 ;
  assign n7393 = n7112 & n30919 ;
  assign n6414 = n6272 & n6411 ;
  assign n6205 = n30415 & n6190 ;
  assign n6246 = n5017 & n6244 ;
  assign n7394 = n6205 | n6246 ;
  assign n7395 = n30530 & n6217 ;
  assign n7396 = n7394 | n7395 ;
  assign n7397 = n6414 | n7396 ;
  assign n30920 = ~n7397 ;
  assign n7398 = x11 & n30920 ;
  assign n7399 = n30180 & n7397 ;
  assign n7400 = n7398 | n7399 ;
  assign n7392 = n7112 & n7391 ;
  assign n7401 = n7112 | n7391 ;
  assign n30921 = ~n7392 ;
  assign n7402 = n30921 & n7401 ;
  assign n7403 = n7400 | n7402 ;
  assign n30922 = ~n7393 ;
  assign n7404 = n30922 & n7403 ;
  assign n7405 = n7110 & n7404 ;
  assign n6993 = n6991 & n6992 ;
  assign n7406 = n6991 | n6992 ;
  assign n30923 = ~n6993 ;
  assign n7407 = n30923 & n7406 ;
  assign n7408 = n7110 | n7404 ;
  assign n30924 = ~n7405 ;
  assign n7409 = n30924 & n7408 ;
  assign n7411 = n7407 & n7409 ;
  assign n7412 = n7405 | n7411 ;
  assign n7414 = n7014 | n7412 ;
  assign n30925 = ~n7412 ;
  assign n7413 = n7014 & n30925 ;
  assign n30926 = ~n7014 ;
  assign n7415 = n30926 & n7412 ;
  assign n7416 = n7413 | n7415 ;
  assign n30927 = ~n7407 ;
  assign n7410 = n30927 & n7409 ;
  assign n30928 = ~n7409 ;
  assign n7417 = n7407 & n30928 ;
  assign n7418 = n7410 | n7417 ;
  assign n7419 = n7400 & n7402 ;
  assign n30929 = ~n7419 ;
  assign n7420 = n7403 & n30929 ;
  assign n7088 = n6445 & n7068 ;
  assign n7421 = n69 & n30545 ;
  assign n7422 = n30535 & n7041 ;
  assign n7423 = n7421 | n7422 ;
  assign n7424 = n7088 | n7423 ;
  assign n7425 = x8 | n7424 ;
  assign n7426 = x8 & n7424 ;
  assign n30930 = ~n7426 ;
  assign n7427 = n7425 & n30930 ;
  assign n30931 = ~n7427 ;
  assign n7429 = n7420 & n30931 ;
  assign n7428 = n7420 & n7427 ;
  assign n7430 = n7420 | n7427 ;
  assign n30932 = ~n7428 ;
  assign n7431 = n30932 & n7430 ;
  assign n30933 = ~n7389 ;
  assign n7432 = n7387 & n30933 ;
  assign n7433 = n7390 | n7432 ;
  assign n6293 = n30410 & n6272 ;
  assign n6234 = n30415 & n6217 ;
  assign n6256 = n30405 & n6244 ;
  assign n7434 = n6234 | n6256 ;
  assign n7435 = n5017 & n6190 ;
  assign n7436 = n7434 | n7435 ;
  assign n7437 = n6293 | n7436 ;
  assign n7438 = x11 | n7437 ;
  assign n7439 = x11 & n7437 ;
  assign n30934 = ~n7439 ;
  assign n7440 = n7438 & n30934 ;
  assign n7442 = n7433 | n7440 ;
  assign n30935 = ~n7433 ;
  assign n7441 = n30935 & n7440 ;
  assign n30936 = ~n7440 ;
  assign n7443 = n7433 & n30936 ;
  assign n7444 = n7441 | n7443 ;
  assign n30937 = ~n7377 ;
  assign n7445 = n7125 & n30937 ;
  assign n7446 = n7378 | n7445 ;
  assign n7375 = n7373 & n7374 ;
  assign n7447 = n7373 | n7374 ;
  assign n30938 = ~n7375 ;
  assign n7448 = n30938 & n7447 ;
  assign n5947 = n5723 & n5937 ;
  assign n5979 = n30282 & n5970 ;
  assign n6032 = n30361 & n6018 ;
  assign n7449 = n5979 | n6032 ;
  assign n7450 = n4033 & n5994 ;
  assign n7451 = n7449 | n7450 ;
  assign n7452 = n5947 | n7451 ;
  assign n7453 = x14 | n7452 ;
  assign n7454 = x14 & n7452 ;
  assign n30939 = ~n7454 ;
  assign n7455 = n7453 & n30939 ;
  assign n7457 = n7448 | n7455 ;
  assign n30940 = ~n7149 ;
  assign n7458 = n30940 & n7371 ;
  assign n7459 = n7372 | n7458 ;
  assign n7460 = n7368 | n7369 ;
  assign n30941 = ~n7370 ;
  assign n7461 = n30941 & n7460 ;
  assign n7462 = n7169 | n7362 ;
  assign n30942 = ~n7363 ;
  assign n7463 = n30942 & n7462 ;
  assign n4702 = n30238 & n4686 ;
  assign n4717 = n30082 & n4706 ;
  assign n4734 = n1445 & n4726 ;
  assign n7464 = n4717 | n4734 ;
  assign n7465 = n1219 & n4748 ;
  assign n7466 = n7464 | n7465 ;
  assign n7467 = n4702 | n7466 ;
  assign n7468 = x20 | n7467 ;
  assign n7469 = x20 & n7467 ;
  assign n30943 = ~n7469 ;
  assign n7470 = n7468 & n30943 ;
  assign n7472 = n7463 | n7470 ;
  assign n30944 = ~n7463 ;
  assign n7471 = n30944 & n7470 ;
  assign n30945 = ~n7470 ;
  assign n7473 = n7463 & n30945 ;
  assign n7474 = n7471 | n7473 ;
  assign n7475 = n7358 & n7360 ;
  assign n30946 = ~n7475 ;
  assign n7476 = n7361 & n30946 ;
  assign n4696 = n30203 & n4686 ;
  assign n4709 = n1445 & n4706 ;
  assign n4731 = n1556 & n4726 ;
  assign n7477 = n4709 | n4731 ;
  assign n7478 = n30082 & n4748 ;
  assign n7479 = n7477 | n7478 ;
  assign n7480 = n4696 | n7479 ;
  assign n30947 = ~n7480 ;
  assign n7481 = x20 & n30947 ;
  assign n7482 = n30374 & n7480 ;
  assign n7483 = n7481 | n7482 ;
  assign n30948 = ~n7483 ;
  assign n7484 = n7476 & n30948 ;
  assign n30949 = ~n7476 ;
  assign n7485 = n30949 & n7483 ;
  assign n7486 = n7484 | n7485 ;
  assign n30950 = ~n7191 ;
  assign n7356 = n30950 & n7355 ;
  assign n7487 = n7356 | n7357 ;
  assign n4701 = n30209 & n4686 ;
  assign n4722 = n1556 & n4706 ;
  assign n4729 = n30196 & n4726 ;
  assign n7488 = n4722 | n4729 ;
  assign n7489 = n1445 & n4748 ;
  assign n7490 = n7488 | n7489 ;
  assign n7491 = n4701 | n7490 ;
  assign n30951 = ~n7491 ;
  assign n7492 = x20 & n30951 ;
  assign n7493 = n30374 & n7491 ;
  assign n7494 = n7492 | n7493 ;
  assign n7495 = n7487 | n7494 ;
  assign n7496 = n7487 & n7494 ;
  assign n30952 = ~n7496 ;
  assign n7497 = n7495 & n30952 ;
  assign n30953 = ~n7352 ;
  assign n7353 = n7204 & n30953 ;
  assign n30954 = ~n7204 ;
  assign n7498 = n30954 & n7352 ;
  assign n7499 = n7353 | n7498 ;
  assign n4700 = n3307 & n4686 ;
  assign n4736 = n30105 & n4726 ;
  assign n4752 = n1556 & n4748 ;
  assign n7500 = n4736 | n4752 ;
  assign n7501 = n30196 & n4706 ;
  assign n7502 = n7500 | n7501 ;
  assign n7503 = n4700 | n7502 ;
  assign n30955 = ~n7503 ;
  assign n7504 = x20 & n30955 ;
  assign n7505 = n30374 & n7503 ;
  assign n7506 = n7504 | n7505 ;
  assign n30956 = ~n7506 ;
  assign n7507 = n7499 & n30956 ;
  assign n30957 = ~n7499 ;
  assign n7508 = n30957 & n7506 ;
  assign n7509 = n7507 | n7508 ;
  assign n30958 = ~n7216 ;
  assign n7350 = n30958 & n7349 ;
  assign n30959 = ~n7349 ;
  assign n7510 = n7216 & n30959 ;
  assign n7511 = n7350 | n7510 ;
  assign n4703 = n30233 & n4686 ;
  assign n4742 = n1812 & n4726 ;
  assign n4751 = n30196 & n4748 ;
  assign n7512 = n4742 | n4751 ;
  assign n7513 = n30105 & n4706 ;
  assign n7514 = n7512 | n7513 ;
  assign n7515 = n4703 | n7514 ;
  assign n7516 = x20 | n7515 ;
  assign n7517 = x20 & n7515 ;
  assign n30960 = ~n7517 ;
  assign n7518 = n7516 & n30960 ;
  assign n30961 = ~n7518 ;
  assign n7520 = n7511 & n30961 ;
  assign n7519 = n7511 & n7518 ;
  assign n7521 = n7511 | n7518 ;
  assign n30962 = ~n7519 ;
  assign n7522 = n30962 & n7521 ;
  assign n7347 = n7228 & n7346 ;
  assign n7523 = n7228 | n7346 ;
  assign n30963 = ~n7347 ;
  assign n7524 = n30963 & n7523 ;
  assign n4687 = n4230 & n4686 ;
  assign n4718 = n1812 & n4706 ;
  assign n4756 = n30105 & n4748 ;
  assign n7525 = n4718 | n4756 ;
  assign n7526 = n30108 & n4726 ;
  assign n7527 = n7525 | n7526 ;
  assign n7528 = n4687 | n7527 ;
  assign n7529 = x20 | n7528 ;
  assign n7530 = x20 & n7528 ;
  assign n30964 = ~n7530 ;
  assign n7531 = n7529 & n30964 ;
  assign n7533 = n7524 | n7531 ;
  assign n30965 = ~n7524 ;
  assign n7532 = n30965 & n7531 ;
  assign n30966 = ~n7531 ;
  assign n7534 = n7524 & n30966 ;
  assign n7535 = n7532 | n7534 ;
  assign n30967 = ~n7344 ;
  assign n7536 = n7343 & n30967 ;
  assign n7537 = n7345 | n7536 ;
  assign n4691 = n3592 & n4686 ;
  assign n4744 = n30114 & n4726 ;
  assign n4749 = n1812 & n4748 ;
  assign n7538 = n4744 | n4749 ;
  assign n7539 = n30108 & n4706 ;
  assign n7540 = n7538 | n7539 ;
  assign n7541 = n4691 | n7540 ;
  assign n7542 = x20 | n7541 ;
  assign n7543 = x20 & n7541 ;
  assign n30968 = ~n7543 ;
  assign n7544 = n7542 & n30968 ;
  assign n7546 = n7537 | n7544 ;
  assign n30969 = ~n7537 ;
  assign n7545 = n30969 & n7544 ;
  assign n30970 = ~n7544 ;
  assign n7547 = n7537 & n30970 ;
  assign n7548 = n7545 | n7547 ;
  assign n7337 = n7248 & n7336 ;
  assign n7549 = n7248 | n7336 ;
  assign n30971 = ~n7337 ;
  assign n7550 = n30971 & n7549 ;
  assign n4699 = n30310 & n4686 ;
  assign n4723 = n30114 & n4706 ;
  assign n4745 = n30123 & n4726 ;
  assign n7551 = n4723 | n4745 ;
  assign n7552 = n30108 & n4748 ;
  assign n7553 = n7551 | n7552 ;
  assign n7554 = n4699 | n7553 ;
  assign n7555 = x20 | n7554 ;
  assign n7556 = x20 & n7554 ;
  assign n30972 = ~n7556 ;
  assign n7557 = n7555 & n30972 ;
  assign n7559 = n7550 | n7557 ;
  assign n30973 = ~n7550 ;
  assign n7558 = n30973 & n7557 ;
  assign n30974 = ~n7557 ;
  assign n7560 = n7550 & n30974 ;
  assign n7561 = n7558 | n7560 ;
  assign n7335 = n7260 | n7333 ;
  assign n7562 = n7260 & n7333 ;
  assign n30975 = ~n7562 ;
  assign n7563 = n7335 & n30975 ;
  assign n5256 = n4686 & n5251 ;
  assign n4711 = n30123 & n4706 ;
  assign n4761 = n30114 & n4748 ;
  assign n7564 = n4711 | n4761 ;
  assign n7565 = n2102 & n4726 ;
  assign n7566 = n7564 | n7565 ;
  assign n7567 = n5256 | n7566 ;
  assign n7568 = x20 | n7567 ;
  assign n7569 = x20 & n7567 ;
  assign n30976 = ~n7569 ;
  assign n7570 = n7568 & n30976 ;
  assign n7572 = n7563 | n7570 ;
  assign n7571 = n7563 & n7570 ;
  assign n30977 = ~n7571 ;
  assign n7573 = n30977 & n7572 ;
  assign n7574 = n7329 | n7331 ;
  assign n30978 = ~n7332 ;
  assign n7575 = n30978 & n7574 ;
  assign n5270 = n4686 & n30440 ;
  assign n4708 = n2102 & n4706 ;
  assign n4746 = n2216 & n4726 ;
  assign n7576 = n4708 | n4746 ;
  assign n7577 = n30123 & n4748 ;
  assign n7578 = n7576 | n7577 ;
  assign n7579 = n5270 | n7578 ;
  assign n7580 = x20 | n7579 ;
  assign n7581 = x20 & n7579 ;
  assign n30979 = ~n7581 ;
  assign n7582 = n7580 & n30979 ;
  assign n7584 = n7575 | n7582 ;
  assign n7328 = n7286 | n7326 ;
  assign n7585 = n7286 & n7326 ;
  assign n30980 = ~n7585 ;
  assign n7586 = n7328 & n30980 ;
  assign n4689 = n4352 & n4686 ;
  assign n4707 = n2216 & n4706 ;
  assign n4730 = n2295 & n4726 ;
  assign n7587 = n4707 | n4730 ;
  assign n7588 = n2102 & n4748 ;
  assign n7589 = n7587 | n7588 ;
  assign n7590 = n4689 | n7589 ;
  assign n7591 = x20 | n7590 ;
  assign n7592 = x20 & n7590 ;
  assign n30981 = ~n7592 ;
  assign n7593 = n7591 & n30981 ;
  assign n7595 = n7586 | n7593 ;
  assign n30982 = ~n7586 ;
  assign n7594 = n30982 & n7593 ;
  assign n30983 = ~n7593 ;
  assign n7596 = n7586 & n30983 ;
  assign n7597 = n7594 | n7596 ;
  assign n30984 = ~n7321 ;
  assign n7324 = n30984 & n7323 ;
  assign n30985 = ~n7323 ;
  assign n7598 = n7321 & n30985 ;
  assign n7599 = n7324 | n7598 ;
  assign n5340 = n4686 & n30444 ;
  assign n4713 = n2295 & n4706 ;
  assign n4762 = n2216 & n4748 ;
  assign n7600 = n4713 | n4762 ;
  assign n7601 = n30445 & n4726 ;
  assign n7602 = n7600 | n7601 ;
  assign n7603 = n5340 | n7602 ;
  assign n7604 = x20 | n7603 ;
  assign n7605 = x20 & n7603 ;
  assign n30986 = ~n7605 ;
  assign n7606 = n7604 & n30986 ;
  assign n7608 = n7599 & n7606 ;
  assign n30987 = ~n7599 ;
  assign n7607 = n30987 & n7606 ;
  assign n30988 = ~n7606 ;
  assign n7609 = n7599 & n30988 ;
  assign n7610 = n7607 | n7609 ;
  assign n30989 = ~n6890 ;
  assign n7302 = n30989 & n7301 ;
  assign n30990 = ~n7301 ;
  assign n7611 = n6890 & n30990 ;
  assign n7612 = n7302 | n7611 ;
  assign n30991 = ~n7310 ;
  assign n7613 = n30991 & n7612 ;
  assign n30992 = ~n7612 ;
  assign n7614 = n7310 & n30992 ;
  assign n7615 = n7613 | n7614 ;
  assign n5398 = n4686 & n5392 ;
  assign n4728 = n30157 & n4726 ;
  assign n4763 = n2295 & n4748 ;
  assign n7616 = n4728 | n4763 ;
  assign n7617 = n30445 & n4706 ;
  assign n7618 = n7616 | n7617 ;
  assign n7619 = n5398 | n7618 ;
  assign n7620 = x20 | n7619 ;
  assign n7621 = x20 & n7619 ;
  assign n30993 = ~n7621 ;
  assign n7622 = n7620 & n30993 ;
  assign n7624 = n7615 | n7622 ;
  assign n7625 = n7295 & n7299 ;
  assign n30994 = ~n7625 ;
  assign n7626 = n7300 & n30994 ;
  assign n5449 = n4686 & n30452 ;
  assign n4719 = n30157 & n4706 ;
  assign n4764 = n30445 & n4748 ;
  assign n7627 = n4719 | n4764 ;
  assign n7628 = n30453 & n4726 ;
  assign n7629 = n7627 | n7628 ;
  assign n7630 = n5449 | n7629 ;
  assign n7631 = x20 | n7630 ;
  assign n7632 = x20 & n7630 ;
  assign n30995 = ~n7632 ;
  assign n7633 = n7631 & n30995 ;
  assign n7675 = n7626 | n7633 ;
  assign n30996 = ~n7292 ;
  assign n7293 = n7288 & n30996 ;
  assign n30997 = ~n7288 ;
  assign n7635 = n30997 & n7292 ;
  assign n7636 = n7293 | n7635 ;
  assign n5501 = n4686 & n30458 ;
  assign n4737 = n2639 & n4726 ;
  assign n4759 = n30157 & n4748 ;
  assign n7637 = n4737 | n4759 ;
  assign n7638 = n30453 & n4706 ;
  assign n7639 = n7637 | n7638 ;
  assign n7640 = n5501 | n7639 ;
  assign n7641 = x20 | n7640 ;
  assign n7642 = x20 & n7640 ;
  assign n30998 = ~n7642 ;
  assign n7643 = n7641 & n30998 ;
  assign n7644 = n7636 & n7643 ;
  assign n7645 = n30463 & n4683 ;
  assign n7646 = x20 & n7645 ;
  assign n6577 = n4686 & n6573 ;
  assign n7647 = n30463 & n4706 ;
  assign n7648 = n30155 & n4748 ;
  assign n7649 = n7647 | n7648 ;
  assign n7650 = n6577 | n7649 ;
  assign n7652 = n7646 | n7650 ;
  assign n7653 = x20 & n7652 ;
  assign n5572 = n4686 & n5567 ;
  assign n4721 = n30155 & n4706 ;
  assign n4765 = n2639 & n4748 ;
  assign n7654 = n4721 | n4765 ;
  assign n7655 = n30463 & n4726 ;
  assign n7656 = n7654 | n7655 ;
  assign n7657 = n5572 | n7656 ;
  assign n7658 = n7653 | n7657 ;
  assign n30999 = ~n7658 ;
  assign n7659 = x20 & n30999 ;
  assign n7661 = n7287 | n7659 ;
  assign n5637 = n4686 & n5631 ;
  assign n4720 = n2639 & n4706 ;
  assign n4766 = n30453 & n4748 ;
  assign n7662 = n4720 | n4766 ;
  assign n7663 = n30155 & n4726 ;
  assign n7664 = n7662 | n7663 ;
  assign n7665 = n5637 | n7664 ;
  assign n31000 = ~n7665 ;
  assign n7666 = x20 & n31000 ;
  assign n7667 = n30374 & n7665 ;
  assign n7668 = n7666 | n7667 ;
  assign n7669 = n7661 & n7668 ;
  assign n7670 = n7636 | n7643 ;
  assign n31001 = ~n7644 ;
  assign n7671 = n31001 & n7670 ;
  assign n7673 = n7669 & n7671 ;
  assign n7674 = n7644 | n7673 ;
  assign n7634 = n7626 & n7633 ;
  assign n31002 = ~n7634 ;
  assign n7676 = n31002 & n7675 ;
  assign n31003 = ~n7674 ;
  assign n7677 = n31003 & n7676 ;
  assign n31004 = ~n7677 ;
  assign n7678 = n7675 & n31004 ;
  assign n7623 = n7615 & n7622 ;
  assign n31005 = ~n7623 ;
  assign n7679 = n31005 & n7624 ;
  assign n31006 = ~n7678 ;
  assign n7680 = n31006 & n7679 ;
  assign n31007 = ~n7680 ;
  assign n7681 = n7624 & n31007 ;
  assign n7682 = n7610 & n7681 ;
  assign n7684 = n7608 | n7682 ;
  assign n31008 = ~n7684 ;
  assign n7686 = n7597 & n31008 ;
  assign n31009 = ~n7686 ;
  assign n7687 = n7595 & n31009 ;
  assign n7583 = n7575 & n7582 ;
  assign n31010 = ~n7583 ;
  assign n7688 = n31010 & n7584 ;
  assign n31011 = ~n7687 ;
  assign n7689 = n31011 & n7688 ;
  assign n31012 = ~n7689 ;
  assign n7690 = n7584 & n31012 ;
  assign n31013 = ~n7690 ;
  assign n7692 = n7573 & n31013 ;
  assign n31014 = ~n7692 ;
  assign n7693 = n7572 & n31014 ;
  assign n31015 = ~n7693 ;
  assign n7695 = n7561 & n31015 ;
  assign n31016 = ~n7695 ;
  assign n7696 = n7559 & n31016 ;
  assign n31017 = ~n7696 ;
  assign n7698 = n7548 & n31017 ;
  assign n31018 = ~n7698 ;
  assign n7699 = n7546 & n31018 ;
  assign n31019 = ~n7699 ;
  assign n7700 = n7535 & n31019 ;
  assign n31020 = ~n7700 ;
  assign n7701 = n7533 & n31020 ;
  assign n7703 = n7522 | n7701 ;
  assign n31021 = ~n7520 ;
  assign n7704 = n31021 & n7703 ;
  assign n7706 = n7509 | n7704 ;
  assign n31022 = ~n7507 ;
  assign n7707 = n31022 & n7706 ;
  assign n31023 = ~n7707 ;
  assign n7709 = n7497 & n31023 ;
  assign n31024 = ~n7709 ;
  assign n7710 = n7495 & n31024 ;
  assign n7712 = n7486 | n7710 ;
  assign n31025 = ~n7484 ;
  assign n7713 = n31025 & n7712 ;
  assign n31026 = ~n7713 ;
  assign n7715 = n7474 & n31026 ;
  assign n31027 = ~n7715 ;
  assign n7716 = n7472 & n31027 ;
  assign n7718 = n7461 | n7716 ;
  assign n4692 = n30212 & n4686 ;
  assign n4747 = n30082 & n4726 ;
  assign n4753 = n30074 & n4748 ;
  assign n7719 = n4747 | n4753 ;
  assign n7720 = n1219 & n4706 ;
  assign n7721 = n7719 | n7720 ;
  assign n7722 = n4692 | n7721 ;
  assign n31028 = ~n7722 ;
  assign n7723 = x20 & n31028 ;
  assign n7724 = n30374 & n7722 ;
  assign n7725 = n7723 | n7724 ;
  assign n7717 = n7461 & n7716 ;
  assign n31029 = ~n7717 ;
  assign n7726 = n31029 & n7718 ;
  assign n31030 = ~n7725 ;
  assign n7727 = n31030 & n7726 ;
  assign n31031 = ~n7727 ;
  assign n7728 = n7718 & n31031 ;
  assign n7730 = n7459 | n7728 ;
  assign n3874 = n37300 & n30263 ;
  assign n5158 = n3700 & n5144 ;
  assign n5180 = n3764 & n5166 ;
  assign n7731 = n5158 | n5180 ;
  assign n7732 = n30264 & n5191 ;
  assign n7733 = n7731 | n7732 ;
  assign n7734 = n3874 | n7733 ;
  assign n7735 = x17 | n7734 ;
  assign n7736 = x17 & n7734 ;
  assign n31032 = ~n7736 ;
  assign n7737 = n7735 & n31032 ;
  assign n31033 = ~n7459 ;
  assign n7729 = n31033 & n7728 ;
  assign n31034 = ~n7728 ;
  assign n7738 = n7459 & n31034 ;
  assign n7739 = n7729 | n7738 ;
  assign n31035 = ~n7737 ;
  assign n7741 = n31035 & n7739 ;
  assign n31036 = ~n7741 ;
  assign n7742 = n7730 & n31036 ;
  assign n31037 = ~n7448 ;
  assign n7456 = n31037 & n7455 ;
  assign n31038 = ~n7455 ;
  assign n7743 = n7448 & n31038 ;
  assign n7744 = n7456 | n7743 ;
  assign n31039 = ~n7742 ;
  assign n7745 = n31039 & n7744 ;
  assign n31040 = ~n7745 ;
  assign n7746 = n7457 & n31040 ;
  assign n31041 = ~n7746 ;
  assign n7748 = n7446 & n31041 ;
  assign n6274 = n30512 & n6272 ;
  assign n6203 = n30405 & n6190 ;
  assign n6253 = n4811 & n6244 ;
  assign n7749 = n6203 | n6253 ;
  assign n7750 = n5017 & n6217 ;
  assign n7751 = n7749 | n7750 ;
  assign n7752 = n6274 | n7751 ;
  assign n7753 = x11 | n7752 ;
  assign n7754 = x11 & n7752 ;
  assign n31042 = ~n7754 ;
  assign n7755 = n7753 & n31042 ;
  assign n31043 = ~n7446 ;
  assign n7747 = n31043 & n7746 ;
  assign n7756 = n7747 | n7748 ;
  assign n7757 = n7755 | n7756 ;
  assign n31044 = ~n7748 ;
  assign n7758 = n31044 & n7757 ;
  assign n31045 = ~n7758 ;
  assign n7760 = n7444 & n31045 ;
  assign n31046 = ~n7760 ;
  assign n7761 = n7442 & n31046 ;
  assign n7763 = n7431 | n7761 ;
  assign n31047 = ~n7429 ;
  assign n7764 = n31047 & n7763 ;
  assign n7766 = n7418 | n7764 ;
  assign n7765 = n7418 & n7764 ;
  assign n31048 = ~n7765 ;
  assign n7767 = n31048 & n7766 ;
  assign n31049 = ~n7431 ;
  assign n7762 = n31049 & n7761 ;
  assign n31050 = ~n7761 ;
  assign n7768 = n7431 & n31050 ;
  assign n7769 = n7762 | n7768 ;
  assign n7759 = n7444 & n7758 ;
  assign n7770 = n7444 | n7758 ;
  assign n31051 = ~n7759 ;
  assign n7771 = n31051 & n7770 ;
  assign n7087 = n30540 & n7068 ;
  assign n31052 = ~n7016 ;
  assign n7017 = n67 & n31052 ;
  assign n7032 = n30545 & n7017 ;
  assign n7055 = n30530 & n7041 ;
  assign n7772 = n7032 | n7055 ;
  assign n7773 = n69 & n30535 ;
  assign n7774 = n7772 | n7773 ;
  assign n7775 = n7087 | n7774 ;
  assign n31053 = ~n7775 ;
  assign n7776 = x8 & n31053 ;
  assign n7777 = n30185 & n7775 ;
  assign n7778 = n7776 | n7777 ;
  assign n7779 = n7771 | n7778 ;
  assign n7780 = n7771 & n7778 ;
  assign n31054 = ~n7780 ;
  assign n7781 = n7779 & n31054 ;
  assign n7782 = n7755 & n7756 ;
  assign n31055 = ~n7782 ;
  assign n7783 = n7757 & n31055 ;
  assign n7092 = n30587 & n7068 ;
  assign n7024 = n30535 & n7017 ;
  assign n7044 = n30415 & n7041 ;
  assign n7784 = n7024 | n7044 ;
  assign n7785 = n69 & n30530 ;
  assign n7786 = n7784 | n7785 ;
  assign n7787 = n7092 | n7786 ;
  assign n7788 = x8 | n7787 ;
  assign n7789 = x8 & n7787 ;
  assign n31056 = ~n7789 ;
  assign n7790 = n7788 & n31056 ;
  assign n31057 = ~n7790 ;
  assign n7792 = n7783 & n31057 ;
  assign n7791 = n7783 & n7790 ;
  assign n7793 = n7783 | n7790 ;
  assign n31058 = ~n7791 ;
  assign n7794 = n31058 & n7793 ;
  assign n31059 = ~n7744 ;
  assign n7795 = n7742 & n31059 ;
  assign n7796 = n7745 | n7795 ;
  assign n6277 = n30578 & n6272 ;
  assign n6196 = n4811 & n6190 ;
  assign n6236 = n30405 & n6217 ;
  assign n7797 = n6196 | n6236 ;
  assign n7798 = n4664 & n6244 ;
  assign n7799 = n7797 | n7798 ;
  assign n7800 = n6277 | n7799 ;
  assign n7801 = x11 | n7800 ;
  assign n7802 = x11 & n7800 ;
  assign n31060 = ~n7802 ;
  assign n7803 = n7801 & n31060 ;
  assign n7805 = n7796 | n7803 ;
  assign n7740 = n7737 & n7739 ;
  assign n7806 = n7737 | n7739 ;
  assign n31061 = ~n7740 ;
  assign n7807 = n31061 & n7806 ;
  assign n5952 = n30286 & n5937 ;
  assign n5997 = n4093 & n5994 ;
  assign n6028 = n30282 & n6018 ;
  assign n7808 = n5997 | n6028 ;
  assign n7809 = n4033 & n5970 ;
  assign n7810 = n7808 | n7809 ;
  assign n7811 = n5952 | n7810 ;
  assign n7812 = x14 | n7811 ;
  assign n7813 = x14 & n7811 ;
  assign n31062 = ~n7813 ;
  assign n7814 = n7812 & n31062 ;
  assign n7816 = n7807 | n7814 ;
  assign n7815 = n7807 & n7814 ;
  assign n31063 = ~n7815 ;
  assign n7817 = n31063 & n7816 ;
  assign n31064 = ~n7726 ;
  assign n7818 = n7725 & n31064 ;
  assign n7819 = n7727 | n7818 ;
  assign n3788 = n37300 & n3787 ;
  assign n5149 = n3764 & n5144 ;
  assign n5171 = n1074 & n5166 ;
  assign n7820 = n5149 | n5171 ;
  assign n7821 = n3700 & n5191 ;
  assign n7822 = n7820 | n7821 ;
  assign n7823 = n3788 | n7822 ;
  assign n31065 = ~n7823 ;
  assign n7824 = x17 & n31065 ;
  assign n7825 = n30580 & n7823 ;
  assign n7826 = n7824 | n7825 ;
  assign n7827 = n7819 | n7826 ;
  assign n7828 = n7819 & n7826 ;
  assign n31066 = ~n7828 ;
  assign n7829 = n7827 & n31066 ;
  assign n7714 = n7474 & n7713 ;
  assign n7830 = n7474 | n7713 ;
  assign n31067 = ~n7714 ;
  assign n7831 = n31067 & n7830 ;
  assign n4424 = n37300 & n4420 ;
  assign n5150 = n1074 & n5144 ;
  assign n5196 = n3764 & n5191 ;
  assign n7832 = n5150 | n5196 ;
  assign n7833 = n30074 & n5166 ;
  assign n7834 = n7832 | n7833 ;
  assign n7835 = n4424 | n7834 ;
  assign n31068 = ~n7835 ;
  assign n7836 = x17 & n31068 ;
  assign n7837 = n30580 & n7835 ;
  assign n7838 = n7836 | n7837 ;
  assign n7839 = n7831 | n7838 ;
  assign n7840 = n7831 & n7838 ;
  assign n31069 = ~n7840 ;
  assign n7841 = n7839 & n31069 ;
  assign n31070 = ~n7486 ;
  assign n7711 = n31070 & n7710 ;
  assign n31071 = ~n7710 ;
  assign n7842 = n7486 & n31071 ;
  assign n7843 = n7711 | n7842 ;
  assign n2847 = n37300 & n30173 ;
  assign n5174 = n1219 & n5166 ;
  assign n5197 = n1074 & n5191 ;
  assign n7844 = n5174 | n5197 ;
  assign n7845 = n30074 & n5144 ;
  assign n7846 = n7844 | n7845 ;
  assign n7847 = n2847 | n7846 ;
  assign n7848 = x17 | n7847 ;
  assign n7849 = x17 & n7847 ;
  assign n31072 = ~n7849 ;
  assign n7850 = n7848 & n31072 ;
  assign n31073 = ~n7850 ;
  assign n7852 = n7843 & n31073 ;
  assign n31074 = ~n7843 ;
  assign n7851 = n31074 & n7850 ;
  assign n7853 = n7851 | n7852 ;
  assign n7708 = n7497 & n7707 ;
  assign n7854 = n7497 | n7707 ;
  assign n31075 = ~n7708 ;
  assign n7855 = n31075 & n7854 ;
  assign n3398 = n37300 & n30212 ;
  assign n5163 = n1219 & n5144 ;
  assign n5195 = n30074 & n5191 ;
  assign n7856 = n5163 | n5195 ;
  assign n7857 = n30082 & n5166 ;
  assign n7858 = n7856 | n7857 ;
  assign n7859 = n3398 | n7858 ;
  assign n7860 = x17 | n7859 ;
  assign n7861 = x17 & n7859 ;
  assign n31076 = ~n7861 ;
  assign n7862 = n7860 & n31076 ;
  assign n7864 = n7855 | n7862 ;
  assign n7863 = n7855 & n7862 ;
  assign n31077 = ~n7863 ;
  assign n7865 = n31077 & n7864 ;
  assign n31078 = ~n7704 ;
  assign n7705 = n7509 & n31078 ;
  assign n31079 = ~n7509 ;
  assign n7866 = n31079 & n7704 ;
  assign n7867 = n7705 | n7866 ;
  assign n3629 = n37300 & n30238 ;
  assign n5172 = n1445 & n5166 ;
  assign n5199 = n1219 & n5191 ;
  assign n7868 = n5172 | n5199 ;
  assign n7869 = n30082 & n5144 ;
  assign n7870 = n7868 | n7869 ;
  assign n7871 = n3629 | n7870 ;
  assign n7872 = x17 | n7871 ;
  assign n7873 = x17 & n7871 ;
  assign n31080 = ~n7873 ;
  assign n7874 = n7872 & n31080 ;
  assign n31081 = ~n7867 ;
  assign n7875 = n31081 & n7874 ;
  assign n31082 = ~n7522 ;
  assign n7702 = n31082 & n7701 ;
  assign n31083 = ~n7701 ;
  assign n7876 = n7522 & n31083 ;
  assign n7877 = n7702 | n7876 ;
  assign n3374 = n37300 & n30203 ;
  assign n5151 = n1445 & n5144 ;
  assign n5170 = n1556 & n5166 ;
  assign n7878 = n5151 | n5170 ;
  assign n7879 = n30082 & n5191 ;
  assign n7880 = n7878 | n7879 ;
  assign n7881 = n3374 | n7880 ;
  assign n7882 = x17 | n7881 ;
  assign n7883 = x17 & n7881 ;
  assign n31084 = ~n7883 ;
  assign n7884 = n7882 & n31084 ;
  assign n31085 = ~n7884 ;
  assign n7886 = n7877 & n31085 ;
  assign n31086 = ~n7877 ;
  assign n7885 = n31086 & n7884 ;
  assign n7887 = n7885 | n7886 ;
  assign n31087 = ~n7535 ;
  assign n7888 = n31087 & n7699 ;
  assign n7889 = n7700 | n7888 ;
  assign n3387 = n37300 & n30209 ;
  assign n5154 = n1556 & n5144 ;
  assign n5192 = n1445 & n5191 ;
  assign n7890 = n5154 | n5192 ;
  assign n7891 = n30196 & n5166 ;
  assign n7892 = n7890 | n7891 ;
  assign n7893 = n3387 | n7892 ;
  assign n31088 = ~n7893 ;
  assign n7894 = x17 & n31088 ;
  assign n7895 = n30580 & n7893 ;
  assign n7896 = n7894 | n7895 ;
  assign n7898 = n7889 | n7896 ;
  assign n31089 = ~n7896 ;
  assign n7897 = n7889 & n31089 ;
  assign n31090 = ~n7889 ;
  assign n7899 = n31090 & n7896 ;
  assign n7900 = n7897 | n7899 ;
  assign n3310 = n37300 & n3307 ;
  assign n5182 = n30105 & n5166 ;
  assign n5206 = n1556 & n5191 ;
  assign n7901 = n5182 | n5206 ;
  assign n7902 = n30196 & n5144 ;
  assign n7903 = n7901 | n7902 ;
  assign n7904 = n3310 | n7903 ;
  assign n7905 = x17 | n7904 ;
  assign n7906 = x17 & n7904 ;
  assign n31091 = ~n7906 ;
  assign n7907 = n7905 & n31091 ;
  assign n7697 = n7548 & n7696 ;
  assign n7908 = n7548 | n7696 ;
  assign n31092 = ~n7697 ;
  assign n7909 = n31092 & n7908 ;
  assign n7911 = n7907 | n7909 ;
  assign n31093 = ~n7909 ;
  assign n7910 = n7907 & n31093 ;
  assign n31094 = ~n7907 ;
  assign n7912 = n31094 & n7909 ;
  assign n7913 = n7910 | n7912 ;
  assign n7694 = n7561 & n7693 ;
  assign n7914 = n7561 | n7693 ;
  assign n31095 = ~n7694 ;
  assign n7915 = n31095 & n7914 ;
  assign n3612 = n37300 & n30233 ;
  assign n5187 = n1812 & n5166 ;
  assign n5207 = n30196 & n5191 ;
  assign n7916 = n5187 | n5207 ;
  assign n7917 = n30105 & n5144 ;
  assign n7918 = n7916 | n7917 ;
  assign n7919 = n3612 | n7918 ;
  assign n7920 = x17 | n7919 ;
  assign n7921 = x17 & n7919 ;
  assign n31096 = ~n7921 ;
  assign n7922 = n7920 & n31096 ;
  assign n7924 = n7915 | n7922 ;
  assign n7923 = n7915 & n7922 ;
  assign n31097 = ~n7923 ;
  assign n7925 = n31097 & n7924 ;
  assign n7691 = n7573 & n7690 ;
  assign n7926 = n7573 | n7690 ;
  assign n31098 = ~n7691 ;
  assign n7927 = n31098 & n7926 ;
  assign n4235 = n37300 & n4230 ;
  assign n5147 = n1812 & n5144 ;
  assign n5193 = n30105 & n5191 ;
  assign n7928 = n5147 | n5193 ;
  assign n7929 = n30108 & n5166 ;
  assign n7930 = n7928 | n7929 ;
  assign n7931 = n4235 | n7930 ;
  assign n7932 = x17 | n7931 ;
  assign n7933 = x17 & n7931 ;
  assign n31099 = ~n7933 ;
  assign n7934 = n7932 & n31099 ;
  assign n7936 = n7927 | n7934 ;
  assign n31100 = ~n7927 ;
  assign n7935 = n31100 & n7934 ;
  assign n31101 = ~n7934 ;
  assign n7937 = n7927 & n31101 ;
  assign n7938 = n7935 | n7937 ;
  assign n31102 = ~n7688 ;
  assign n7939 = n7687 & n31102 ;
  assign n7940 = n7689 | n7939 ;
  assign n3595 = n37300 & n3592 ;
  assign n5184 = n30114 & n5166 ;
  assign n5209 = n1812 & n5191 ;
  assign n7941 = n5184 | n5209 ;
  assign n7942 = n30108 & n5144 ;
  assign n7943 = n7941 | n7942 ;
  assign n7944 = n3595 | n7943 ;
  assign n7945 = x17 | n7944 ;
  assign n7946 = x17 & n7944 ;
  assign n31103 = ~n7946 ;
  assign n7947 = n7945 & n31103 ;
  assign n7949 = n7940 | n7947 ;
  assign n31104 = ~n7940 ;
  assign n7948 = n31104 & n7947 ;
  assign n31105 = ~n7947 ;
  assign n7950 = n7940 & n31105 ;
  assign n7951 = n7948 | n7950 ;
  assign n7685 = n7597 | n7684 ;
  assign n7952 = n7597 & n7684 ;
  assign n31106 = ~n7952 ;
  assign n7953 = n7685 & n31106 ;
  assign n4382 = n37300 & n30310 ;
  assign n5145 = n30114 & n5144 ;
  assign n5185 = n30123 & n5166 ;
  assign n7954 = n5145 | n5185 ;
  assign n7955 = n30108 & n5191 ;
  assign n7956 = n7954 | n7955 ;
  assign n7957 = n4382 | n7956 ;
  assign n7958 = x17 | n7957 ;
  assign n7959 = x17 & n7957 ;
  assign n31107 = ~n7959 ;
  assign n7960 = n7958 & n31107 ;
  assign n7962 = n7953 | n7960 ;
  assign n31108 = ~n7953 ;
  assign n7961 = n31108 & n7960 ;
  assign n31109 = ~n7960 ;
  assign n7963 = n7953 & n31109 ;
  assign n7964 = n7961 | n7963 ;
  assign n31110 = ~n7610 ;
  assign n7683 = n31110 & n7681 ;
  assign n31111 = ~n7681 ;
  assign n7965 = n7610 & n31111 ;
  assign n7966 = n7683 | n7965 ;
  assign n5257 = n37300 & n5251 ;
  assign n5160 = n30123 & n5144 ;
  assign n5210 = n30114 & n5191 ;
  assign n7967 = n5160 | n5210 ;
  assign n7968 = n2102 & n5166 ;
  assign n7969 = n7967 | n7968 ;
  assign n7970 = n5257 | n7969 ;
  assign n7971 = x17 | n7970 ;
  assign n7972 = x17 & n7970 ;
  assign n31112 = ~n7972 ;
  assign n7973 = n7971 & n31112 ;
  assign n7975 = n7966 & n7973 ;
  assign n31113 = ~n7966 ;
  assign n7974 = n31113 & n7973 ;
  assign n31114 = ~n7973 ;
  assign n7976 = n7966 & n31114 ;
  assign n7977 = n7974 | n7976 ;
  assign n5275 = n37300 & n30440 ;
  assign n5157 = n2102 & n5144 ;
  assign n5183 = n2216 & n5166 ;
  assign n7978 = n5157 | n5183 ;
  assign n7979 = n30123 & n5191 ;
  assign n7980 = n7978 | n7979 ;
  assign n7981 = n5275 | n7980 ;
  assign n7982 = x17 | n7981 ;
  assign n7983 = x17 & n7981 ;
  assign n31115 = ~n7983 ;
  assign n7984 = n7982 & n31115 ;
  assign n31116 = ~n7676 ;
  assign n7985 = n7674 & n31116 ;
  assign n7986 = n7677 | n7985 ;
  assign n4354 = n37300 & n4352 ;
  assign n5161 = n2216 & n5144 ;
  assign n5186 = n2295 & n5166 ;
  assign n7987 = n5161 | n5186 ;
  assign n7988 = n2102 & n5191 ;
  assign n7989 = n7987 | n7988 ;
  assign n7990 = n4354 | n7989 ;
  assign n7991 = x17 | n7990 ;
  assign n7992 = x17 & n7990 ;
  assign n31117 = ~n7992 ;
  assign n7993 = n7991 & n31117 ;
  assign n7995 = n7986 | n7993 ;
  assign n31118 = ~n7986 ;
  assign n7994 = n31118 & n7993 ;
  assign n31119 = ~n7993 ;
  assign n7996 = n7986 & n31119 ;
  assign n7997 = n7994 | n7996 ;
  assign n31120 = ~n7669 ;
  assign n7672 = n31120 & n7671 ;
  assign n31121 = ~n7671 ;
  assign n7998 = n7669 & n31121 ;
  assign n7999 = n7672 | n7998 ;
  assign n5341 = n37300 & n30444 ;
  assign n5159 = n2295 & n5144 ;
  assign n5188 = n30445 & n5166 ;
  assign n8000 = n5159 | n5188 ;
  assign n8001 = n2216 & n5191 ;
  assign n8002 = n8000 | n8001 ;
  assign n8003 = n5341 | n8002 ;
  assign n31122 = ~n8003 ;
  assign n8004 = x17 & n31122 ;
  assign n8005 = n30580 & n8003 ;
  assign n8006 = n8004 | n8005 ;
  assign n8007 = n7999 | n8006 ;
  assign n8008 = n7999 & n8006 ;
  assign n31123 = ~n8008 ;
  assign n8009 = n8007 & n31123 ;
  assign n5397 = n37300 & n5392 ;
  assign n5167 = n30157 & n5166 ;
  assign n5211 = n2295 & n5191 ;
  assign n8010 = n5167 | n5211 ;
  assign n8011 = n30445 & n5144 ;
  assign n8012 = n8010 | n8011 ;
  assign n8013 = n5397 | n8012 ;
  assign n8014 = x17 | n8013 ;
  assign n8015 = x17 & n8013 ;
  assign n31124 = ~n8015 ;
  assign n8016 = n8014 & n31124 ;
  assign n31125 = ~n7287 ;
  assign n7660 = n31125 & n7659 ;
  assign n31126 = ~n7659 ;
  assign n8017 = n7287 & n31126 ;
  assign n8018 = n7660 | n8017 ;
  assign n31127 = ~n7668 ;
  assign n8019 = n31127 & n8018 ;
  assign n31128 = ~n8018 ;
  assign n8020 = n7668 & n31128 ;
  assign n8021 = n8019 | n8020 ;
  assign n8023 = n8016 | n8021 ;
  assign n8024 = n7653 & n7657 ;
  assign n31129 = ~n8024 ;
  assign n8025 = n7658 & n31129 ;
  assign n5451 = n37300 & n30452 ;
  assign n5155 = n30157 & n5144 ;
  assign n5212 = n30445 & n5191 ;
  assign n8026 = n5155 | n5212 ;
  assign n8027 = n30453 & n5166 ;
  assign n8028 = n8026 | n8027 ;
  assign n8029 = n5451 | n8028 ;
  assign n8030 = x17 | n8029 ;
  assign n8031 = x17 & n8029 ;
  assign n31130 = ~n8031 ;
  assign n8032 = n8030 & n31130 ;
  assign n8034 = n8025 | n8032 ;
  assign n31131 = ~n7650 ;
  assign n7651 = n7646 & n31131 ;
  assign n31132 = ~n7646 ;
  assign n8035 = n31132 & n7650 ;
  assign n8036 = n7651 | n8035 ;
  assign n5502 = n37300 & n30458 ;
  assign n5189 = n2639 & n5166 ;
  assign n5208 = n30157 & n5191 ;
  assign n8037 = n5189 | n5208 ;
  assign n8038 = n30453 & n5144 ;
  assign n8039 = n8037 | n8038 ;
  assign n8040 = n5502 | n8039 ;
  assign n8041 = x17 | n8040 ;
  assign n8042 = x17 & n8040 ;
  assign n31133 = ~n8042 ;
  assign n8043 = n8041 & n31133 ;
  assign n8044 = n8036 & n8043 ;
  assign n8045 = n37297 & n30463 ;
  assign n8046 = x17 & n8045 ;
  assign n6579 = n37300 & n6573 ;
  assign n8047 = n30463 & n5144 ;
  assign n8048 = n30155 & n5191 ;
  assign n8049 = n8047 | n8048 ;
  assign n8050 = n6579 | n8049 ;
  assign n8052 = n8046 | n8050 ;
  assign n8053 = x17 & n8052 ;
  assign n5573 = n37300 & n5567 ;
  assign n5173 = n30463 & n5166 ;
  assign n8054 = n30155 & n5144 ;
  assign n8055 = n2639 & n5191 ;
  assign n8056 = n8054 | n8055 ;
  assign n8057 = n5173 | n8056 ;
  assign n8058 = n5573 | n8057 ;
  assign n8060 = n8053 | n8058 ;
  assign n31134 = ~n8060 ;
  assign n8061 = x17 & n31134 ;
  assign n8063 = n7645 | n8061 ;
  assign n5634 = n37300 & n5631 ;
  assign n5148 = n2639 & n5144 ;
  assign n5194 = n30453 & n5191 ;
  assign n8064 = n5148 | n5194 ;
  assign n8065 = n30155 & n5166 ;
  assign n8066 = n8064 | n8065 ;
  assign n8067 = n5634 | n8066 ;
  assign n31135 = ~n8067 ;
  assign n8068 = x17 & n31135 ;
  assign n8069 = n30580 & n8067 ;
  assign n8070 = n8068 | n8069 ;
  assign n8071 = n8063 & n8070 ;
  assign n8072 = n8036 | n8043 ;
  assign n31136 = ~n8044 ;
  assign n8073 = n31136 & n8072 ;
  assign n8075 = n8071 & n8073 ;
  assign n8076 = n8044 | n8075 ;
  assign n8033 = n8025 & n8032 ;
  assign n31137 = ~n8033 ;
  assign n8077 = n31137 & n8034 ;
  assign n31138 = ~n8076 ;
  assign n8079 = n31138 & n8077 ;
  assign n31139 = ~n8079 ;
  assign n8080 = n8034 & n31139 ;
  assign n8022 = n8016 & n8021 ;
  assign n31140 = ~n8022 ;
  assign n8081 = n31140 & n8023 ;
  assign n31141 = ~n8080 ;
  assign n8082 = n31141 & n8081 ;
  assign n31142 = ~n8082 ;
  assign n8083 = n8023 & n31142 ;
  assign n31143 = ~n8083 ;
  assign n8085 = n8009 & n31143 ;
  assign n31144 = ~n8085 ;
  assign n8086 = n8007 & n31144 ;
  assign n31145 = ~n8086 ;
  assign n8087 = n7997 & n31145 ;
  assign n31146 = ~n8087 ;
  assign n8088 = n7995 & n31146 ;
  assign n8090 = n7984 | n8088 ;
  assign n31147 = ~n7679 ;
  assign n8091 = n7678 & n31147 ;
  assign n8092 = n7680 | n8091 ;
  assign n8089 = n7984 & n8088 ;
  assign n31148 = ~n8089 ;
  assign n8093 = n31148 & n8090 ;
  assign n31149 = ~n8092 ;
  assign n8094 = n31149 & n8093 ;
  assign n31150 = ~n8094 ;
  assign n8095 = n8090 & n31150 ;
  assign n8097 = n7977 & n8095 ;
  assign n8098 = n7975 | n8097 ;
  assign n31151 = ~n8098 ;
  assign n8100 = n7964 & n31151 ;
  assign n31152 = ~n8100 ;
  assign n8101 = n7962 & n31152 ;
  assign n31153 = ~n8101 ;
  assign n8102 = n7951 & n31153 ;
  assign n31154 = ~n8102 ;
  assign n8103 = n7949 & n31154 ;
  assign n31155 = ~n8103 ;
  assign n8105 = n7938 & n31155 ;
  assign n31156 = ~n8105 ;
  assign n8106 = n7936 & n31156 ;
  assign n31157 = ~n8106 ;
  assign n8108 = n7925 & n31157 ;
  assign n31158 = ~n8108 ;
  assign n8109 = n7924 & n31158 ;
  assign n31159 = ~n8109 ;
  assign n8110 = n7913 & n31159 ;
  assign n31160 = ~n8110 ;
  assign n8111 = n7911 & n31160 ;
  assign n31161 = ~n8111 ;
  assign n8113 = n7900 & n31161 ;
  assign n31162 = ~n8113 ;
  assign n8114 = n7898 & n31162 ;
  assign n8116 = n7887 | n8114 ;
  assign n31163 = ~n7886 ;
  assign n8117 = n31163 & n8116 ;
  assign n31164 = ~n7874 ;
  assign n8118 = n7867 & n31164 ;
  assign n8119 = n7875 | n8118 ;
  assign n31165 = ~n8119 ;
  assign n8121 = n8117 & n31165 ;
  assign n8122 = n7875 | n8121 ;
  assign n31166 = ~n8122 ;
  assign n8124 = n7865 & n31166 ;
  assign n31167 = ~n8124 ;
  assign n8125 = n7864 & n31167 ;
  assign n8127 = n7853 | n8125 ;
  assign n31168 = ~n7852 ;
  assign n8128 = n31168 & n8127 ;
  assign n31169 = ~n8128 ;
  assign n8130 = n7841 & n31169 ;
  assign n31170 = ~n8130 ;
  assign n8131 = n7839 & n31170 ;
  assign n31171 = ~n8131 ;
  assign n8133 = n7829 & n31171 ;
  assign n31172 = ~n8133 ;
  assign n8134 = n7827 & n31172 ;
  assign n31173 = ~n8134 ;
  assign n8136 = n7817 & n31173 ;
  assign n31174 = ~n8136 ;
  assign n8137 = n7816 & n31174 ;
  assign n7804 = n7796 & n7803 ;
  assign n31175 = ~n7804 ;
  assign n8138 = n31175 & n7805 ;
  assign n31176 = ~n8137 ;
  assign n8140 = n31176 & n8138 ;
  assign n31177 = ~n8140 ;
  assign n8141 = n7805 & n31177 ;
  assign n8143 = n7794 | n8141 ;
  assign n31178 = ~n7792 ;
  assign n8144 = n31178 & n8143 ;
  assign n31179 = ~n8144 ;
  assign n8146 = n7781 & n31179 ;
  assign n31180 = ~n8146 ;
  assign n8147 = n7779 & n31180 ;
  assign n31181 = ~n8147 ;
  assign n8149 = n7769 & n31181 ;
  assign n8148 = n7769 & n8147 ;
  assign n8150 = n7769 | n8147 ;
  assign n31182 = ~n8148 ;
  assign n8151 = n31182 & n8150 ;
  assign n8145 = n7781 & n8144 ;
  assign n8152 = n7781 | n8144 ;
  assign n31183 = ~n8145 ;
  assign n8153 = n31183 & n8152 ;
  assign n8142 = n7794 & n8141 ;
  assign n31184 = ~n8142 ;
  assign n8154 = n31184 & n8143 ;
  assign n37291 = x4 & x5 ;
  assign n8155 = x4 | x5 ;
  assign n31185 = ~n37291 ;
  assign n8156 = n31185 & n8155 ;
  assign n8157 = n738 & n8156 ;
  assign n8176 = n30597 & n8157 ;
  assign n31186 = ~n741 ;
  assign n8195 = n31186 & n8156 ;
  assign n8224 = n8176 | n8195 ;
  assign n8225 = n30545 & n8224 ;
  assign n8226 = x5 & n8225 ;
  assign n8227 = x5 | n8225 ;
  assign n31187 = ~n8226 ;
  assign n8228 = n31187 & n8227 ;
  assign n31188 = ~n8228 ;
  assign n8230 = n8154 & n31188 ;
  assign n8229 = n8154 & n8228 ;
  assign n8231 = n8154 | n8228 ;
  assign n31189 = ~n8229 ;
  assign n8232 = n31189 & n8231 ;
  assign n8139 = n8137 & n8138 ;
  assign n8233 = n8137 | n8138 ;
  assign n31190 = ~n8139 ;
  assign n8234 = n31190 & n8233 ;
  assign n7083 = n6411 & n7068 ;
  assign n4935 = n69 & n30415 ;
  assign n7051 = n5017 & n7041 ;
  assign n8235 = n4935 | n7051 ;
  assign n8236 = n30530 & n7017 ;
  assign n8237 = n8235 | n8236 ;
  assign n8238 = n7083 | n8237 ;
  assign n8239 = x8 | n8238 ;
  assign n8240 = x8 & n8238 ;
  assign n31191 = ~n8240 ;
  assign n8241 = n8239 & n31191 ;
  assign n8243 = n8234 | n8241 ;
  assign n8135 = n7817 & n8134 ;
  assign n8244 = n7817 | n8134 ;
  assign n31192 = ~n8135 ;
  assign n8245 = n31192 & n8244 ;
  assign n6290 = n30385 & n6272 ;
  assign n6228 = n4811 & n6217 ;
  assign n6255 = n30361 & n6244 ;
  assign n8246 = n6228 | n6255 ;
  assign n8247 = n4664 & n6190 ;
  assign n8248 = n8246 | n8247 ;
  assign n8249 = n6290 | n8248 ;
  assign n8250 = x11 | n8249 ;
  assign n8251 = x11 & n8249 ;
  assign n31193 = ~n8251 ;
  assign n8252 = n8250 & n31193 ;
  assign n8254 = n8245 | n8252 ;
  assign n31194 = ~n8245 ;
  assign n8253 = n31194 & n8252 ;
  assign n31195 = ~n8252 ;
  assign n8255 = n8245 & n31195 ;
  assign n8256 = n8253 | n8255 ;
  assign n8132 = n7829 & n8131 ;
  assign n8257 = n7829 | n8131 ;
  assign n31196 = ~n8132 ;
  assign n8258 = n31196 & n8257 ;
  assign n5938 = n4442 & n5937 ;
  assign n5978 = n4093 & n5970 ;
  assign n6026 = n4033 & n6018 ;
  assign n8259 = n5978 | n6026 ;
  assign n8260 = n30264 & n5994 ;
  assign n8261 = n8259 | n8260 ;
  assign n8262 = n5938 | n8261 ;
  assign n8263 = x14 | n8262 ;
  assign n8264 = x14 & n8262 ;
  assign n31197 = ~n8264 ;
  assign n8265 = n8263 & n31197 ;
  assign n8267 = n8258 | n8265 ;
  assign n8266 = n8258 & n8265 ;
  assign n31198 = ~n8266 ;
  assign n8268 = n31198 & n8267 ;
  assign n8129 = n7841 & n8128 ;
  assign n8269 = n7841 | n8128 ;
  assign n31199 = ~n8129 ;
  assign n8270 = n31199 & n8269 ;
  assign n5951 = n30349 & n5937 ;
  assign n5998 = n3700 & n5994 ;
  assign n6021 = n4093 & n6018 ;
  assign n8271 = n5998 | n6021 ;
  assign n8272 = n30264 & n5970 ;
  assign n8273 = n8271 | n8272 ;
  assign n8274 = n5951 | n8273 ;
  assign n31200 = ~n8274 ;
  assign n8275 = x14 & n31200 ;
  assign n8276 = n30547 & n8274 ;
  assign n8277 = n8275 | n8276 ;
  assign n8278 = n8270 | n8277 ;
  assign n8279 = n8270 & n8277 ;
  assign n31201 = ~n8279 ;
  assign n8280 = n8278 & n31201 ;
  assign n31202 = ~n7853 ;
  assign n8126 = n31202 & n8125 ;
  assign n31203 = ~n8125 ;
  assign n8281 = n7853 & n31203 ;
  assign n8282 = n8126 | n8281 ;
  assign n5946 = n30263 & n5937 ;
  assign n5975 = n3700 & n5970 ;
  assign n6004 = n3764 & n5994 ;
  assign n8283 = n5975 | n6004 ;
  assign n8284 = n30264 & n6018 ;
  assign n8285 = n8283 | n8284 ;
  assign n8286 = n5946 | n8285 ;
  assign n8287 = x14 | n8286 ;
  assign n8288 = x14 & n8286 ;
  assign n31204 = ~n8288 ;
  assign n8289 = n8287 & n31204 ;
  assign n31205 = ~n8289 ;
  assign n8291 = n8282 & n31205 ;
  assign n31206 = ~n8282 ;
  assign n8290 = n31206 & n8289 ;
  assign n8292 = n8290 | n8291 ;
  assign n8123 = n7865 | n8122 ;
  assign n8293 = n7865 & n8122 ;
  assign n31207 = ~n8293 ;
  assign n8294 = n8123 & n31207 ;
  assign n5956 = n3787 & n5937 ;
  assign n5977 = n3764 & n5970 ;
  assign n6003 = n1074 & n5994 ;
  assign n8295 = n5977 | n6003 ;
  assign n8296 = n3700 & n6018 ;
  assign n8297 = n8295 | n8296 ;
  assign n8298 = n5956 | n8297 ;
  assign n31208 = ~n8298 ;
  assign n8299 = x14 & n31208 ;
  assign n8300 = n30547 & n8298 ;
  assign n8301 = n8299 | n8300 ;
  assign n8302 = n8294 | n8301 ;
  assign n8303 = n8294 & n8301 ;
  assign n31209 = ~n8303 ;
  assign n8304 = n8302 & n31209 ;
  assign n8120 = n8117 | n8119 ;
  assign n8305 = n8117 & n8119 ;
  assign n31210 = ~n8305 ;
  assign n8306 = n8120 & n31210 ;
  assign n5959 = n4420 & n5937 ;
  assign n5971 = n1074 & n5970 ;
  assign n6020 = n3764 & n6018 ;
  assign n8307 = n5971 | n6020 ;
  assign n8308 = n30074 & n5994 ;
  assign n8309 = n8307 | n8308 ;
  assign n8310 = n5959 | n8309 ;
  assign n31211 = ~n8310 ;
  assign n8311 = x14 & n31211 ;
  assign n8312 = n30547 & n8310 ;
  assign n8313 = n8311 | n8312 ;
  assign n31212 = ~n8313 ;
  assign n8314 = n8306 & n31212 ;
  assign n31213 = ~n8306 ;
  assign n8315 = n31213 & n8313 ;
  assign n8316 = n8314 | n8315 ;
  assign n8115 = n7887 & n8114 ;
  assign n31214 = ~n8115 ;
  assign n8317 = n31214 & n8116 ;
  assign n5966 = n30173 & n5937 ;
  assign n6012 = n1219 & n5994 ;
  assign n6019 = n1074 & n6018 ;
  assign n8318 = n6012 | n6019 ;
  assign n8319 = n30074 & n5970 ;
  assign n8320 = n8318 | n8319 ;
  assign n8321 = n5966 | n8320 ;
  assign n8322 = x14 | n8321 ;
  assign n8323 = x14 & n8321 ;
  assign n31215 = ~n8323 ;
  assign n8324 = n8322 & n31215 ;
  assign n31216 = ~n8324 ;
  assign n8326 = n8317 & n31216 ;
  assign n8325 = n8317 & n8324 ;
  assign n8327 = n8317 | n8324 ;
  assign n31217 = ~n8325 ;
  assign n8328 = n31217 & n8327 ;
  assign n31218 = ~n7900 ;
  assign n8112 = n31218 & n8111 ;
  assign n8329 = n8112 | n8113 ;
  assign n5954 = n30212 & n5937 ;
  assign n6011 = n30082 & n5994 ;
  assign n6024 = n30074 & n6018 ;
  assign n8330 = n6011 | n6024 ;
  assign n8331 = n1219 & n5970 ;
  assign n8332 = n8330 | n8331 ;
  assign n8333 = n5954 | n8332 ;
  assign n8334 = x14 | n8333 ;
  assign n8335 = x14 & n8333 ;
  assign n31219 = ~n8335 ;
  assign n8336 = n8334 & n31219 ;
  assign n8338 = n8329 | n8336 ;
  assign n8337 = n8329 & n8336 ;
  assign n31220 = ~n8337 ;
  assign n8339 = n31220 & n8338 ;
  assign n5957 = n30238 & n5937 ;
  assign n5972 = n30082 & n5970 ;
  assign n6023 = n1219 & n6018 ;
  assign n8340 = n5972 | n6023 ;
  assign n8341 = n1445 & n5994 ;
  assign n8342 = n8340 | n8341 ;
  assign n8343 = n5957 | n8342 ;
  assign n8344 = x14 | n8343 ;
  assign n8345 = x14 & n8343 ;
  assign n31221 = ~n8345 ;
  assign n8346 = n8344 & n31221 ;
  assign n8107 = n7925 & n8106 ;
  assign n8347 = n7925 | n8106 ;
  assign n31222 = ~n8107 ;
  assign n8348 = n31222 & n8347 ;
  assign n31223 = ~n7938 ;
  assign n8104 = n31223 & n8103 ;
  assign n8349 = n8104 | n8105 ;
  assign n5943 = n30209 & n5937 ;
  assign n5973 = n1556 & n5970 ;
  assign n6034 = n1445 & n6018 ;
  assign n8350 = n5973 | n6034 ;
  assign n8351 = n30196 & n5994 ;
  assign n8352 = n8350 | n8351 ;
  assign n8353 = n5943 | n8352 ;
  assign n31224 = ~n8353 ;
  assign n8354 = x14 & n31224 ;
  assign n8355 = n30547 & n8353 ;
  assign n8356 = n8354 | n8355 ;
  assign n8357 = n8349 | n8356 ;
  assign n8358 = n8349 & n8356 ;
  assign n31225 = ~n8358 ;
  assign n8359 = n8357 & n31225 ;
  assign n31226 = ~n7951 ;
  assign n8360 = n31226 & n8101 ;
  assign n8361 = n8102 | n8360 ;
  assign n5955 = n3307 & n5937 ;
  assign n5985 = n30196 & n5970 ;
  assign n6027 = n1556 & n6018 ;
  assign n8362 = n5985 | n6027 ;
  assign n8363 = n30105 & n5994 ;
  assign n8364 = n8362 | n8363 ;
  assign n8365 = n5955 | n8364 ;
  assign n31227 = ~n8365 ;
  assign n8366 = x14 & n31227 ;
  assign n8367 = n30547 & n8365 ;
  assign n8368 = n8366 | n8367 ;
  assign n8369 = n8361 | n8368 ;
  assign n8370 = n8361 & n8368 ;
  assign n31228 = ~n8370 ;
  assign n8371 = n8369 & n31228 ;
  assign n8099 = n7964 | n8098 ;
  assign n8372 = n7964 & n8098 ;
  assign n31229 = ~n8372 ;
  assign n8373 = n8099 & n31229 ;
  assign n5960 = n4230 & n5937 ;
  assign n5988 = n1812 & n5970 ;
  assign n6035 = n30105 & n6018 ;
  assign n8374 = n5988 | n6035 ;
  assign n8375 = n30108 & n5994 ;
  assign n8376 = n8374 | n8375 ;
  assign n8377 = n5960 | n8376 ;
  assign n8378 = x14 | n8377 ;
  assign n8379 = x14 & n8377 ;
  assign n31230 = ~n8379 ;
  assign n8380 = n8378 & n31230 ;
  assign n31231 = ~n8093 ;
  assign n8381 = n8092 & n31231 ;
  assign n8382 = n8094 | n8381 ;
  assign n5939 = n3592 & n5937 ;
  assign n5996 = n30114 & n5994 ;
  assign n6038 = n1812 & n6018 ;
  assign n8383 = n5996 | n6038 ;
  assign n8384 = n30108 & n5970 ;
  assign n8385 = n8383 | n8384 ;
  assign n8386 = n5939 | n8385 ;
  assign n31232 = ~n8386 ;
  assign n8387 = x14 & n31232 ;
  assign n8388 = n30547 & n8386 ;
  assign n8389 = n8387 | n8388 ;
  assign n8390 = n8382 | n8389 ;
  assign n8391 = n8382 & n8389 ;
  assign n31233 = ~n8391 ;
  assign n8392 = n8390 & n31233 ;
  assign n31234 = ~n7997 ;
  assign n8393 = n31234 & n8086 ;
  assign n8394 = n8087 | n8393 ;
  assign n5965 = n30310 & n5937 ;
  assign n5976 = n30114 & n5970 ;
  assign n5995 = n30123 & n5994 ;
  assign n8395 = n5976 | n5995 ;
  assign n8396 = n30108 & n6018 ;
  assign n8397 = n8395 | n8396 ;
  assign n8398 = n5965 | n8397 ;
  assign n31235 = ~n8398 ;
  assign n8399 = x14 & n31235 ;
  assign n8400 = n30547 & n8398 ;
  assign n8401 = n8399 | n8400 ;
  assign n8402 = n8394 | n8401 ;
  assign n8403 = n8394 & n8401 ;
  assign n31236 = ~n8403 ;
  assign n8404 = n8402 & n31236 ;
  assign n31237 = ~n8009 ;
  assign n8084 = n31237 & n8083 ;
  assign n8405 = n8084 | n8085 ;
  assign n5961 = n5251 & n5937 ;
  assign n5974 = n30123 & n5970 ;
  assign n6039 = n30114 & n6018 ;
  assign n8406 = n5974 | n6039 ;
  assign n8407 = n2102 & n5994 ;
  assign n8408 = n8406 | n8407 ;
  assign n8409 = n5961 | n8408 ;
  assign n31238 = ~n8409 ;
  assign n8410 = x14 & n31238 ;
  assign n8411 = n30547 & n8409 ;
  assign n8412 = n8410 | n8411 ;
  assign n8414 = n8405 | n8412 ;
  assign n31239 = ~n8412 ;
  assign n8413 = n8405 & n31239 ;
  assign n31240 = ~n8405 ;
  assign n8415 = n31240 & n8412 ;
  assign n8416 = n8413 | n8415 ;
  assign n31241 = ~n8081 ;
  assign n8417 = n8080 & n31241 ;
  assign n8418 = n8082 | n8417 ;
  assign n5967 = n30440 & n5937 ;
  assign n5986 = n2102 & n5970 ;
  assign n6014 = n2216 & n5994 ;
  assign n8419 = n5986 | n6014 ;
  assign n8420 = n30123 & n6018 ;
  assign n8421 = n8419 | n8420 ;
  assign n8422 = n5967 | n8421 ;
  assign n8423 = x14 | n8422 ;
  assign n8424 = x14 & n8422 ;
  assign n31242 = ~n8424 ;
  assign n8425 = n8423 & n31242 ;
  assign n8427 = n8418 | n8425 ;
  assign n8426 = n8418 & n8425 ;
  assign n31243 = ~n8426 ;
  assign n8428 = n31243 & n8427 ;
  assign n31244 = ~n8077 ;
  assign n8078 = n8076 & n31244 ;
  assign n8429 = n8078 | n8079 ;
  assign n5958 = n4352 & n5937 ;
  assign n6000 = n2295 & n5994 ;
  assign n6037 = n2102 & n6018 ;
  assign n8430 = n6000 | n6037 ;
  assign n8431 = n2216 & n5970 ;
  assign n8432 = n8430 | n8431 ;
  assign n8433 = n5958 | n8432 ;
  assign n8434 = x14 | n8433 ;
  assign n8435 = x14 & n8433 ;
  assign n31245 = ~n8435 ;
  assign n8436 = n8434 & n31245 ;
  assign n8438 = n8429 | n8436 ;
  assign n31246 = ~n8429 ;
  assign n8437 = n31246 & n8436 ;
  assign n31247 = ~n8436 ;
  assign n8439 = n8429 & n31247 ;
  assign n8440 = n8437 | n8439 ;
  assign n31248 = ~n8071 ;
  assign n8074 = n31248 & n8073 ;
  assign n31249 = ~n8073 ;
  assign n8441 = n8071 & n31249 ;
  assign n8442 = n8074 | n8441 ;
  assign n5968 = n30444 & n5937 ;
  assign n5987 = n2295 & n5970 ;
  assign n6025 = n2216 & n6018 ;
  assign n8443 = n5987 | n6025 ;
  assign n8444 = n30445 & n5994 ;
  assign n8445 = n8443 | n8444 ;
  assign n8446 = n5968 | n8445 ;
  assign n8447 = x14 | n8446 ;
  assign n8448 = x14 & n8446 ;
  assign n31250 = ~n8448 ;
  assign n8449 = n8447 & n31250 ;
  assign n8450 = n8442 & n8449 ;
  assign n8451 = n8442 | n8449 ;
  assign n31251 = ~n8450 ;
  assign n8452 = n31251 & n8451 ;
  assign n31252 = ~n7645 ;
  assign n8062 = n31252 & n8061 ;
  assign n31253 = ~n8061 ;
  assign n8453 = n7645 & n31253 ;
  assign n8454 = n8062 | n8453 ;
  assign n31254 = ~n8070 ;
  assign n8455 = n31254 & n8454 ;
  assign n31255 = ~n8454 ;
  assign n8456 = n8070 & n31255 ;
  assign n8457 = n8455 | n8456 ;
  assign n5962 = n5392 & n5937 ;
  assign n6008 = n30157 & n5994 ;
  assign n6022 = n2295 & n6018 ;
  assign n8458 = n6008 | n6022 ;
  assign n8459 = n30445 & n5970 ;
  assign n8460 = n8458 | n8459 ;
  assign n8461 = n5962 | n8460 ;
  assign n8462 = x14 | n8461 ;
  assign n8463 = x14 & n8461 ;
  assign n31256 = ~n8463 ;
  assign n8464 = n8462 & n31256 ;
  assign n8466 = n8457 | n8464 ;
  assign n5963 = n30452 & n5937 ;
  assign n5989 = n30157 & n5970 ;
  assign n6015 = n30453 & n5994 ;
  assign n8467 = n5989 | n6015 ;
  assign n8468 = n30445 & n6018 ;
  assign n8469 = n8467 | n8468 ;
  assign n8470 = n5963 | n8469 ;
  assign n8471 = x14 | n8470 ;
  assign n8472 = x14 & n8470 ;
  assign n31257 = ~n8472 ;
  assign n8473 = n8471 & n31257 ;
  assign n31258 = ~n8053 ;
  assign n8059 = n31258 & n8058 ;
  assign n31259 = ~n8058 ;
  assign n8474 = n8053 & n31259 ;
  assign n8475 = n8059 | n8474 ;
  assign n8477 = n8473 | n8475 ;
  assign n31260 = ~n8050 ;
  assign n8051 = n8046 & n31260 ;
  assign n31261 = ~n8046 ;
  assign n8478 = n31261 & n8050 ;
  assign n8479 = n8051 | n8478 ;
  assign n5945 = n30458 & n5937 ;
  assign n6010 = n2639 & n5994 ;
  assign n6033 = n30157 & n6018 ;
  assign n8480 = n6010 | n6033 ;
  assign n8481 = n30453 & n5970 ;
  assign n8482 = n8480 | n8481 ;
  assign n8483 = n5945 | n8482 ;
  assign n8484 = x14 | n8483 ;
  assign n8485 = x14 & n8483 ;
  assign n31262 = ~n8485 ;
  assign n8486 = n8484 & n31262 ;
  assign n8487 = n8479 & n8486 ;
  assign n8488 = n30463 & n5934 ;
  assign n8489 = x14 & n8488 ;
  assign n6580 = n5937 & n6573 ;
  assign n8490 = n30463 & n5970 ;
  assign n8491 = n30155 & n6018 ;
  assign n8492 = n8490 | n8491 ;
  assign n8493 = n6580 | n8492 ;
  assign n8495 = n8489 | n8493 ;
  assign n8496 = x14 & n8495 ;
  assign n5950 = n5567 & n5937 ;
  assign n5990 = n30155 & n5970 ;
  assign n6040 = n2639 & n6018 ;
  assign n8497 = n5990 | n6040 ;
  assign n8498 = n30463 & n5994 ;
  assign n8499 = n8497 | n8498 ;
  assign n8500 = n5950 | n8499 ;
  assign n8501 = n8496 | n8500 ;
  assign n31263 = ~n8501 ;
  assign n8502 = x14 & n31263 ;
  assign n8504 = n8045 | n8502 ;
  assign n5942 = n5631 & n5937 ;
  assign n5991 = n2639 & n5970 ;
  assign n6041 = n30453 & n6018 ;
  assign n8505 = n5991 | n6041 ;
  assign n8506 = n30155 & n5994 ;
  assign n8507 = n8505 | n8506 ;
  assign n8508 = n5942 | n8507 ;
  assign n31264 = ~n8508 ;
  assign n8509 = x14 & n31264 ;
  assign n8510 = n30547 & n8508 ;
  assign n8511 = n8509 | n8510 ;
  assign n8512 = n8504 & n8511 ;
  assign n8513 = n8479 | n8486 ;
  assign n31265 = ~n8487 ;
  assign n8514 = n31265 & n8513 ;
  assign n8516 = n8512 & n8514 ;
  assign n8517 = n8487 | n8516 ;
  assign n8476 = n8473 & n8475 ;
  assign n31266 = ~n8476 ;
  assign n8518 = n31266 & n8477 ;
  assign n31267 = ~n8517 ;
  assign n8520 = n31267 & n8518 ;
  assign n31268 = ~n8520 ;
  assign n8521 = n8477 & n31268 ;
  assign n8465 = n8457 & n8464 ;
  assign n31269 = ~n8465 ;
  assign n8522 = n31269 & n8466 ;
  assign n31270 = ~n8521 ;
  assign n8523 = n31270 & n8522 ;
  assign n31271 = ~n8523 ;
  assign n8524 = n8466 & n31271 ;
  assign n8525 = n8452 & n8524 ;
  assign n8526 = n8450 | n8525 ;
  assign n31272 = ~n8526 ;
  assign n8527 = n8440 & n31272 ;
  assign n31273 = ~n8527 ;
  assign n8528 = n8438 & n31273 ;
  assign n31274 = ~n8528 ;
  assign n8530 = n8428 & n31274 ;
  assign n31275 = ~n8530 ;
  assign n8531 = n8427 & n31275 ;
  assign n31276 = ~n8531 ;
  assign n8532 = n8416 & n31276 ;
  assign n31277 = ~n8532 ;
  assign n8533 = n8414 & n31277 ;
  assign n31278 = ~n8533 ;
  assign n8535 = n8404 & n31278 ;
  assign n31279 = ~n8535 ;
  assign n8536 = n8402 & n31279 ;
  assign n31280 = ~n8536 ;
  assign n8537 = n8392 & n31280 ;
  assign n31281 = ~n8537 ;
  assign n8538 = n8390 & n31281 ;
  assign n8540 = n8380 | n8538 ;
  assign n31282 = ~n7977 ;
  assign n8096 = n31282 & n8095 ;
  assign n31283 = ~n8095 ;
  assign n8541 = n7977 & n31283 ;
  assign n8542 = n8096 | n8541 ;
  assign n8539 = n8380 & n8538 ;
  assign n31284 = ~n8539 ;
  assign n8543 = n31284 & n8540 ;
  assign n31285 = ~n8542 ;
  assign n8544 = n31285 & n8543 ;
  assign n31286 = ~n8544 ;
  assign n8545 = n8540 & n31286 ;
  assign n8547 = n8373 | n8545 ;
  assign n5944 = n30233 & n5937 ;
  assign n6016 = n1812 & n5994 ;
  assign n6029 = n30196 & n6018 ;
  assign n8548 = n6016 | n6029 ;
  assign n8549 = n30105 & n5970 ;
  assign n8550 = n8548 | n8549 ;
  assign n8551 = n5944 | n8550 ;
  assign n31287 = ~n8551 ;
  assign n8552 = x14 & n31287 ;
  assign n8553 = n30547 & n8551 ;
  assign n8554 = n8552 | n8553 ;
  assign n8546 = n8373 & n8545 ;
  assign n31288 = ~n8546 ;
  assign n8555 = n31288 & n8547 ;
  assign n31289 = ~n8554 ;
  assign n8556 = n31289 & n8555 ;
  assign n31290 = ~n8556 ;
  assign n8557 = n8547 & n31290 ;
  assign n31291 = ~n8557 ;
  assign n8559 = n8371 & n31291 ;
  assign n31292 = ~n8559 ;
  assign n8560 = n8369 & n31292 ;
  assign n31293 = ~n8560 ;
  assign n8561 = n8359 & n31293 ;
  assign n31294 = ~n8561 ;
  assign n8562 = n8357 & n31294 ;
  assign n8564 = n8348 | n8562 ;
  assign n5941 = n30203 & n5937 ;
  assign n6017 = n1556 & n5994 ;
  assign n6042 = n30082 & n6018 ;
  assign n8565 = n6017 | n6042 ;
  assign n8566 = n1445 & n5970 ;
  assign n8567 = n8565 | n8566 ;
  assign n8568 = n5941 | n8567 ;
  assign n31295 = ~n8568 ;
  assign n8569 = x14 & n31295 ;
  assign n8570 = n30547 & n8568 ;
  assign n8571 = n8569 | n8570 ;
  assign n8563 = n8348 & n8562 ;
  assign n31296 = ~n8563 ;
  assign n8572 = n31296 & n8564 ;
  assign n31297 = ~n8571 ;
  assign n8573 = n31297 & n8572 ;
  assign n31298 = ~n8573 ;
  assign n8574 = n8564 & n31298 ;
  assign n8576 = n8346 | n8574 ;
  assign n31299 = ~n7913 ;
  assign n8577 = n31299 & n8109 ;
  assign n8578 = n8110 | n8577 ;
  assign n8575 = n8346 & n8574 ;
  assign n31300 = ~n8575 ;
  assign n8579 = n31300 & n8576 ;
  assign n31301 = ~n8578 ;
  assign n8580 = n31301 & n8579 ;
  assign n31302 = ~n8580 ;
  assign n8581 = n8576 & n31302 ;
  assign n31303 = ~n8581 ;
  assign n8583 = n8339 & n31303 ;
  assign n31304 = ~n8583 ;
  assign n8584 = n8338 & n31304 ;
  assign n8585 = n8328 | n8584 ;
  assign n31305 = ~n8326 ;
  assign n8586 = n31305 & n8585 ;
  assign n8588 = n8316 | n8586 ;
  assign n31306 = ~n8314 ;
  assign n8589 = n31306 & n8588 ;
  assign n31307 = ~n8589 ;
  assign n8591 = n8304 & n31307 ;
  assign n31308 = ~n8591 ;
  assign n8592 = n8302 & n31308 ;
  assign n8594 = n8292 | n8592 ;
  assign n31309 = ~n8291 ;
  assign n8595 = n31309 & n8594 ;
  assign n31310 = ~n8595 ;
  assign n8597 = n8280 & n31310 ;
  assign n31311 = ~n8597 ;
  assign n8598 = n8278 & n31311 ;
  assign n31312 = ~n8598 ;
  assign n8600 = n8268 & n31312 ;
  assign n31313 = ~n8600 ;
  assign n8601 = n8267 & n31313 ;
  assign n31314 = ~n8601 ;
  assign n8603 = n8256 & n31314 ;
  assign n31315 = ~n8603 ;
  assign n8604 = n8254 & n31315 ;
  assign n8242 = n8234 & n8241 ;
  assign n31316 = ~n8242 ;
  assign n8605 = n31316 & n8243 ;
  assign n31317 = ~n8604 ;
  assign n8606 = n31317 & n8605 ;
  assign n31318 = ~n8606 ;
  assign n8607 = n8243 & n31318 ;
  assign n8609 = n8232 | n8607 ;
  assign n31319 = ~n8230 ;
  assign n8610 = n31319 & n8609 ;
  assign n8612 = n8153 | n8610 ;
  assign n31320 = ~n8153 ;
  assign n8611 = n31320 & n8610 ;
  assign n31321 = ~n8610 ;
  assign n8613 = n8153 & n31321 ;
  assign n8614 = n8611 | n8613 ;
  assign n31322 = ~n8232 ;
  assign n8608 = n31322 & n8607 ;
  assign n31323 = ~n8607 ;
  assign n8615 = n8232 & n31323 ;
  assign n8616 = n8608 | n8615 ;
  assign n31324 = ~n8605 ;
  assign n8617 = n8604 & n31324 ;
  assign n8618 = n8606 | n8617 ;
  assign n31325 = ~n8256 ;
  assign n8602 = n31325 & n8601 ;
  assign n8619 = n8602 | n8603 ;
  assign n8599 = n8268 & n8598 ;
  assign n8620 = n8268 | n8598 ;
  assign n31326 = ~n8599 ;
  assign n8621 = n31326 & n8620 ;
  assign n6273 = n4674 & n6272 ;
  assign n6204 = n30361 & n6190 ;
  assign n6254 = n30282 & n6244 ;
  assign n8622 = n6204 | n6254 ;
  assign n8623 = n4664 & n6217 ;
  assign n8624 = n8622 | n8623 ;
  assign n8625 = n6273 | n8624 ;
  assign n31327 = ~n8625 ;
  assign n8626 = x11 & n31327 ;
  assign n8627 = n30180 & n8625 ;
  assign n8628 = n8626 | n8627 ;
  assign n8630 = n8621 & n8628 ;
  assign n8596 = n8280 & n8595 ;
  assign n8631 = n8280 | n8595 ;
  assign n31328 = ~n8596 ;
  assign n8632 = n31328 & n8631 ;
  assign n6284 = n5723 & n6272 ;
  assign n6199 = n30282 & n6190 ;
  assign n6237 = n30361 & n6217 ;
  assign n8633 = n6199 | n6237 ;
  assign n8634 = n4033 & n6244 ;
  assign n8635 = n8633 | n8634 ;
  assign n8636 = n6284 | n8635 ;
  assign n8637 = x11 | n8636 ;
  assign n8638 = x11 & n8636 ;
  assign n31329 = ~n8638 ;
  assign n8639 = n8637 & n31329 ;
  assign n8641 = n8632 | n8639 ;
  assign n8640 = n8632 & n8639 ;
  assign n31330 = ~n8640 ;
  assign n8642 = n31330 & n8641 ;
  assign n31331 = ~n8292 ;
  assign n8593 = n31331 & n8592 ;
  assign n31332 = ~n8592 ;
  assign n8643 = n8292 & n31332 ;
  assign n8644 = n8593 | n8643 ;
  assign n6287 = n30286 & n6272 ;
  assign n6231 = n30282 & n6217 ;
  assign n6249 = n4093 & n6244 ;
  assign n8645 = n6231 | n6249 ;
  assign n8646 = n4033 & n6190 ;
  assign n8647 = n8645 | n8646 ;
  assign n8648 = n6287 | n8647 ;
  assign n8649 = x11 | n8648 ;
  assign n8650 = x11 & n8648 ;
  assign n31333 = ~n8650 ;
  assign n8651 = n8649 & n31333 ;
  assign n31334 = ~n8651 ;
  assign n8653 = n8644 & n31334 ;
  assign n31335 = ~n8644 ;
  assign n8652 = n31335 & n8651 ;
  assign n8654 = n8652 | n8653 ;
  assign n8590 = n8304 & n8589 ;
  assign n8655 = n8304 | n8589 ;
  assign n31336 = ~n8590 ;
  assign n8656 = n31336 & n8655 ;
  assign n6294 = n4442 & n6272 ;
  assign n6207 = n4093 & n6190 ;
  assign n6245 = n30264 & n6244 ;
  assign n8657 = n6207 | n6245 ;
  assign n8658 = n4033 & n6217 ;
  assign n8659 = n8657 | n8658 ;
  assign n8660 = n6294 | n8659 ;
  assign n8661 = x11 | n8660 ;
  assign n8662 = x11 & n8660 ;
  assign n31337 = ~n8662 ;
  assign n8663 = n8661 & n31337 ;
  assign n8665 = n8656 | n8663 ;
  assign n31338 = ~n8316 ;
  assign n8587 = n31338 & n8586 ;
  assign n31339 = ~n8586 ;
  assign n8666 = n8316 & n31339 ;
  assign n8667 = n8587 | n8666 ;
  assign n6299 = n30349 & n6272 ;
  assign n6242 = n4093 & n6217 ;
  assign n6247 = n3700 & n6244 ;
  assign n8668 = n6242 | n6247 ;
  assign n8669 = n30264 & n6190 ;
  assign n8670 = n8668 | n8669 ;
  assign n8671 = n6299 | n8670 ;
  assign n31340 = ~n8671 ;
  assign n8672 = x11 & n31340 ;
  assign n8673 = n30180 & n8671 ;
  assign n8674 = n8672 | n8673 ;
  assign n31341 = ~n8674 ;
  assign n8676 = n8667 & n31341 ;
  assign n8675 = n8667 | n8674 ;
  assign n8677 = n8667 & n8674 ;
  assign n31342 = ~n8677 ;
  assign n8678 = n8675 & n31342 ;
  assign n6295 = n30263 & n6272 ;
  assign n6197 = n3700 & n6190 ;
  assign n6251 = n3764 & n6244 ;
  assign n8679 = n6197 | n6251 ;
  assign n8680 = n30264 & n6217 ;
  assign n8681 = n8679 | n8680 ;
  assign n8682 = n6295 | n8681 ;
  assign n8683 = x11 | n8682 ;
  assign n8684 = x11 & n8682 ;
  assign n31343 = ~n8684 ;
  assign n8685 = n8683 & n31343 ;
  assign n8582 = n8339 & n8581 ;
  assign n8686 = n8339 | n8581 ;
  assign n31344 = ~n8582 ;
  assign n8687 = n31344 & n8686 ;
  assign n6296 = n3787 & n6272 ;
  assign n6195 = n3764 & n6190 ;
  assign n6263 = n1074 & n6244 ;
  assign n8688 = n6195 | n6263 ;
  assign n8689 = n3700 & n6217 ;
  assign n8690 = n8688 | n8689 ;
  assign n8691 = n6296 | n8690 ;
  assign n31345 = ~n8691 ;
  assign n8692 = x11 & n31345 ;
  assign n8693 = n30180 & n8691 ;
  assign n8694 = n8692 | n8693 ;
  assign n8696 = n8687 | n8694 ;
  assign n31346 = ~n8694 ;
  assign n8695 = n8687 & n31346 ;
  assign n31347 = ~n8687 ;
  assign n8697 = n31347 & n8694 ;
  assign n8698 = n8695 | n8697 ;
  assign n6298 = n4420 & n6272 ;
  assign n6201 = n1074 & n6190 ;
  assign n6221 = n3764 & n6217 ;
  assign n8699 = n6201 | n6221 ;
  assign n8700 = n30074 & n6244 ;
  assign n8701 = n8699 | n8700 ;
  assign n8702 = n6298 | n8701 ;
  assign n31348 = ~n8702 ;
  assign n8703 = x11 & n31348 ;
  assign n8704 = n30180 & n8702 ;
  assign n8705 = n8703 | n8704 ;
  assign n31349 = ~n8572 ;
  assign n8706 = n8571 & n31349 ;
  assign n8707 = n8573 | n8706 ;
  assign n6301 = n30173 & n6272 ;
  assign n6243 = n1074 & n6217 ;
  assign n6250 = n1219 & n6244 ;
  assign n8708 = n6243 | n6250 ;
  assign n8709 = n30074 & n6190 ;
  assign n8710 = n8708 | n8709 ;
  assign n8711 = n6301 | n8710 ;
  assign n8712 = x11 | n8711 ;
  assign n8713 = x11 & n8711 ;
  assign n31350 = ~n8713 ;
  assign n8714 = n8712 & n31350 ;
  assign n8716 = n8707 | n8714 ;
  assign n8715 = n8707 & n8714 ;
  assign n31351 = ~n8715 ;
  assign n8717 = n31351 & n8716 ;
  assign n31352 = ~n8359 ;
  assign n8718 = n31352 & n8560 ;
  assign n8719 = n8561 | n8718 ;
  assign n6289 = n30212 & n6272 ;
  assign n6194 = n1219 & n6190 ;
  assign n6238 = n30074 & n6217 ;
  assign n8720 = n6194 | n6238 ;
  assign n8721 = n30082 & n6244 ;
  assign n8722 = n8720 | n8721 ;
  assign n8723 = n6289 | n8722 ;
  assign n8724 = x11 | n8723 ;
  assign n8725 = x11 & n8723 ;
  assign n31353 = ~n8725 ;
  assign n8726 = n8724 & n31353 ;
  assign n8728 = n8719 | n8726 ;
  assign n31354 = ~n8719 ;
  assign n8727 = n31354 & n8726 ;
  assign n31355 = ~n8726 ;
  assign n8729 = n8719 & n31355 ;
  assign n8730 = n8727 | n8729 ;
  assign n31356 = ~n8371 ;
  assign n8558 = n31356 & n8557 ;
  assign n8731 = n8558 | n8559 ;
  assign n6297 = n30238 & n6272 ;
  assign n6232 = n1219 & n6217 ;
  assign n6258 = n1445 & n6244 ;
  assign n8732 = n6232 | n6258 ;
  assign n8733 = n30082 & n6190 ;
  assign n8734 = n8732 | n8733 ;
  assign n8735 = n6297 | n8734 ;
  assign n8736 = x11 | n8735 ;
  assign n8737 = x11 & n8735 ;
  assign n31357 = ~n8737 ;
  assign n8738 = n8736 & n31357 ;
  assign n8740 = n8731 | n8738 ;
  assign n31358 = ~n8731 ;
  assign n8739 = n31358 & n8738 ;
  assign n31359 = ~n8738 ;
  assign n8741 = n8731 & n31359 ;
  assign n8742 = n8739 | n8741 ;
  assign n31360 = ~n8555 ;
  assign n8743 = n8554 & n31360 ;
  assign n8744 = n8556 | n8743 ;
  assign n6300 = n30203 & n6272 ;
  assign n6241 = n30082 & n6217 ;
  assign n6259 = n1556 & n6244 ;
  assign n8745 = n6241 | n6259 ;
  assign n8746 = n1445 & n6190 ;
  assign n8747 = n8745 | n8746 ;
  assign n8748 = n6300 | n8747 ;
  assign n31361 = ~n8748 ;
  assign n8749 = x11 & n31361 ;
  assign n8750 = n30180 & n8748 ;
  assign n8751 = n8749 | n8750 ;
  assign n8752 = n8744 | n8751 ;
  assign n8753 = n8744 & n8751 ;
  assign n31362 = ~n8753 ;
  assign n8754 = n8752 & n31362 ;
  assign n31363 = ~n8543 ;
  assign n8755 = n8542 & n31363 ;
  assign n8756 = n8544 | n8755 ;
  assign n6304 = n30209 & n6272 ;
  assign n6192 = n1556 & n6190 ;
  assign n6230 = n1445 & n6217 ;
  assign n8757 = n6192 | n6230 ;
  assign n8758 = n30196 & n6244 ;
  assign n8759 = n8757 | n8758 ;
  assign n8760 = n6304 | n8759 ;
  assign n8761 = x11 | n8760 ;
  assign n8762 = x11 & n8760 ;
  assign n31364 = ~n8762 ;
  assign n8763 = n8761 & n31364 ;
  assign n8765 = n8756 | n8763 ;
  assign n31365 = ~n8756 ;
  assign n8764 = n31365 & n8763 ;
  assign n31366 = ~n8763 ;
  assign n8766 = n8756 & n31366 ;
  assign n8767 = n8764 | n8766 ;
  assign n31367 = ~n8392 ;
  assign n8768 = n31367 & n8536 ;
  assign n8769 = n8537 | n8768 ;
  assign n6303 = n3307 & n6272 ;
  assign n6200 = n30196 & n6190 ;
  assign n6225 = n1556 & n6217 ;
  assign n8770 = n6200 | n6225 ;
  assign n8771 = n30105 & n6244 ;
  assign n8772 = n8770 | n8771 ;
  assign n8773 = n6303 | n8772 ;
  assign n31368 = ~n8773 ;
  assign n8774 = x11 & n31368 ;
  assign n8775 = n30180 & n8773 ;
  assign n8776 = n8774 | n8775 ;
  assign n8777 = n8769 | n8776 ;
  assign n8778 = n8769 & n8776 ;
  assign n31369 = ~n8778 ;
  assign n8779 = n8777 & n31369 ;
  assign n31370 = ~n8404 ;
  assign n8534 = n31370 & n8533 ;
  assign n8780 = n8534 | n8535 ;
  assign n6285 = n30233 & n6272 ;
  assign n6223 = n30196 & n6217 ;
  assign n6252 = n1812 & n6244 ;
  assign n8781 = n6223 | n6252 ;
  assign n8782 = n30105 & n6190 ;
  assign n8783 = n8781 | n8782 ;
  assign n8784 = n6285 | n8783 ;
  assign n8785 = x11 | n8784 ;
  assign n8786 = x11 & n8784 ;
  assign n31371 = ~n8786 ;
  assign n8787 = n8785 & n31371 ;
  assign n8789 = n8780 | n8787 ;
  assign n31372 = ~n8780 ;
  assign n8788 = n31372 & n8787 ;
  assign n31373 = ~n8787 ;
  assign n8790 = n8780 & n31373 ;
  assign n8791 = n8788 | n8790 ;
  assign n31374 = ~n8416 ;
  assign n8792 = n31374 & n8531 ;
  assign n8793 = n8532 | n8792 ;
  assign n6282 = n4230 & n6272 ;
  assign n6210 = n1812 & n6190 ;
  assign n6219 = n30105 & n6217 ;
  assign n8794 = n6210 | n6219 ;
  assign n8795 = n30108 & n6244 ;
  assign n8796 = n8794 | n8795 ;
  assign n8797 = n6282 | n8796 ;
  assign n8798 = x11 | n8797 ;
  assign n8799 = x11 & n8797 ;
  assign n31375 = ~n8799 ;
  assign n8800 = n8798 & n31375 ;
  assign n8802 = n8793 | n8800 ;
  assign n31376 = ~n8793 ;
  assign n8801 = n31376 & n8800 ;
  assign n31377 = ~n8800 ;
  assign n8803 = n8793 & n31377 ;
  assign n8804 = n8801 | n8803 ;
  assign n31378 = ~n8428 ;
  assign n8529 = n31378 & n8528 ;
  assign n8805 = n8529 | n8530 ;
  assign n6305 = n3592 & n6272 ;
  assign n6229 = n1812 & n6217 ;
  assign n6260 = n30114 & n6244 ;
  assign n8806 = n6229 | n6260 ;
  assign n8807 = n30108 & n6190 ;
  assign n8808 = n8806 | n8807 ;
  assign n8809 = n6305 | n8808 ;
  assign n31379 = ~n8809 ;
  assign n8810 = x11 & n31379 ;
  assign n8811 = n30180 & n8809 ;
  assign n8812 = n8810 | n8811 ;
  assign n8813 = n8805 | n8812 ;
  assign n8814 = n8805 & n8812 ;
  assign n31380 = ~n8814 ;
  assign n8815 = n8813 & n31380 ;
  assign n31381 = ~n8440 ;
  assign n8816 = n31381 & n8526 ;
  assign n8817 = n8527 | n8816 ;
  assign n6291 = n30310 & n6272 ;
  assign n6208 = n30114 & n6190 ;
  assign n6262 = n30123 & n6244 ;
  assign n8818 = n6208 | n6262 ;
  assign n8819 = n30108 & n6217 ;
  assign n8820 = n8818 | n8819 ;
  assign n8821 = n6291 | n8820 ;
  assign n8822 = x11 | n8821 ;
  assign n8823 = x11 & n8821 ;
  assign n31382 = ~n8823 ;
  assign n8824 = n8822 & n31382 ;
  assign n8826 = n8817 | n8824 ;
  assign n31383 = ~n8817 ;
  assign n8825 = n31383 & n8824 ;
  assign n31384 = ~n8824 ;
  assign n8827 = n8817 & n31384 ;
  assign n8828 = n8825 | n8827 ;
  assign n8829 = n8452 | n8524 ;
  assign n31385 = ~n8525 ;
  assign n8830 = n31385 & n8829 ;
  assign n6306 = n5251 & n6272 ;
  assign n6198 = n30123 & n6190 ;
  assign n6227 = n30114 & n6217 ;
  assign n8831 = n6198 | n6227 ;
  assign n8832 = n2102 & n6244 ;
  assign n8833 = n8831 | n8832 ;
  assign n8834 = n6306 | n8833 ;
  assign n8835 = x11 | n8834 ;
  assign n8836 = x11 & n8834 ;
  assign n31386 = ~n8836 ;
  assign n8837 = n8835 & n31386 ;
  assign n8838 = n8830 & n8837 ;
  assign n31387 = ~n8522 ;
  assign n8839 = n8521 & n31387 ;
  assign n8840 = n8523 | n8839 ;
  assign n6283 = n30440 & n6272 ;
  assign n6202 = n2102 & n6190 ;
  assign n6226 = n30123 & n6217 ;
  assign n8841 = n6202 | n6226 ;
  assign n8842 = n2216 & n6244 ;
  assign n8843 = n8841 | n8842 ;
  assign n8844 = n6283 | n8843 ;
  assign n8845 = x11 | n8844 ;
  assign n8846 = x11 & n8844 ;
  assign n31388 = ~n8846 ;
  assign n8847 = n8845 & n31388 ;
  assign n8849 = n8840 | n8847 ;
  assign n31389 = ~n8840 ;
  assign n8848 = n31389 & n8847 ;
  assign n31390 = ~n8847 ;
  assign n8850 = n8840 & n31390 ;
  assign n8851 = n8848 | n8850 ;
  assign n31391 = ~n8518 ;
  assign n8519 = n8517 & n31391 ;
  assign n8852 = n8519 | n8520 ;
  assign n6276 = n4352 & n6272 ;
  assign n6209 = n2216 & n6190 ;
  assign n6261 = n2295 & n6244 ;
  assign n8853 = n6209 | n6261 ;
  assign n8854 = n2102 & n6217 ;
  assign n8855 = n8853 | n8854 ;
  assign n8856 = n6276 | n8855 ;
  assign n8857 = x11 | n8856 ;
  assign n8858 = x11 & n8856 ;
  assign n31392 = ~n8858 ;
  assign n8859 = n8857 & n31392 ;
  assign n8861 = n8852 | n8859 ;
  assign n31393 = ~n8852 ;
  assign n8860 = n31393 & n8859 ;
  assign n31394 = ~n8859 ;
  assign n8862 = n8852 & n31394 ;
  assign n8863 = n8860 | n8862 ;
  assign n31395 = ~n8512 ;
  assign n8515 = n31395 & n8514 ;
  assign n31396 = ~n8514 ;
  assign n8864 = n8512 & n31396 ;
  assign n8865 = n8515 | n8864 ;
  assign n6275 = n30444 & n6272 ;
  assign n6211 = n2295 & n6190 ;
  assign n6224 = n2216 & n6217 ;
  assign n8866 = n6211 | n6224 ;
  assign n8867 = n30445 & n6244 ;
  assign n8868 = n8866 | n8867 ;
  assign n8869 = n6275 | n8868 ;
  assign n8870 = x11 | n8869 ;
  assign n8871 = x11 & n8869 ;
  assign n31397 = ~n8871 ;
  assign n8872 = n8870 & n31397 ;
  assign n8874 = n8865 | n8872 ;
  assign n31398 = ~n8045 ;
  assign n8503 = n31398 & n8502 ;
  assign n31399 = ~n8502 ;
  assign n8875 = n8045 & n31399 ;
  assign n8876 = n8503 | n8875 ;
  assign n31400 = ~n8511 ;
  assign n8877 = n31400 & n8876 ;
  assign n31401 = ~n8876 ;
  assign n8878 = n8511 & n31401 ;
  assign n8879 = n8877 | n8878 ;
  assign n6281 = n5392 & n6272 ;
  assign n6222 = n2295 & n6217 ;
  assign n6264 = n30157 & n6244 ;
  assign n8880 = n6222 | n6264 ;
  assign n8881 = n30445 & n6190 ;
  assign n8882 = n8880 | n8881 ;
  assign n8883 = n6281 | n8882 ;
  assign n8884 = x11 | n8883 ;
  assign n8885 = x11 & n8883 ;
  assign n31402 = ~n8885 ;
  assign n8886 = n8884 & n31402 ;
  assign n8888 = n8879 | n8886 ;
  assign n8887 = n8879 & n8886 ;
  assign n31403 = ~n8887 ;
  assign n8889 = n31403 & n8888 ;
  assign n8890 = n8496 & n8500 ;
  assign n31404 = ~n8890 ;
  assign n8891 = n8501 & n31404 ;
  assign n6280 = n30452 & n6272 ;
  assign n6191 = n30157 & n6190 ;
  assign n6239 = n30445 & n6217 ;
  assign n8892 = n6191 | n6239 ;
  assign n8893 = n30453 & n6244 ;
  assign n8894 = n8892 | n8893 ;
  assign n8895 = n6280 | n8894 ;
  assign n8896 = x11 | n8895 ;
  assign n8897 = x11 & n8895 ;
  assign n31405 = ~n8897 ;
  assign n8898 = n8896 & n31405 ;
  assign n8900 = n8891 | n8898 ;
  assign n31406 = ~n8493 ;
  assign n8494 = n8489 & n31406 ;
  assign n31407 = ~n8489 ;
  assign n8901 = n31407 & n8493 ;
  assign n8902 = n8494 | n8901 ;
  assign n6286 = n30458 & n6272 ;
  assign n6220 = n30157 & n6217 ;
  assign n6248 = n2639 & n6244 ;
  assign n8903 = n6220 | n6248 ;
  assign n8904 = n30453 & n6190 ;
  assign n8905 = n8903 | n8904 ;
  assign n8906 = n6286 | n8905 ;
  assign n8907 = x11 | n8906 ;
  assign n8908 = x11 & n8906 ;
  assign n31408 = ~n8908 ;
  assign n8909 = n8907 & n31408 ;
  assign n8910 = n8902 & n8909 ;
  assign n8911 = n30463 & n6188 ;
  assign n8912 = x11 & n8911 ;
  assign n6578 = n6272 & n6573 ;
  assign n8913 = n30463 & n6190 ;
  assign n8914 = n30155 & n6217 ;
  assign n8915 = n8913 | n8914 ;
  assign n8916 = n6578 | n8915 ;
  assign n8918 = n8912 | n8916 ;
  assign n8919 = x11 & n8918 ;
  assign n6279 = n5567 & n6272 ;
  assign n6193 = n30155 & n6190 ;
  assign n6235 = n2639 & n6217 ;
  assign n8920 = n6193 | n6235 ;
  assign n8921 = n30463 & n6244 ;
  assign n8922 = n8920 | n8921 ;
  assign n8923 = n6279 | n8922 ;
  assign n8924 = n8919 | n8923 ;
  assign n31409 = ~n8924 ;
  assign n8925 = x11 & n31409 ;
  assign n8927 = n8488 | n8925 ;
  assign n6278 = n5631 & n6272 ;
  assign n6206 = n2639 & n6190 ;
  assign n6218 = n30453 & n6217 ;
  assign n8928 = n6206 | n6218 ;
  assign n8929 = n30155 & n6244 ;
  assign n8930 = n8928 | n8929 ;
  assign n8931 = n6278 | n8930 ;
  assign n31410 = ~n8931 ;
  assign n8932 = x11 & n31410 ;
  assign n8933 = n30180 & n8931 ;
  assign n8934 = n8932 | n8933 ;
  assign n8935 = n8927 & n8934 ;
  assign n8936 = n8902 | n8909 ;
  assign n31411 = ~n8910 ;
  assign n8937 = n31411 & n8936 ;
  assign n8939 = n8935 & n8937 ;
  assign n8940 = n8910 | n8939 ;
  assign n8899 = n8891 & n8898 ;
  assign n31412 = ~n8899 ;
  assign n8941 = n31412 & n8900 ;
  assign n31413 = ~n8940 ;
  assign n8942 = n31413 & n8941 ;
  assign n31414 = ~n8942 ;
  assign n8943 = n8900 & n31414 ;
  assign n31415 = ~n8943 ;
  assign n8945 = n8889 & n31415 ;
  assign n31416 = ~n8945 ;
  assign n8946 = n8888 & n31416 ;
  assign n8873 = n8865 & n8872 ;
  assign n31417 = ~n8873 ;
  assign n8947 = n31417 & n8874 ;
  assign n31418 = ~n8946 ;
  assign n8948 = n31418 & n8947 ;
  assign n31419 = ~n8948 ;
  assign n8949 = n8874 & n31419 ;
  assign n31420 = ~n8949 ;
  assign n8951 = n8863 & n31420 ;
  assign n31421 = ~n8951 ;
  assign n8952 = n8861 & n31421 ;
  assign n31422 = ~n8952 ;
  assign n8955 = n8851 & n31422 ;
  assign n31423 = ~n8955 ;
  assign n8956 = n8849 & n31423 ;
  assign n8957 = n8830 | n8837 ;
  assign n8958 = n8956 & n8957 ;
  assign n8959 = n8838 | n8958 ;
  assign n31424 = ~n8959 ;
  assign n8962 = n8828 & n31424 ;
  assign n31425 = ~n8962 ;
  assign n8963 = n8826 & n31425 ;
  assign n31426 = ~n8963 ;
  assign n8965 = n8815 & n31426 ;
  assign n31427 = ~n8965 ;
  assign n8966 = n8813 & n31427 ;
  assign n31428 = ~n8966 ;
  assign n8967 = n8804 & n31428 ;
  assign n31429 = ~n8967 ;
  assign n8968 = n8802 & n31429 ;
  assign n31430 = ~n8968 ;
  assign n8971 = n8791 & n31430 ;
  assign n31431 = ~n8971 ;
  assign n8972 = n8789 & n31431 ;
  assign n31432 = ~n8972 ;
  assign n8973 = n8779 & n31432 ;
  assign n31433 = ~n8973 ;
  assign n8974 = n8777 & n31433 ;
  assign n31434 = ~n8974 ;
  assign n8977 = n8767 & n31434 ;
  assign n31435 = ~n8977 ;
  assign n8978 = n8765 & n31435 ;
  assign n31436 = ~n8978 ;
  assign n8979 = n8754 & n31436 ;
  assign n31437 = ~n8979 ;
  assign n8980 = n8752 & n31437 ;
  assign n31438 = ~n8980 ;
  assign n8982 = n8742 & n31438 ;
  assign n31439 = ~n8982 ;
  assign n8983 = n8740 & n31439 ;
  assign n31440 = ~n8983 ;
  assign n8984 = n8730 & n31440 ;
  assign n31441 = ~n8984 ;
  assign n8985 = n8728 & n31441 ;
  assign n31442 = ~n8985 ;
  assign n8987 = n8717 & n31442 ;
  assign n31443 = ~n8987 ;
  assign n8988 = n8716 & n31443 ;
  assign n8990 = n8705 & n8988 ;
  assign n31444 = ~n8579 ;
  assign n8991 = n8578 & n31444 ;
  assign n8992 = n8580 | n8991 ;
  assign n8989 = n8705 | n8988 ;
  assign n31445 = ~n8990 ;
  assign n8993 = n8989 & n31445 ;
  assign n8994 = n8992 & n8993 ;
  assign n8995 = n8990 | n8994 ;
  assign n31446 = ~n8995 ;
  assign n8996 = n8698 & n31446 ;
  assign n31447 = ~n8996 ;
  assign n8997 = n8696 & n31447 ;
  assign n8998 = n8685 & n8997 ;
  assign n8999 = n8328 & n8584 ;
  assign n31448 = ~n8999 ;
  assign n9000 = n8585 & n31448 ;
  assign n9001 = n8685 | n8997 ;
  assign n31449 = ~n8998 ;
  assign n9002 = n31449 & n9001 ;
  assign n31450 = ~n9000 ;
  assign n9003 = n31450 & n9002 ;
  assign n9004 = n8998 | n9003 ;
  assign n9006 = n8678 | n9004 ;
  assign n31451 = ~n8676 ;
  assign n9007 = n31451 & n9006 ;
  assign n8664 = n8656 & n8663 ;
  assign n31452 = ~n8664 ;
  assign n9008 = n31452 & n8665 ;
  assign n31453 = ~n9007 ;
  assign n9009 = n31453 & n9008 ;
  assign n31454 = ~n9009 ;
  assign n9010 = n8665 & n31454 ;
  assign n9012 = n8654 | n9010 ;
  assign n31455 = ~n8653 ;
  assign n9013 = n31455 & n9012 ;
  assign n31456 = ~n9013 ;
  assign n9015 = n8642 & n31456 ;
  assign n31457 = ~n9015 ;
  assign n9016 = n8641 & n31457 ;
  assign n8629 = n8621 | n8628 ;
  assign n31458 = ~n8630 ;
  assign n9017 = n8629 & n31458 ;
  assign n9019 = n9016 & n9017 ;
  assign n9020 = n8630 | n9019 ;
  assign n9021 = n8619 | n9020 ;
  assign n7097 = n30410 & n7068 ;
  assign n7027 = n30415 & n7017 ;
  assign n7054 = n30405 & n7041 ;
  assign n9022 = n7027 | n7054 ;
  assign n9023 = n69 & n5017 ;
  assign n9024 = n9022 | n9023 ;
  assign n9025 = n7097 | n9024 ;
  assign n31459 = ~n9025 ;
  assign n9026 = x8 & n31459 ;
  assign n9027 = n30185 & n9025 ;
  assign n9028 = n9026 | n9027 ;
  assign n9029 = n8619 & n9020 ;
  assign n31460 = ~n9029 ;
  assign n9030 = n9021 & n31460 ;
  assign n31461 = ~n9028 ;
  assign n9031 = n31461 & n9030 ;
  assign n31462 = ~n9031 ;
  assign n9032 = n9021 & n31462 ;
  assign n9034 = n8618 | n9032 ;
  assign n8182 = n6445 & n8157 ;
  assign n9035 = n740 & n30545 ;
  assign n9036 = n30535 & n8195 ;
  assign n9037 = n9035 | n9036 ;
  assign n9038 = n8182 | n9037 ;
  assign n31463 = ~n9038 ;
  assign n9039 = x5 & n31463 ;
  assign n9040 = n30053 & n9038 ;
  assign n9041 = n9039 | n9040 ;
  assign n9033 = n8618 & n9032 ;
  assign n31464 = ~n9033 ;
  assign n9042 = n31464 & n9034 ;
  assign n31465 = ~n9041 ;
  assign n9043 = n31465 & n9042 ;
  assign n31466 = ~n9043 ;
  assign n9044 = n9034 & n31466 ;
  assign n31467 = ~n9044 ;
  assign n9046 = n8616 & n31467 ;
  assign n31468 = ~n8616 ;
  assign n9045 = n31468 & n9044 ;
  assign n9047 = n9045 | n9046 ;
  assign n31469 = ~n9042 ;
  assign n9048 = n9041 & n31469 ;
  assign n9049 = n9043 | n9048 ;
  assign n31470 = ~n9030 ;
  assign n9050 = n9028 & n31470 ;
  assign n9051 = n9031 | n9050 ;
  assign n8185 = n30540 & n8157 ;
  assign n8211 = n30530 & n8195 ;
  assign n31471 = ~n8156 ;
  assign n9052 = n738 & n31471 ;
  assign n9065 = n30545 & n9052 ;
  assign n9074 = n8211 | n9065 ;
  assign n9075 = n740 & n30535 ;
  assign n9076 = n9074 | n9075 ;
  assign n9077 = n8185 | n9076 ;
  assign n31472 = ~n9077 ;
  assign n9078 = x5 & n31472 ;
  assign n9079 = n30053 & n9077 ;
  assign n9080 = n9078 | n9079 ;
  assign n9081 = n9051 | n9080 ;
  assign n31473 = ~n9016 ;
  assign n9018 = n31473 & n9017 ;
  assign n31474 = ~n9017 ;
  assign n9082 = n9016 & n31474 ;
  assign n9083 = n9018 | n9082 ;
  assign n7081 = n30512 & n7068 ;
  assign n5110 = n69 & n30405 ;
  assign n7042 = n4811 & n7041 ;
  assign n9084 = n5110 | n7042 ;
  assign n9085 = n5017 & n7017 ;
  assign n9086 = n9084 | n9085 ;
  assign n9087 = n7081 | n9086 ;
  assign n9088 = x8 | n9087 ;
  assign n9089 = x8 & n9087 ;
  assign n31475 = ~n9089 ;
  assign n9090 = n9088 & n31475 ;
  assign n9092 = n9083 | n9090 ;
  assign n31476 = ~n9083 ;
  assign n9091 = n31476 & n9090 ;
  assign n31477 = ~n9090 ;
  assign n9093 = n9083 & n31477 ;
  assign n9094 = n9091 | n9093 ;
  assign n9014 = n8642 & n9013 ;
  assign n9095 = n8642 | n9013 ;
  assign n31478 = ~n9014 ;
  assign n9096 = n31478 & n9095 ;
  assign n7080 = n30578 & n7068 ;
  assign n4827 = n69 & n4811 ;
  assign n7064 = n4664 & n7041 ;
  assign n9097 = n4827 | n7064 ;
  assign n9098 = n30405 & n7017 ;
  assign n9099 = n9097 | n9098 ;
  assign n9100 = n7080 | n9099 ;
  assign n9101 = x8 | n9100 ;
  assign n9102 = x8 & n9100 ;
  assign n31479 = ~n9102 ;
  assign n9103 = n9101 & n31479 ;
  assign n9105 = n9096 | n9103 ;
  assign n9104 = n9096 & n9103 ;
  assign n31480 = ~n9104 ;
  assign n9106 = n31480 & n9105 ;
  assign n31481 = ~n8654 ;
  assign n9011 = n31481 & n9010 ;
  assign n31482 = ~n9010 ;
  assign n9107 = n8654 & n31482 ;
  assign n9108 = n9011 | n9107 ;
  assign n7100 = n30385 & n7068 ;
  assign n7026 = n4811 & n7017 ;
  assign n7049 = n30361 & n7041 ;
  assign n9109 = n7026 | n7049 ;
  assign n9110 = n69 & n4664 ;
  assign n9111 = n9109 | n9110 ;
  assign n9112 = n7100 | n9111 ;
  assign n9113 = x8 | n9112 ;
  assign n9114 = x8 & n9112 ;
  assign n31483 = ~n9114 ;
  assign n9115 = n9113 & n31483 ;
  assign n31484 = ~n9115 ;
  assign n9117 = n9108 & n31484 ;
  assign n31485 = ~n9108 ;
  assign n9116 = n31485 & n9115 ;
  assign n9118 = n9116 | n9117 ;
  assign n31486 = ~n9008 ;
  assign n9119 = n9007 & n31486 ;
  assign n9120 = n9009 | n9119 ;
  assign n7079 = n4674 & n7068 ;
  assign n4574 = n69 & n30361 ;
  assign n7046 = n30282 & n7041 ;
  assign n9121 = n4574 | n7046 ;
  assign n9122 = n4664 & n7017 ;
  assign n9123 = n9121 | n9122 ;
  assign n9124 = n7079 | n9123 ;
  assign n31487 = ~n9124 ;
  assign n9125 = x8 & n31487 ;
  assign n9126 = n30185 & n9124 ;
  assign n9127 = n9125 | n9126 ;
  assign n9128 = n9120 | n9127 ;
  assign n9129 = n9120 & n9127 ;
  assign n31488 = ~n9129 ;
  assign n9130 = n9128 & n31488 ;
  assign n31489 = ~n9004 ;
  assign n9005 = n8678 & n31489 ;
  assign n31490 = ~n8678 ;
  assign n9131 = n31490 & n9004 ;
  assign n9132 = n9005 | n9131 ;
  assign n7072 = n5723 & n7068 ;
  assign n3941 = n69 & n30282 ;
  assign n7031 = n30361 & n7017 ;
  assign n9133 = n3941 | n7031 ;
  assign n9134 = n4033 & n7041 ;
  assign n9135 = n9133 | n9134 ;
  assign n9136 = n7072 | n9135 ;
  assign n9137 = x8 | n9136 ;
  assign n9138 = x8 & n9136 ;
  assign n31491 = ~n9138 ;
  assign n9139 = n9137 & n31491 ;
  assign n31492 = ~n9139 ;
  assign n9141 = n9132 & n31492 ;
  assign n31493 = ~n9132 ;
  assign n9140 = n31493 & n9139 ;
  assign n9142 = n9140 | n9141 ;
  assign n31494 = ~n9002 ;
  assign n9143 = n9000 & n31494 ;
  assign n9144 = n9003 | n9143 ;
  assign n7089 = n30286 & n7068 ;
  assign n7022 = n30282 & n7017 ;
  assign n7047 = n4093 & n7041 ;
  assign n9145 = n7022 | n7047 ;
  assign n9146 = n69 & n4033 ;
  assign n9147 = n9145 | n9146 ;
  assign n9148 = n7089 | n9147 ;
  assign n9149 = x8 | n9148 ;
  assign n9150 = x8 & n9148 ;
  assign n31495 = ~n9150 ;
  assign n9151 = n9149 & n31495 ;
  assign n31496 = ~n9151 ;
  assign n9153 = n9144 & n31496 ;
  assign n31497 = ~n8698 ;
  assign n9154 = n31497 & n8995 ;
  assign n9155 = n8996 | n9154 ;
  assign n7103 = n4442 & n7068 ;
  assign n4102 = n69 & n4093 ;
  assign n7025 = n4033 & n7017 ;
  assign n9156 = n4102 | n7025 ;
  assign n9157 = n30264 & n7041 ;
  assign n9158 = n9156 | n9157 ;
  assign n9159 = n7103 | n9158 ;
  assign n31498 = ~n9159 ;
  assign n9160 = x8 & n31498 ;
  assign n9161 = n30185 & n9159 ;
  assign n9162 = n9160 | n9161 ;
  assign n9163 = n9155 | n9162 ;
  assign n9164 = n9155 & n9162 ;
  assign n31499 = ~n9164 ;
  assign n9165 = n9163 & n31499 ;
  assign n9166 = n8992 | n8993 ;
  assign n31500 = ~n8994 ;
  assign n9167 = n31500 & n9166 ;
  assign n7094 = n30349 & n7068 ;
  assign n7020 = n4093 & n7017 ;
  assign n7058 = n3700 & n7041 ;
  assign n9168 = n7020 | n7058 ;
  assign n9169 = n69 & n30264 ;
  assign n9170 = n9168 | n9169 ;
  assign n9171 = n7094 | n9170 ;
  assign n9172 = x8 | n9171 ;
  assign n9173 = x8 & n9171 ;
  assign n31501 = ~n9173 ;
  assign n9174 = n9172 & n31501 ;
  assign n9176 = n9167 | n9174 ;
  assign n9175 = n9167 & n9174 ;
  assign n31502 = ~n9175 ;
  assign n9177 = n31502 & n9176 ;
  assign n31503 = ~n8717 ;
  assign n8986 = n31503 & n8985 ;
  assign n9178 = n8986 | n8987 ;
  assign n7096 = n30263 & n7068 ;
  assign n3701 = n69 & n3700 ;
  assign n7053 = n3764 & n7041 ;
  assign n9179 = n3701 | n7053 ;
  assign n9180 = n30264 & n7017 ;
  assign n9181 = n9179 | n9180 ;
  assign n9182 = n7096 | n9181 ;
  assign n9183 = x8 | n9182 ;
  assign n9184 = x8 & n9182 ;
  assign n31504 = ~n9184 ;
  assign n9185 = n9183 & n31504 ;
  assign n9187 = n9178 | n9185 ;
  assign n9186 = n9178 & n9185 ;
  assign n31505 = ~n9186 ;
  assign n9188 = n31505 & n9187 ;
  assign n31506 = ~n8730 ;
  assign n9189 = n31506 & n8983 ;
  assign n9190 = n8984 | n9189 ;
  assign n7084 = n3787 & n7068 ;
  assign n3767 = n69 & n3764 ;
  assign n7050 = n1074 & n7041 ;
  assign n9191 = n3767 | n7050 ;
  assign n9192 = n3700 & n7017 ;
  assign n9193 = n9191 | n9192 ;
  assign n9194 = n7084 | n9193 ;
  assign n31507 = ~n9194 ;
  assign n9195 = x8 & n31507 ;
  assign n9196 = n30185 & n9194 ;
  assign n9197 = n9195 | n9196 ;
  assign n9198 = n9190 | n9197 ;
  assign n9199 = n9190 & n9197 ;
  assign n31508 = ~n9199 ;
  assign n9200 = n9198 & n31508 ;
  assign n31509 = ~n8742 ;
  assign n8981 = n31509 & n8980 ;
  assign n9201 = n8981 | n8982 ;
  assign n7101 = n4420 & n7068 ;
  assign n1079 = n69 & n1074 ;
  assign n7019 = n3764 & n7017 ;
  assign n9202 = n1079 | n7019 ;
  assign n9203 = n30074 & n7041 ;
  assign n9204 = n9202 | n9203 ;
  assign n9205 = n7101 | n9204 ;
  assign n31510 = ~n9205 ;
  assign n9206 = x8 & n31510 ;
  assign n9207 = n30185 & n9205 ;
  assign n9208 = n9206 | n9207 ;
  assign n9210 = n9201 | n9208 ;
  assign n31511 = ~n9208 ;
  assign n9209 = n9201 & n31511 ;
  assign n31512 = ~n9201 ;
  assign n9211 = n31512 & n9208 ;
  assign n9212 = n9209 | n9211 ;
  assign n31513 = ~n8754 ;
  assign n9213 = n31513 & n8978 ;
  assign n9214 = n8979 | n9213 ;
  assign n7090 = n30173 & n7068 ;
  assign n7023 = n1074 & n7017 ;
  assign n7052 = n1219 & n7041 ;
  assign n9215 = n7023 | n7052 ;
  assign n9216 = n69 & n30074 ;
  assign n9217 = n9215 | n9216 ;
  assign n9218 = n7090 | n9217 ;
  assign n9219 = x8 | n9218 ;
  assign n9220 = x8 & n9218 ;
  assign n31514 = ~n9220 ;
  assign n9221 = n9219 & n31514 ;
  assign n9223 = n9214 | n9221 ;
  assign n9222 = n9214 & n9221 ;
  assign n31515 = ~n9222 ;
  assign n9224 = n31515 & n9223 ;
  assign n8975 = n8767 & n8974 ;
  assign n9225 = n8767 | n8974 ;
  assign n31516 = ~n8975 ;
  assign n9226 = n31516 & n9225 ;
  assign n7082 = n30212 & n7068 ;
  assign n7029 = n30074 & n7017 ;
  assign n7059 = n30082 & n7041 ;
  assign n9227 = n7029 | n7059 ;
  assign n9228 = n69 & n1219 ;
  assign n9229 = n9227 | n9228 ;
  assign n9230 = n7082 | n9229 ;
  assign n9231 = x8 | n9230 ;
  assign n9232 = x8 & n9230 ;
  assign n31517 = ~n9232 ;
  assign n9233 = n9231 & n31517 ;
  assign n9234 = n9226 | n9233 ;
  assign n31518 = ~n8767 ;
  assign n8976 = n31518 & n8974 ;
  assign n9235 = n8976 | n8977 ;
  assign n31519 = ~n9235 ;
  assign n9236 = n9233 & n31519 ;
  assign n31520 = ~n9233 ;
  assign n9237 = n31520 & n9235 ;
  assign n9238 = n9236 | n9237 ;
  assign n31521 = ~n8779 ;
  assign n9239 = n31521 & n8972 ;
  assign n9240 = n8973 | n9239 ;
  assign n7099 = n30238 & n7068 ;
  assign n1338 = n69 & n30082 ;
  assign n7048 = n1445 & n7041 ;
  assign n9241 = n1338 | n7048 ;
  assign n9242 = n1219 & n7017 ;
  assign n9243 = n9241 | n9242 ;
  assign n9244 = n7099 | n9243 ;
  assign n9245 = x8 | n9244 ;
  assign n9246 = x8 & n9244 ;
  assign n31522 = ~n9246 ;
  assign n9247 = n9245 & n31522 ;
  assign n9248 = n9240 | n9247 ;
  assign n9251 = n8779 & n8972 ;
  assign n9252 = n8779 | n8972 ;
  assign n31523 = ~n9251 ;
  assign n9253 = n31523 & n9252 ;
  assign n9254 = n9247 & n9253 ;
  assign n9255 = n9247 | n9253 ;
  assign n31524 = ~n9254 ;
  assign n9256 = n31524 & n9255 ;
  assign n8969 = n8791 & n8968 ;
  assign n9257 = n8791 | n8968 ;
  assign n31525 = ~n8969 ;
  assign n9258 = n31525 & n9257 ;
  assign n7095 = n30203 & n7068 ;
  assign n7018 = n30082 & n7017 ;
  assign n7061 = n1556 & n7041 ;
  assign n9259 = n7018 | n7061 ;
  assign n9260 = n69 & n1445 ;
  assign n9261 = n9259 | n9260 ;
  assign n9262 = n7095 | n9261 ;
  assign n31526 = ~n9262 ;
  assign n9263 = x8 & n31526 ;
  assign n9264 = n30185 & n9262 ;
  assign n9265 = n9263 | n9264 ;
  assign n9267 = n9258 | n9265 ;
  assign n31527 = ~n9265 ;
  assign n9266 = n9258 & n31527 ;
  assign n31528 = ~n9258 ;
  assign n9268 = n31528 & n9265 ;
  assign n9269 = n9266 | n9268 ;
  assign n31529 = ~n8804 ;
  assign n9249 = n31529 & n8966 ;
  assign n9270 = n8967 | n9249 ;
  assign n7093 = n30209 & n7068 ;
  assign n1557 = n69 & n1556 ;
  assign n7035 = n1445 & n7017 ;
  assign n9271 = n1557 | n7035 ;
  assign n9272 = n30196 & n7041 ;
  assign n9273 = n9271 | n9272 ;
  assign n9274 = n7093 | n9273 ;
  assign n31530 = ~n9274 ;
  assign n9275 = x8 & n31530 ;
  assign n9276 = n30185 & n9274 ;
  assign n9277 = n9275 | n9276 ;
  assign n9278 = n9270 | n9277 ;
  assign n9279 = n9270 & n9277 ;
  assign n31531 = ~n9279 ;
  assign n9280 = n9278 & n31531 ;
  assign n8964 = n8815 | n8963 ;
  assign n9281 = n8815 & n8963 ;
  assign n31532 = ~n9281 ;
  assign n9282 = n8964 & n31532 ;
  assign n7102 = n3307 & n7068 ;
  assign n7036 = n1556 & n7017 ;
  assign n7043 = n30105 & n7041 ;
  assign n9283 = n7036 | n7043 ;
  assign n9284 = n69 & n30196 ;
  assign n9285 = n9283 | n9284 ;
  assign n9286 = n7102 | n9285 ;
  assign n9287 = x8 | n9286 ;
  assign n9288 = x8 & n9286 ;
  assign n31533 = ~n9288 ;
  assign n9289 = n9287 & n31533 ;
  assign n9291 = n9282 | n9289 ;
  assign n31534 = ~n8815 ;
  assign n9292 = n31534 & n8963 ;
  assign n9293 = n8965 | n9292 ;
  assign n31535 = ~n9293 ;
  assign n9294 = n9289 & n31535 ;
  assign n31536 = ~n9289 ;
  assign n9295 = n31536 & n9293 ;
  assign n9296 = n9294 | n9295 ;
  assign n31537 = ~n8828 ;
  assign n8960 = n31537 & n8959 ;
  assign n9297 = n8960 | n8962 ;
  assign n7091 = n30233 & n7068 ;
  assign n7033 = n30196 & n7017 ;
  assign n7060 = n1812 & n7041 ;
  assign n9298 = n7033 | n7060 ;
  assign n9299 = n69 & n30105 ;
  assign n9300 = n9298 | n9299 ;
  assign n9301 = n7091 | n9300 ;
  assign n9302 = x8 | n9301 ;
  assign n9303 = x8 & n9301 ;
  assign n31538 = ~n9303 ;
  assign n9304 = n9302 & n31538 ;
  assign n9306 = n9297 | n9304 ;
  assign n8961 = n8828 & n8959 ;
  assign n9307 = n8828 | n8959 ;
  assign n31539 = ~n8961 ;
  assign n9308 = n31539 & n9307 ;
  assign n9309 = n9304 & n9308 ;
  assign n9310 = n9304 | n9308 ;
  assign n31540 = ~n9309 ;
  assign n9311 = n31540 & n9310 ;
  assign n31541 = ~n8838 ;
  assign n9312 = n31541 & n8957 ;
  assign n31542 = ~n8956 ;
  assign n9313 = n31542 & n9312 ;
  assign n31543 = ~n9312 ;
  assign n9314 = n8956 & n31543 ;
  assign n9315 = n9313 | n9314 ;
  assign n7085 = n4230 & n7068 ;
  assign n1816 = n69 & n1812 ;
  assign n7037 = n30105 & n7017 ;
  assign n9316 = n1816 | n7037 ;
  assign n9317 = n30108 & n7041 ;
  assign n9318 = n9316 | n9317 ;
  assign n9319 = n7085 | n9318 ;
  assign n9320 = x8 | n9319 ;
  assign n9321 = x8 & n9319 ;
  assign n31544 = ~n9321 ;
  assign n9322 = n9320 & n31544 ;
  assign n9324 = n9315 | n9322 ;
  assign n31545 = ~n9315 ;
  assign n9325 = n31545 & n9322 ;
  assign n31546 = ~n9322 ;
  assign n9326 = n9315 & n31546 ;
  assign n9327 = n9325 | n9326 ;
  assign n31547 = ~n8851 ;
  assign n8953 = n31547 & n8952 ;
  assign n9328 = n8953 | n8955 ;
  assign n7098 = n3592 & n7068 ;
  assign n7034 = n1812 & n7017 ;
  assign n7062 = n30114 & n7041 ;
  assign n9329 = n7034 | n7062 ;
  assign n9330 = n69 & n30108 ;
  assign n9331 = n9329 | n9330 ;
  assign n9332 = n7098 | n9331 ;
  assign n9333 = x8 | n9332 ;
  assign n9334 = x8 & n9332 ;
  assign n31548 = ~n9334 ;
  assign n9335 = n9333 & n31548 ;
  assign n9337 = n9328 | n9335 ;
  assign n8954 = n8851 & n8952 ;
  assign n9338 = n8851 | n8952 ;
  assign n31549 = ~n8954 ;
  assign n9339 = n31549 & n9338 ;
  assign n9340 = n9335 & n9339 ;
  assign n9341 = n9335 | n9339 ;
  assign n31550 = ~n9340 ;
  assign n9342 = n31550 & n9341 ;
  assign n7104 = n30310 & n7068 ;
  assign n1961 = n69 & n30114 ;
  assign n7045 = n30123 & n7041 ;
  assign n9343 = n1961 | n7045 ;
  assign n9344 = n30108 & n7017 ;
  assign n9345 = n9343 | n9344 ;
  assign n9346 = n7104 | n9345 ;
  assign n9347 = x8 | n9346 ;
  assign n9348 = x8 & n9346 ;
  assign n31551 = ~n9348 ;
  assign n9349 = n9347 & n31551 ;
  assign n31552 = ~n8947 ;
  assign n9350 = n8946 & n31552 ;
  assign n9351 = n8948 | n9350 ;
  assign n7105 = n5251 & n7068 ;
  assign n2062 = n69 & n30123 ;
  assign n7038 = n30114 & n7017 ;
  assign n9352 = n2062 | n7038 ;
  assign n9353 = n2102 & n7041 ;
  assign n9354 = n9352 | n9353 ;
  assign n9355 = n7105 | n9354 ;
  assign n31553 = ~n9355 ;
  assign n9356 = x8 & n31553 ;
  assign n9357 = n30185 & n9355 ;
  assign n9358 = n9356 | n9357 ;
  assign n9359 = n9351 | n9358 ;
  assign n9360 = n9351 & n9358 ;
  assign n31554 = ~n9360 ;
  assign n9361 = n9359 & n31554 ;
  assign n31555 = ~n8889 ;
  assign n8944 = n31555 & n8943 ;
  assign n9362 = n8944 | n8945 ;
  assign n7078 = n30440 & n7068 ;
  assign n2104 = n69 & n2102 ;
  assign n7063 = n2216 & n7041 ;
  assign n9363 = n2104 | n7063 ;
  assign n9364 = n30123 & n7017 ;
  assign n9365 = n9363 | n9364 ;
  assign n9366 = n7078 | n9365 ;
  assign n9367 = x8 | n9366 ;
  assign n9368 = x8 & n9366 ;
  assign n31556 = ~n9368 ;
  assign n9369 = n9367 & n31556 ;
  assign n9371 = n9362 | n9369 ;
  assign n31557 = ~n9362 ;
  assign n9370 = n31557 & n9369 ;
  assign n31558 = ~n9369 ;
  assign n9372 = n9362 & n31558 ;
  assign n9373 = n9370 | n9372 ;
  assign n31559 = ~n8941 ;
  assign n9374 = n8940 & n31559 ;
  assign n9375 = n8942 | n9374 ;
  assign n7076 = n4352 & n7068 ;
  assign n7028 = n2102 & n7017 ;
  assign n7056 = n2295 & n7041 ;
  assign n9376 = n7028 | n7056 ;
  assign n9377 = n69 & n2216 ;
  assign n9378 = n9376 | n9377 ;
  assign n9379 = n7076 | n9378 ;
  assign n9380 = x8 | n9379 ;
  assign n9381 = x8 & n9379 ;
  assign n31560 = ~n9381 ;
  assign n9382 = n9380 & n31560 ;
  assign n9384 = n9375 | n9382 ;
  assign n31561 = ~n9375 ;
  assign n9383 = n31561 & n9382 ;
  assign n31562 = ~n9382 ;
  assign n9385 = n9375 & n31562 ;
  assign n9386 = n9383 | n9385 ;
  assign n31563 = ~n8935 ;
  assign n8938 = n31563 & n8937 ;
  assign n31564 = ~n8937 ;
  assign n9387 = n8935 & n31564 ;
  assign n9388 = n8938 | n9387 ;
  assign n7075 = n30444 & n7068 ;
  assign n2297 = n69 & n2295 ;
  assign n7057 = n30445 & n7041 ;
  assign n9389 = n2297 | n7057 ;
  assign n9390 = n2216 & n7017 ;
  assign n9391 = n9389 | n9390 ;
  assign n9392 = n7075 | n9391 ;
  assign n9393 = x8 | n9392 ;
  assign n9394 = x8 & n9392 ;
  assign n31565 = ~n9394 ;
  assign n9395 = n9393 & n31565 ;
  assign n9397 = n9388 | n9395 ;
  assign n31566 = ~n8488 ;
  assign n8926 = n31566 & n8925 ;
  assign n31567 = ~n8925 ;
  assign n9398 = n8488 & n31567 ;
  assign n9399 = n8926 | n9398 ;
  assign n31568 = ~n8934 ;
  assign n9400 = n31568 & n9399 ;
  assign n31569 = ~n9399 ;
  assign n9401 = n8934 & n31569 ;
  assign n9402 = n9400 | n9401 ;
  assign n7074 = n5392 & n7068 ;
  assign n7039 = n2295 & n7017 ;
  assign n7066 = n30157 & n7041 ;
  assign n9403 = n7039 | n7066 ;
  assign n9404 = n69 & n30445 ;
  assign n9405 = n9403 | n9404 ;
  assign n9406 = n7074 | n9405 ;
  assign n9407 = x8 | n9406 ;
  assign n9408 = x8 & n9406 ;
  assign n31570 = ~n9408 ;
  assign n9409 = n9407 & n31570 ;
  assign n9411 = n9402 | n9409 ;
  assign n31571 = ~n9402 ;
  assign n9410 = n31571 & n9409 ;
  assign n31572 = ~n9409 ;
  assign n9412 = n9402 & n31572 ;
  assign n9413 = n9410 | n9412 ;
  assign n9414 = n8919 & n8923 ;
  assign n31573 = ~n9414 ;
  assign n9415 = n8924 & n31573 ;
  assign n7073 = n30452 & n7068 ;
  assign n2780 = n69 & n30157 ;
  assign n7065 = n30453 & n7041 ;
  assign n9416 = n2780 | n7065 ;
  assign n9417 = n30445 & n7017 ;
  assign n9418 = n9416 | n9417 ;
  assign n9419 = n7073 | n9418 ;
  assign n9420 = x8 | n9419 ;
  assign n9421 = x8 & n9419 ;
  assign n31574 = ~n9421 ;
  assign n9422 = n9420 & n31574 ;
  assign n9424 = n9415 | n9422 ;
  assign n31575 = ~n8916 ;
  assign n8917 = n8912 & n31575 ;
  assign n31576 = ~n8912 ;
  assign n9425 = n31576 & n8916 ;
  assign n9426 = n8917 | n9425 ;
  assign n7071 = n30458 & n7068 ;
  assign n2796 = n69 & n30453 ;
  assign n7040 = n30157 & n7017 ;
  assign n9427 = n2796 | n7040 ;
  assign n9428 = n2639 & n7041 ;
  assign n9429 = n9427 | n9428 ;
  assign n9430 = n7071 | n9429 ;
  assign n31577 = ~n9430 ;
  assign n9431 = x8 & n31577 ;
  assign n9432 = n30185 & n9430 ;
  assign n9433 = n9431 | n9432 ;
  assign n9434 = n9426 | n9433 ;
  assign n9435 = n67 & n30463 ;
  assign n9436 = x8 & n9435 ;
  assign n7070 = n6573 & n7068 ;
  assign n9437 = n69 & n30463 ;
  assign n9438 = n30155 & n7017 ;
  assign n9439 = n9437 | n9438 ;
  assign n9440 = n7070 | n9439 ;
  assign n9442 = n9436 | n9440 ;
  assign n9443 = x8 & n9442 ;
  assign n7077 = n5567 & n7068 ;
  assign n2790 = n69 & n30155 ;
  assign n7030 = n2639 & n7017 ;
  assign n9444 = n2790 | n7030 ;
  assign n9445 = n30463 & n7041 ;
  assign n9446 = n9444 | n9445 ;
  assign n9447 = n7077 | n9446 ;
  assign n9448 = n9443 | n9447 ;
  assign n31578 = ~n9448 ;
  assign n9449 = x8 & n31578 ;
  assign n9451 = n8911 | n9449 ;
  assign n7069 = n5631 & n7068 ;
  assign n7021 = n30453 & n7017 ;
  assign n7067 = n30155 & n7041 ;
  assign n9452 = n7021 | n7067 ;
  assign n9453 = n69 & n2639 ;
  assign n9454 = n9452 | n9453 ;
  assign n9455 = n7069 | n9454 ;
  assign n31579 = ~n9455 ;
  assign n9456 = x8 & n31579 ;
  assign n9457 = n30185 & n9455 ;
  assign n9458 = n9456 | n9457 ;
  assign n9459 = n9451 & n9458 ;
  assign n9460 = n9426 & n9433 ;
  assign n31580 = ~n9460 ;
  assign n9461 = n9434 & n31580 ;
  assign n31581 = ~n9459 ;
  assign n9463 = n31581 & n9461 ;
  assign n31582 = ~n9463 ;
  assign n9464 = n9434 & n31582 ;
  assign n9423 = n9415 & n9422 ;
  assign n31583 = ~n9423 ;
  assign n9465 = n31583 & n9424 ;
  assign n31584 = ~n9464 ;
  assign n9466 = n31584 & n9465 ;
  assign n31585 = ~n9466 ;
  assign n9467 = n9424 & n31585 ;
  assign n31586 = ~n9467 ;
  assign n9469 = n9413 & n31586 ;
  assign n31587 = ~n9469 ;
  assign n9470 = n9411 & n31587 ;
  assign n9396 = n9388 & n9395 ;
  assign n31588 = ~n9396 ;
  assign n9471 = n31588 & n9397 ;
  assign n31589 = ~n9470 ;
  assign n9472 = n31589 & n9471 ;
  assign n31590 = ~n9472 ;
  assign n9473 = n9397 & n31590 ;
  assign n31591 = ~n9473 ;
  assign n9475 = n9386 & n31591 ;
  assign n31592 = ~n9475 ;
  assign n9476 = n9384 & n31592 ;
  assign n31593 = ~n9476 ;
  assign n9477 = n9373 & n31593 ;
  assign n31594 = ~n9477 ;
  assign n9478 = n9371 & n31594 ;
  assign n31595 = ~n9478 ;
  assign n9480 = n9361 & n31595 ;
  assign n31596 = ~n9480 ;
  assign n9481 = n9359 & n31596 ;
  assign n9483 = n9349 & n9481 ;
  assign n8950 = n8863 & n8949 ;
  assign n9484 = n8863 | n8949 ;
  assign n31597 = ~n8950 ;
  assign n9485 = n31597 & n9484 ;
  assign n9482 = n9349 | n9481 ;
  assign n31598 = ~n9483 ;
  assign n9486 = n9482 & n31598 ;
  assign n9487 = n9485 & n9486 ;
  assign n9489 = n9483 | n9487 ;
  assign n31599 = ~n9489 ;
  assign n9490 = n9342 & n31599 ;
  assign n31600 = ~n9490 ;
  assign n9491 = n9337 & n31600 ;
  assign n31601 = ~n9491 ;
  assign n9493 = n9327 & n31601 ;
  assign n31602 = ~n9493 ;
  assign n9494 = n9324 & n31602 ;
  assign n31603 = ~n9494 ;
  assign n9495 = n9311 & n31603 ;
  assign n31604 = ~n9495 ;
  assign n9496 = n9306 & n31604 ;
  assign n31605 = ~n9496 ;
  assign n9497 = n9296 & n31605 ;
  assign n31606 = ~n9497 ;
  assign n9498 = n9291 & n31606 ;
  assign n31607 = ~n9498 ;
  assign n9499 = n9280 & n31607 ;
  assign n31608 = ~n9499 ;
  assign n9500 = n9278 & n31608 ;
  assign n31609 = ~n9500 ;
  assign n9502 = n9269 & n31609 ;
  assign n31610 = ~n9502 ;
  assign n9503 = n9267 & n31610 ;
  assign n31611 = ~n9503 ;
  assign n9504 = n9256 & n31611 ;
  assign n31612 = ~n9504 ;
  assign n9505 = n9248 & n31612 ;
  assign n31613 = ~n9505 ;
  assign n9507 = n9238 & n31613 ;
  assign n31614 = ~n9507 ;
  assign n9508 = n9234 & n31614 ;
  assign n31615 = ~n9508 ;
  assign n9509 = n9224 & n31615 ;
  assign n31616 = ~n9509 ;
  assign n9510 = n9223 & n31616 ;
  assign n31617 = ~n9510 ;
  assign n9512 = n9212 & n31617 ;
  assign n31618 = ~n9512 ;
  assign n9513 = n9210 & n31618 ;
  assign n31619 = ~n9513 ;
  assign n9514 = n9200 & n31619 ;
  assign n31620 = ~n9514 ;
  assign n9515 = n9198 & n31620 ;
  assign n31621 = ~n9515 ;
  assign n9517 = n9188 & n31621 ;
  assign n31622 = ~n9517 ;
  assign n9518 = n9187 & n31622 ;
  assign n31623 = ~n9518 ;
  assign n9519 = n9177 & n31623 ;
  assign n31624 = ~n9519 ;
  assign n9520 = n9176 & n31624 ;
  assign n31625 = ~n9520 ;
  assign n9522 = n9165 & n31625 ;
  assign n31626 = ~n9522 ;
  assign n9523 = n9163 & n31626 ;
  assign n31627 = ~n9144 ;
  assign n9152 = n31627 & n9151 ;
  assign n9524 = n9152 | n9153 ;
  assign n9525 = n9523 | n9524 ;
  assign n31628 = ~n9153 ;
  assign n9526 = n31628 & n9525 ;
  assign n9528 = n9142 | n9526 ;
  assign n31629 = ~n9141 ;
  assign n9529 = n31629 & n9528 ;
  assign n31630 = ~n9529 ;
  assign n9531 = n9130 & n31630 ;
  assign n31631 = ~n9531 ;
  assign n9532 = n9128 & n31631 ;
  assign n9534 = n9118 | n9532 ;
  assign n31632 = ~n9117 ;
  assign n9535 = n31632 & n9534 ;
  assign n31633 = ~n9535 ;
  assign n9537 = n9106 & n31633 ;
  assign n31634 = ~n9537 ;
  assign n9538 = n9105 & n31634 ;
  assign n31635 = ~n9538 ;
  assign n9540 = n9094 & n31635 ;
  assign n31636 = ~n9540 ;
  assign n9541 = n9092 & n31636 ;
  assign n9542 = n9051 & n9080 ;
  assign n31637 = ~n9542 ;
  assign n9543 = n9081 & n31637 ;
  assign n31638 = ~n9541 ;
  assign n9544 = n31638 & n9543 ;
  assign n31639 = ~n9544 ;
  assign n9545 = n9081 & n31639 ;
  assign n9547 = n9049 | n9545 ;
  assign n31640 = ~n9049 ;
  assign n9546 = n31640 & n9545 ;
  assign n31641 = ~n9545 ;
  assign n9548 = n9049 & n31641 ;
  assign n9549 = n9546 | n9548 ;
  assign n31642 = ~n9543 ;
  assign n9550 = n9541 & n31642 ;
  assign n9551 = n9544 | n9550 ;
  assign n31643 = ~n733 ;
  assign n9552 = x2 & n31643 ;
  assign n31644 = ~x1 ;
  assign n9559 = n31644 & x2 ;
  assign n37292 = x1 & x2 ;
  assign n9560 = x1 | x2 ;
  assign n31645 = ~n37292 ;
  assign n9561 = n31645 & n9560 ;
  assign n9562 = x0 & n9561 ;
  assign n9581 = n9559 | n9562 ;
  assign n9582 = n30597 & n9581 ;
  assign n9583 = n9552 | n9582 ;
  assign n9584 = n30545 & n9583 ;
  assign n9585 = x2 & n9584 ;
  assign n9586 = x2 | n9584 ;
  assign n31646 = ~n9585 ;
  assign n9587 = n31646 & n9586 ;
  assign n8169 = n30587 & n8157 ;
  assign n5872 = n740 & n30530 ;
  assign n8221 = n30415 & n8195 ;
  assign n9588 = n5872 | n8221 ;
  assign n9589 = n30535 & n9052 ;
  assign n9590 = n9588 | n9589 ;
  assign n9591 = n8169 | n9590 ;
  assign n9592 = x5 | n9591 ;
  assign n9593 = x5 & n9591 ;
  assign n31647 = ~n9593 ;
  assign n9594 = n9592 & n31647 ;
  assign n9595 = n9587 & n9594 ;
  assign n9539 = n9094 & n9538 ;
  assign n9596 = n9094 | n9538 ;
  assign n31648 = ~n9539 ;
  assign n9597 = n31648 & n9596 ;
  assign n9598 = n9587 | n9594 ;
  assign n31649 = ~n9595 ;
  assign n9599 = n31649 & n9598 ;
  assign n9601 = n9597 & n9599 ;
  assign n9602 = n9595 | n9601 ;
  assign n9604 = n9551 | n9602 ;
  assign n31650 = ~n9602 ;
  assign n9603 = n9551 & n31650 ;
  assign n31651 = ~n9551 ;
  assign n9605 = n31651 & n9602 ;
  assign n9606 = n9603 | n9605 ;
  assign n31652 = ~n9597 ;
  assign n9600 = n31652 & n9599 ;
  assign n31653 = ~n9599 ;
  assign n9607 = n9597 & n31653 ;
  assign n9608 = n9600 | n9607 ;
  assign n31654 = ~n9106 ;
  assign n9536 = n31654 & n9535 ;
  assign n9609 = n9536 | n9537 ;
  assign n8190 = n6411 & n8157 ;
  assign n4932 = n740 & n30415 ;
  assign n8223 = n5017 & n8195 ;
  assign n9610 = n4932 | n8223 ;
  assign n9611 = n30530 & n9052 ;
  assign n9612 = n9610 | n9611 ;
  assign n9613 = n8190 | n9612 ;
  assign n31655 = ~n9613 ;
  assign n9614 = x5 & n31655 ;
  assign n9615 = n30053 & n9613 ;
  assign n9616 = n9614 | n9615 ;
  assign n9617 = n9609 | n9616 ;
  assign n9618 = n9609 & n9616 ;
  assign n31656 = ~n9618 ;
  assign n9619 = n9617 & n31656 ;
  assign n31657 = ~n9118 ;
  assign n9533 = n31657 & n9532 ;
  assign n31658 = ~n9532 ;
  assign n9620 = n9118 & n31658 ;
  assign n9621 = n9533 | n9620 ;
  assign n8159 = n30410 & n8157 ;
  assign n8206 = n30405 & n8195 ;
  assign n9063 = n30415 & n9052 ;
  assign n9622 = n8206 | n9063 ;
  assign n9623 = n740 & n5017 ;
  assign n9624 = n9622 | n9623 ;
  assign n9625 = n8159 | n9624 ;
  assign n9626 = x5 | n9625 ;
  assign n9627 = x5 & n9625 ;
  assign n31659 = ~n9627 ;
  assign n9628 = n9626 & n31659 ;
  assign n31660 = ~n9628 ;
  assign n9630 = n9621 & n31660 ;
  assign n31661 = ~n9621 ;
  assign n9629 = n31661 & n9628 ;
  assign n9631 = n9629 | n9630 ;
  assign n9530 = n9130 & n9529 ;
  assign n9632 = n9130 | n9529 ;
  assign n31662 = ~n9530 ;
  assign n9633 = n31662 & n9632 ;
  assign n8173 = n30512 & n8157 ;
  assign n5107 = n740 & n30405 ;
  assign n8202 = n4811 & n8195 ;
  assign n9634 = n5107 | n8202 ;
  assign n9635 = n5017 & n9052 ;
  assign n9636 = n9634 | n9635 ;
  assign n9637 = n8173 | n9636 ;
  assign n31663 = ~n9637 ;
  assign n9638 = x5 & n31663 ;
  assign n9639 = n30053 & n9637 ;
  assign n9640 = n9638 | n9639 ;
  assign n9641 = n9633 | n9640 ;
  assign n9642 = n9633 & n9640 ;
  assign n31664 = ~n9642 ;
  assign n9643 = n9641 & n31664 ;
  assign n31665 = ~n9142 ;
  assign n9527 = n31665 & n9526 ;
  assign n31666 = ~n9526 ;
  assign n9644 = n9142 & n31666 ;
  assign n9645 = n9527 | n9644 ;
  assign n8178 = n30578 & n8157 ;
  assign n4821 = n740 & n4811 ;
  assign n8196 = n4664 & n8195 ;
  assign n9646 = n4821 | n8196 ;
  assign n9647 = n30405 & n9052 ;
  assign n9648 = n9646 | n9647 ;
  assign n9649 = n8178 | n9648 ;
  assign n31667 = ~n9649 ;
  assign n9650 = x5 & n31667 ;
  assign n9651 = n30053 & n9649 ;
  assign n9652 = n9650 | n9651 ;
  assign n31668 = ~n9652 ;
  assign n9653 = n9645 & n31668 ;
  assign n31669 = ~n9645 ;
  assign n9654 = n31669 & n9652 ;
  assign n9655 = n9653 | n9654 ;
  assign n9656 = n9523 & n9524 ;
  assign n31670 = ~n9656 ;
  assign n9657 = n9525 & n31670 ;
  assign n9521 = n9165 & n9520 ;
  assign n9658 = n9165 | n9520 ;
  assign n31671 = ~n9521 ;
  assign n9659 = n31671 & n9658 ;
  assign n8168 = n4674 & n8157 ;
  assign n4577 = n740 & n30361 ;
  assign n8205 = n30282 & n8195 ;
  assign n9660 = n4577 | n8205 ;
  assign n9661 = n4664 & n9052 ;
  assign n9662 = n9660 | n9661 ;
  assign n9663 = n8168 | n9662 ;
  assign n31672 = ~n9663 ;
  assign n9664 = x5 & n31672 ;
  assign n9665 = n30053 & n9663 ;
  assign n9666 = n9664 | n9665 ;
  assign n9667 = n9659 | n9666 ;
  assign n8174 = n5723 & n8157 ;
  assign n3942 = n740 & n30282 ;
  assign n9066 = n30361 & n9052 ;
  assign n9668 = n3942 | n9066 ;
  assign n9669 = n4033 & n8195 ;
  assign n9670 = n9668 | n9669 ;
  assign n9671 = n8174 | n9670 ;
  assign n9672 = x5 | n9671 ;
  assign n9673 = x5 & n9671 ;
  assign n31673 = ~n9673 ;
  assign n9674 = n9672 & n31673 ;
  assign n9516 = n9188 & n9515 ;
  assign n9675 = n9188 | n9515 ;
  assign n31674 = ~n9516 ;
  assign n9676 = n31674 & n9675 ;
  assign n8167 = n30286 & n8157 ;
  assign n8208 = n4093 & n8195 ;
  assign n9062 = n30282 & n9052 ;
  assign n9677 = n8208 | n9062 ;
  assign n9678 = n740 & n4033 ;
  assign n9679 = n9677 | n9678 ;
  assign n9680 = n8167 | n9679 ;
  assign n9681 = x5 | n9680 ;
  assign n9682 = x5 & n9680 ;
  assign n31675 = ~n9682 ;
  assign n9683 = n9681 & n31675 ;
  assign n9685 = n9676 | n9683 ;
  assign n31676 = ~n9676 ;
  assign n9684 = n31676 & n9683 ;
  assign n31677 = ~n9683 ;
  assign n9686 = n9676 & n31677 ;
  assign n9687 = n9684 | n9686 ;
  assign n31678 = ~n9200 ;
  assign n9688 = n31678 & n9513 ;
  assign n9689 = n9514 | n9688 ;
  assign n8162 = n4442 & n8157 ;
  assign n4097 = n740 & n4093 ;
  assign n8198 = n30264 & n8195 ;
  assign n9690 = n4097 | n8198 ;
  assign n9691 = n4033 & n9052 ;
  assign n9692 = n9690 | n9691 ;
  assign n9693 = n8162 | n9692 ;
  assign n9694 = x5 | n9693 ;
  assign n9695 = x5 & n9693 ;
  assign n31679 = ~n9695 ;
  assign n9696 = n9694 & n31679 ;
  assign n9697 = n9689 & n9696 ;
  assign n31680 = ~n9212 ;
  assign n9511 = n31680 & n9510 ;
  assign n9698 = n9511 | n9512 ;
  assign n8186 = n30349 & n8157 ;
  assign n8220 = n3700 & n8195 ;
  assign n9061 = n4093 & n9052 ;
  assign n9699 = n8220 | n9061 ;
  assign n9700 = n740 & n30264 ;
  assign n9701 = n9699 | n9700 ;
  assign n9702 = n8186 | n9701 ;
  assign n31681 = ~n9702 ;
  assign n9703 = x5 & n31681 ;
  assign n9704 = n30053 & n9702 ;
  assign n9705 = n9703 | n9704 ;
  assign n9707 = n9698 & n9705 ;
  assign n9706 = n9698 | n9705 ;
  assign n31682 = ~n9224 ;
  assign n9708 = n31682 & n9508 ;
  assign n9709 = n9509 | n9708 ;
  assign n8179 = n30263 & n8157 ;
  assign n3704 = n740 & n3700 ;
  assign n8203 = n3764 & n8195 ;
  assign n9710 = n3704 | n8203 ;
  assign n9711 = n30264 & n9052 ;
  assign n9712 = n9710 | n9711 ;
  assign n9713 = n8179 | n9712 ;
  assign n9714 = x5 | n9713 ;
  assign n9715 = x5 & n9713 ;
  assign n31683 = ~n9715 ;
  assign n9716 = n9714 & n31683 ;
  assign n9718 = n9709 | n9716 ;
  assign n31684 = ~n9709 ;
  assign n9717 = n31684 & n9716 ;
  assign n31685 = ~n9716 ;
  assign n9719 = n9709 & n31685 ;
  assign n9720 = n9717 | n9719 ;
  assign n31686 = ~n9238 ;
  assign n9506 = n31686 & n9505 ;
  assign n9721 = n9506 | n9507 ;
  assign n8180 = n3787 & n8157 ;
  assign n8199 = n1074 & n8195 ;
  assign n9064 = n3700 & n9052 ;
  assign n9722 = n8199 | n9064 ;
  assign n9723 = n740 & n3764 ;
  assign n9724 = n9722 | n9723 ;
  assign n9725 = n8180 | n9724 ;
  assign n31687 = ~n9725 ;
  assign n9726 = x5 & n31687 ;
  assign n9727 = n30053 & n9725 ;
  assign n9728 = n9726 | n9727 ;
  assign n9730 = n9721 | n9728 ;
  assign n31688 = ~n9728 ;
  assign n9729 = n9721 & n31688 ;
  assign n31689 = ~n9721 ;
  assign n9731 = n31689 & n9728 ;
  assign n9732 = n9729 | n9731 ;
  assign n31690 = ~n8791 ;
  assign n8970 = n31690 & n8968 ;
  assign n9733 = n8970 | n8971 ;
  assign n9734 = n9265 | n9733 ;
  assign n9735 = n9265 & n9733 ;
  assign n31691 = ~n9735 ;
  assign n9736 = n9734 & n31691 ;
  assign n9250 = n8804 & n8966 ;
  assign n9737 = n8804 | n8966 ;
  assign n31692 = ~n9250 ;
  assign n9738 = n31692 & n9737 ;
  assign n9740 = n9277 | n9738 ;
  assign n31693 = ~n9277 ;
  assign n9739 = n31693 & n9738 ;
  assign n31694 = ~n9738 ;
  assign n9741 = n9277 & n31694 ;
  assign n9742 = n9739 | n9741 ;
  assign n9743 = n9289 | n9293 ;
  assign n9290 = n9282 & n9289 ;
  assign n31695 = ~n9290 ;
  assign n9744 = n31695 & n9291 ;
  assign n31696 = ~n9297 ;
  assign n9305 = n31696 & n9304 ;
  assign n31697 = ~n9304 ;
  assign n9746 = n9297 & n31697 ;
  assign n9747 = n9305 | n9746 ;
  assign n9323 = n9315 & n9322 ;
  assign n31698 = ~n9328 ;
  assign n9336 = n31698 & n9335 ;
  assign n31699 = ~n9335 ;
  assign n9748 = n9328 & n31699 ;
  assign n9749 = n9336 | n9748 ;
  assign n9750 = n9482 & n9485 ;
  assign n9751 = n9483 | n9750 ;
  assign n31700 = ~n9751 ;
  assign n9752 = n9749 & n31700 ;
  assign n31701 = ~n9752 ;
  assign n9753 = n9341 & n31701 ;
  assign n9754 = n9323 | n9753 ;
  assign n9755 = n9324 & n9754 ;
  assign n31702 = ~n9755 ;
  assign n9757 = n9747 & n31702 ;
  assign n31703 = ~n9757 ;
  assign n9758 = n9310 & n31703 ;
  assign n31704 = ~n9758 ;
  assign n9759 = n9744 & n31704 ;
  assign n31705 = ~n9759 ;
  assign n9760 = n9743 & n31705 ;
  assign n31706 = ~n9760 ;
  assign n9762 = n9742 & n31706 ;
  assign n31707 = ~n9762 ;
  assign n9763 = n9740 & n31707 ;
  assign n31708 = ~n9763 ;
  assign n9764 = n9736 & n31708 ;
  assign n31709 = ~n9764 ;
  assign n9765 = n9734 & n31709 ;
  assign n9766 = n9256 & n9765 ;
  assign n9767 = n9256 | n9765 ;
  assign n31710 = ~n9766 ;
  assign n9768 = n31710 & n9767 ;
  assign n8177 = n4420 & n8157 ;
  assign n1076 = n740 & n1074 ;
  assign n9059 = n3764 & n9052 ;
  assign n9769 = n1076 | n9059 ;
  assign n9770 = n30074 & n8195 ;
  assign n9771 = n9769 | n9770 ;
  assign n9772 = n8177 | n9771 ;
  assign n31711 = ~n9772 ;
  assign n9773 = x5 & n31711 ;
  assign n9774 = n30053 & n9772 ;
  assign n9775 = n9773 | n9774 ;
  assign n9777 = n9768 | n9775 ;
  assign n31712 = ~n9775 ;
  assign n9776 = n9768 & n31712 ;
  assign n31713 = ~n9768 ;
  assign n9778 = n31713 & n9775 ;
  assign n9779 = n9776 | n9778 ;
  assign n31714 = ~n9269 ;
  assign n9501 = n31714 & n9500 ;
  assign n9780 = n9501 | n9502 ;
  assign n8166 = n30173 & n8157 ;
  assign n8212 = n1219 & n8195 ;
  assign n9057 = n1074 & n9052 ;
  assign n9781 = n8212 | n9057 ;
  assign n9782 = n740 & n30074 ;
  assign n9783 = n9781 | n9782 ;
  assign n9784 = n8166 | n9783 ;
  assign n9785 = x5 | n9784 ;
  assign n9786 = x5 & n9784 ;
  assign n31715 = ~n9786 ;
  assign n9787 = n9785 & n31715 ;
  assign n9788 = n9780 & n9787 ;
  assign n9761 = n9280 & n9760 ;
  assign n9789 = n9280 | n9760 ;
  assign n31716 = ~n9761 ;
  assign n9790 = n31716 & n9789 ;
  assign n8187 = n30212 & n8157 ;
  assign n1223 = n740 & n1219 ;
  assign n8207 = n30082 & n8195 ;
  assign n9791 = n1223 | n8207 ;
  assign n9792 = n30074 & n9052 ;
  assign n9793 = n9791 | n9792 ;
  assign n9794 = n8187 | n9793 ;
  assign n31717 = ~n9794 ;
  assign n9795 = x5 & n31717 ;
  assign n9796 = n30053 & n9794 ;
  assign n9797 = n9795 | n9796 ;
  assign n9799 = n9790 | n9797 ;
  assign n31718 = ~n9797 ;
  assign n9798 = n9790 & n31718 ;
  assign n31719 = ~n9790 ;
  assign n9800 = n31719 & n9797 ;
  assign n9801 = n9798 | n9800 ;
  assign n9745 = n9496 & n9744 ;
  assign n9802 = n9496 | n9744 ;
  assign n31720 = ~n9745 ;
  assign n9803 = n31720 & n9802 ;
  assign n8175 = n30238 & n8157 ;
  assign n1340 = n740 & n30082 ;
  assign n8213 = n1445 & n8195 ;
  assign n9804 = n1340 | n8213 ;
  assign n9805 = n1219 & n9052 ;
  assign n9806 = n9804 | n9805 ;
  assign n9807 = n8175 | n9806 ;
  assign n9808 = x5 | n9807 ;
  assign n9809 = x5 & n9807 ;
  assign n31721 = ~n9809 ;
  assign n9810 = n9808 & n31721 ;
  assign n9811 = n9803 & n9810 ;
  assign n31722 = ~n9747 ;
  assign n9756 = n31722 & n9755 ;
  assign n9812 = n9756 | n9757 ;
  assign n8189 = n30203 & n8157 ;
  assign n8216 = n1556 & n8195 ;
  assign n9055 = n30082 & n9052 ;
  assign n9813 = n8216 | n9055 ;
  assign n9814 = n740 & n1445 ;
  assign n9815 = n9813 | n9814 ;
  assign n9816 = n8189 | n9815 ;
  assign n9817 = x5 | n9816 ;
  assign n9818 = x5 & n9816 ;
  assign n31723 = ~n9818 ;
  assign n9819 = n9817 & n31723 ;
  assign n9821 = n9812 | n9819 ;
  assign n31724 = ~n9812 ;
  assign n9820 = n31724 & n9819 ;
  assign n31725 = ~n9819 ;
  assign n9822 = n9812 & n31725 ;
  assign n9823 = n9820 | n9822 ;
  assign n31726 = ~n9327 ;
  assign n9492 = n31726 & n9491 ;
  assign n9824 = n9492 | n9493 ;
  assign n8191 = n30209 & n8157 ;
  assign n1561 = n740 & n1556 ;
  assign n8210 = n30196 & n8195 ;
  assign n9825 = n1561 | n8210 ;
  assign n9826 = n1445 & n9052 ;
  assign n9827 = n9825 | n9826 ;
  assign n9828 = n8191 | n9827 ;
  assign n31727 = ~n9828 ;
  assign n9829 = x5 & n31727 ;
  assign n9830 = n30053 & n9828 ;
  assign n9831 = n9829 | n9830 ;
  assign n9832 = n9824 | n9831 ;
  assign n9833 = n9824 & n9831 ;
  assign n31728 = ~n9833 ;
  assign n9834 = n9832 & n31728 ;
  assign n31729 = ~n9342 ;
  assign n9835 = n31729 & n9489 ;
  assign n9836 = n9490 | n9835 ;
  assign n8192 = n3307 & n8157 ;
  assign n8197 = n30105 & n8195 ;
  assign n9060 = n1556 & n9052 ;
  assign n9837 = n8197 | n9060 ;
  assign n9838 = n740 & n30196 ;
  assign n9839 = n9837 | n9838 ;
  assign n9840 = n8192 | n9839 ;
  assign n9841 = x5 | n9840 ;
  assign n9842 = x5 & n9840 ;
  assign n31730 = ~n9842 ;
  assign n9843 = n9841 & n31730 ;
  assign n9845 = n9836 | n9843 ;
  assign n31731 = ~n9836 ;
  assign n9844 = n31731 & n9843 ;
  assign n31732 = ~n9843 ;
  assign n9846 = n9836 & n31732 ;
  assign n9847 = n9844 | n9846 ;
  assign n31733 = ~n9361 ;
  assign n9479 = n31733 & n9478 ;
  assign n9848 = n9479 | n9480 ;
  assign n8183 = n4230 & n8157 ;
  assign n1814 = n740 & n1812 ;
  assign n9054 = n30105 & n9052 ;
  assign n9849 = n1814 | n9054 ;
  assign n9850 = n30108 & n8195 ;
  assign n9851 = n9849 | n9850 ;
  assign n9852 = n8183 | n9851 ;
  assign n9853 = x5 | n9852 ;
  assign n9854 = x5 & n9852 ;
  assign n31734 = ~n9854 ;
  assign n9855 = n9853 & n31734 ;
  assign n9857 = n9848 | n9855 ;
  assign n31735 = ~n9848 ;
  assign n9856 = n31735 & n9855 ;
  assign n31736 = ~n9855 ;
  assign n9858 = n9848 & n31736 ;
  assign n9859 = n9856 | n9858 ;
  assign n31737 = ~n9373 ;
  assign n9860 = n31737 & n9476 ;
  assign n9861 = n9477 | n9860 ;
  assign n8171 = n3592 & n8157 ;
  assign n8218 = n30114 & n8195 ;
  assign n9053 = n1812 & n9052 ;
  assign n9862 = n8218 | n9053 ;
  assign n9863 = n740 & n30108 ;
  assign n9864 = n9862 | n9863 ;
  assign n9865 = n8171 | n9864 ;
  assign n9866 = x5 | n9865 ;
  assign n9867 = x5 & n9865 ;
  assign n31738 = ~n9867 ;
  assign n9868 = n9866 & n31738 ;
  assign n9870 = n9861 & n9868 ;
  assign n31739 = ~n9861 ;
  assign n9869 = n31739 & n9868 ;
  assign n31740 = ~n9868 ;
  assign n9871 = n9861 & n31740 ;
  assign n9872 = n9869 | n9871 ;
  assign n31741 = ~n9386 ;
  assign n9474 = n31741 & n9473 ;
  assign n9873 = n9474 | n9475 ;
  assign n8170 = n30310 & n8157 ;
  assign n1960 = n740 & n30114 ;
  assign n8215 = n30123 & n8195 ;
  assign n9874 = n1960 | n8215 ;
  assign n9875 = n30108 & n9052 ;
  assign n9876 = n9874 | n9875 ;
  assign n9877 = n8170 | n9876 ;
  assign n9878 = x5 | n9877 ;
  assign n9879 = x5 & n9877 ;
  assign n31742 = ~n9879 ;
  assign n9880 = n9878 & n31742 ;
  assign n9882 = n9873 | n9880 ;
  assign n31743 = ~n9873 ;
  assign n9881 = n31743 & n9880 ;
  assign n31744 = ~n9880 ;
  assign n9883 = n9873 & n31744 ;
  assign n9884 = n9881 | n9883 ;
  assign n31745 = ~n9471 ;
  assign n9885 = n9470 & n31745 ;
  assign n9886 = n9472 | n9885 ;
  assign n8194 = n5251 & n8157 ;
  assign n2061 = n740 & n30123 ;
  assign n9068 = n30114 & n9052 ;
  assign n9887 = n2061 | n9068 ;
  assign n9888 = n2102 & n8195 ;
  assign n9889 = n9887 | n9888 ;
  assign n9890 = n8194 | n9889 ;
  assign n31746 = ~n9890 ;
  assign n9891 = x5 & n31746 ;
  assign n9892 = n30053 & n9890 ;
  assign n9893 = n9891 | n9892 ;
  assign n9895 = n9886 | n9893 ;
  assign n31747 = ~n9893 ;
  assign n9894 = n9886 & n31747 ;
  assign n31748 = ~n9886 ;
  assign n9896 = n31748 & n9893 ;
  assign n9897 = n9894 | n9896 ;
  assign n31749 = ~n9413 ;
  assign n9468 = n31749 & n9467 ;
  assign n9898 = n9468 | n9469 ;
  assign n8184 = n30440 & n8157 ;
  assign n8200 = n2216 & n8195 ;
  assign n9069 = n30123 & n9052 ;
  assign n9899 = n8200 | n9069 ;
  assign n9900 = n740 & n2102 ;
  assign n9901 = n9899 | n9900 ;
  assign n9902 = n8184 | n9901 ;
  assign n9903 = x5 | n9902 ;
  assign n9904 = x5 & n9902 ;
  assign n31750 = ~n9904 ;
  assign n9905 = n9903 & n31750 ;
  assign n9907 = n9898 | n9905 ;
  assign n9906 = n9898 & n9905 ;
  assign n31751 = ~n9465 ;
  assign n9908 = n9464 & n31751 ;
  assign n9909 = n9466 | n9908 ;
  assign n8193 = n4352 & n8157 ;
  assign n2221 = n740 & n2216 ;
  assign n8204 = n2295 & n8195 ;
  assign n9910 = n2221 | n8204 ;
  assign n9911 = n2102 & n9052 ;
  assign n9912 = n9910 | n9911 ;
  assign n9913 = n8193 | n9912 ;
  assign n9914 = x5 | n9913 ;
  assign n9915 = x5 & n9913 ;
  assign n31752 = ~n9915 ;
  assign n9916 = n9914 & n31752 ;
  assign n9918 = n9909 | n9916 ;
  assign n31753 = ~n9909 ;
  assign n9917 = n31753 & n9916 ;
  assign n31754 = ~n9916 ;
  assign n9919 = n9909 & n31754 ;
  assign n9920 = n9917 | n9919 ;
  assign n9462 = n9459 & n9461 ;
  assign n9921 = n9459 | n9461 ;
  assign n31755 = ~n9462 ;
  assign n9922 = n31755 & n9921 ;
  assign n8188 = n30444 & n8157 ;
  assign n2296 = n740 & n2295 ;
  assign n8214 = n30445 & n8195 ;
  assign n9923 = n2296 | n8214 ;
  assign n9924 = n2216 & n9052 ;
  assign n9925 = n9923 | n9924 ;
  assign n9926 = n8188 | n9925 ;
  assign n9927 = x5 | n9926 ;
  assign n9928 = x5 & n9926 ;
  assign n31756 = ~n9928 ;
  assign n9929 = n9927 & n31756 ;
  assign n9931 = n9922 | n9929 ;
  assign n31757 = ~n9922 ;
  assign n9930 = n31757 & n9929 ;
  assign n31758 = ~n9929 ;
  assign n9932 = n9922 & n31758 ;
  assign n9933 = n9930 | n9932 ;
  assign n31759 = ~n8911 ;
  assign n9450 = n31759 & n9449 ;
  assign n31760 = ~n9449 ;
  assign n9934 = n8911 & n31760 ;
  assign n9935 = n9450 | n9934 ;
  assign n31761 = ~n9458 ;
  assign n9936 = n31761 & n9935 ;
  assign n31762 = ~n9935 ;
  assign n9937 = n9458 & n31762 ;
  assign n9938 = n9936 | n9937 ;
  assign n8158 = n5392 & n8157 ;
  assign n8201 = n30157 & n8195 ;
  assign n9070 = n2295 & n9052 ;
  assign n9939 = n8201 | n9070 ;
  assign n9940 = n740 & n30445 ;
  assign n9941 = n9939 | n9940 ;
  assign n9942 = n8158 | n9941 ;
  assign n9943 = x5 | n9942 ;
  assign n9944 = x5 & n9942 ;
  assign n31763 = ~n9944 ;
  assign n9945 = n9943 & n31763 ;
  assign n9947 = n9938 | n9945 ;
  assign n9946 = n9938 & n9945 ;
  assign n9948 = n9443 & n9447 ;
  assign n31764 = ~n9948 ;
  assign n9949 = n9448 & n31764 ;
  assign n8165 = n30452 & n8157 ;
  assign n2783 = n740 & n30157 ;
  assign n9071 = n30445 & n9052 ;
  assign n9950 = n2783 | n9071 ;
  assign n9951 = n30453 & n8195 ;
  assign n9952 = n9950 | n9951 ;
  assign n9953 = n8165 | n9952 ;
  assign n9954 = x5 | n9953 ;
  assign n9955 = x5 & n9953 ;
  assign n31765 = ~n9955 ;
  assign n9956 = n9954 & n31765 ;
  assign n9958 = n9949 | n9956 ;
  assign n31766 = ~n9440 ;
  assign n9441 = n9436 & n31766 ;
  assign n31767 = ~n9436 ;
  assign n9959 = n31767 & n9440 ;
  assign n9960 = n9441 | n9959 ;
  assign n8164 = n30458 & n8157 ;
  assign n8219 = n2639 & n8195 ;
  assign n9058 = n30157 & n9052 ;
  assign n9961 = n8219 | n9058 ;
  assign n9962 = n740 & n30453 ;
  assign n9963 = n9961 | n9962 ;
  assign n9964 = n8164 | n9963 ;
  assign n9965 = x5 | n9964 ;
  assign n9966 = x5 & n9964 ;
  assign n31768 = ~n9966 ;
  assign n9967 = n9965 & n31768 ;
  assign n9968 = n9960 & n9967 ;
  assign n9969 = x5 & n738 ;
  assign n9970 = n30463 & n9969 ;
  assign n8172 = n6573 & n8157 ;
  assign n9971 = n740 & n30463 ;
  assign n9972 = n30155 & n9052 ;
  assign n9973 = n9971 | n9972 ;
  assign n9974 = n8172 | n9973 ;
  assign n9976 = n9970 | n9974 ;
  assign n9977 = x5 & n9976 ;
  assign n8181 = n5567 & n8157 ;
  assign n2791 = n740 & n30155 ;
  assign n9056 = n2639 & n9052 ;
  assign n9978 = n2791 | n9056 ;
  assign n9979 = n30463 & n8195 ;
  assign n9980 = n9978 | n9979 ;
  assign n9981 = n8181 | n9980 ;
  assign n9982 = n9977 | n9981 ;
  assign n31769 = ~n9982 ;
  assign n9983 = x5 & n31769 ;
  assign n9985 = n9435 | n9983 ;
  assign n8161 = n5631 & n8157 ;
  assign n8222 = n30155 & n8195 ;
  assign n9073 = n30453 & n9052 ;
  assign n9986 = n8222 | n9073 ;
  assign n9987 = n740 & n2639 ;
  assign n9988 = n9986 | n9987 ;
  assign n9989 = n8161 | n9988 ;
  assign n31770 = ~n9989 ;
  assign n9990 = x5 & n31770 ;
  assign n9991 = n30053 & n9989 ;
  assign n9992 = n9990 | n9991 ;
  assign n9993 = n9985 & n9992 ;
  assign n9994 = n9960 | n9967 ;
  assign n31771 = ~n9968 ;
  assign n9995 = n31771 & n9994 ;
  assign n9996 = n9993 & n9995 ;
  assign n9997 = n9968 | n9996 ;
  assign n9957 = n9949 & n9956 ;
  assign n31772 = ~n9957 ;
  assign n9998 = n31772 & n9958 ;
  assign n31773 = ~n9997 ;
  assign n9999 = n31773 & n9998 ;
  assign n31774 = ~n9999 ;
  assign n10000 = n9958 & n31774 ;
  assign n10001 = n9946 | n10000 ;
  assign n10002 = n9947 & n10001 ;
  assign n31775 = ~n10002 ;
  assign n10003 = n9933 & n31775 ;
  assign n31776 = ~n10003 ;
  assign n10004 = n9931 & n31776 ;
  assign n31777 = ~n10004 ;
  assign n10006 = n9920 & n31777 ;
  assign n31778 = ~n10006 ;
  assign n10007 = n9918 & n31778 ;
  assign n10008 = n9906 | n10007 ;
  assign n10009 = n9907 & n10008 ;
  assign n31779 = ~n10009 ;
  assign n10011 = n9897 & n31779 ;
  assign n31780 = ~n10011 ;
  assign n10012 = n9895 & n31780 ;
  assign n31781 = ~n10012 ;
  assign n10013 = n9884 & n31781 ;
  assign n31782 = ~n10013 ;
  assign n10014 = n9882 & n31782 ;
  assign n10015 = n9872 & n10014 ;
  assign n10016 = n9870 | n10015 ;
  assign n31783 = ~n10016 ;
  assign n10017 = n9859 & n31783 ;
  assign n31784 = ~n10017 ;
  assign n10018 = n9857 & n31784 ;
  assign n8163 = n30233 & n8157 ;
  assign n8209 = n1812 & n8195 ;
  assign n9067 = n30196 & n9052 ;
  assign n10019 = n8209 | n9067 ;
  assign n10020 = n740 & n30105 ;
  assign n10021 = n10019 | n10020 ;
  assign n10022 = n8163 | n10021 ;
  assign n10023 = x5 | n10022 ;
  assign n10024 = x5 & n10022 ;
  assign n31785 = ~n10024 ;
  assign n10025 = n10023 & n31785 ;
  assign n10027 = n10018 | n10025 ;
  assign n31786 = ~n9485 ;
  assign n9488 = n31786 & n9486 ;
  assign n31787 = ~n9486 ;
  assign n10028 = n9485 & n31787 ;
  assign n10029 = n9488 | n10028 ;
  assign n10026 = n10018 & n10025 ;
  assign n31788 = ~n10026 ;
  assign n10030 = n31788 & n10027 ;
  assign n31789 = ~n10029 ;
  assign n10031 = n31789 & n10030 ;
  assign n31790 = ~n10031 ;
  assign n10032 = n10027 & n31790 ;
  assign n31791 = ~n10032 ;
  assign n10034 = n9847 & n31791 ;
  assign n31792 = ~n10034 ;
  assign n10035 = n9845 & n31792 ;
  assign n31793 = ~n10035 ;
  assign n10036 = n9834 & n31793 ;
  assign n31794 = ~n10036 ;
  assign n10037 = n9832 & n31794 ;
  assign n31795 = ~n10037 ;
  assign n10039 = n9823 & n31795 ;
  assign n31796 = ~n10039 ;
  assign n10040 = n9821 & n31796 ;
  assign n10041 = n9803 | n9810 ;
  assign n10042 = n10040 & n10041 ;
  assign n10043 = n9811 | n10042 ;
  assign n31797 = ~n10043 ;
  assign n10045 = n9801 & n31797 ;
  assign n31798 = ~n10045 ;
  assign n10046 = n9799 & n31798 ;
  assign n10047 = n9780 | n9787 ;
  assign n10048 = n10046 & n10047 ;
  assign n10049 = n9788 | n10048 ;
  assign n31799 = ~n10049 ;
  assign n10051 = n9779 & n31799 ;
  assign n31800 = ~n10051 ;
  assign n10052 = n9777 & n31800 ;
  assign n31801 = ~n10052 ;
  assign n10053 = n9732 & n31801 ;
  assign n31802 = ~n10053 ;
  assign n10054 = n9730 & n31802 ;
  assign n31803 = ~n10054 ;
  assign n10056 = n9720 & n31803 ;
  assign n31804 = ~n10056 ;
  assign n10057 = n9718 & n31804 ;
  assign n10058 = n9706 & n10057 ;
  assign n10059 = n9707 | n10058 ;
  assign n10060 = n9689 | n9696 ;
  assign n31805 = ~n9697 ;
  assign n10061 = n31805 & n10060 ;
  assign n10062 = n10059 & n10061 ;
  assign n10063 = n9697 | n10062 ;
  assign n31806 = ~n10063 ;
  assign n10064 = n9687 & n31806 ;
  assign n31807 = ~n10064 ;
  assign n10065 = n9685 & n31807 ;
  assign n10066 = n9674 & n10065 ;
  assign n31808 = ~n9177 ;
  assign n10067 = n31808 & n9518 ;
  assign n10068 = n9519 | n10067 ;
  assign n10069 = n9674 | n10065 ;
  assign n31809 = ~n10066 ;
  assign n10070 = n31809 & n10069 ;
  assign n10071 = n10068 & n10070 ;
  assign n10072 = n10066 | n10071 ;
  assign n10073 = n9659 & n9666 ;
  assign n31810 = ~n10073 ;
  assign n10074 = n9667 & n31810 ;
  assign n31811 = ~n10072 ;
  assign n10075 = n31811 & n10074 ;
  assign n31812 = ~n10075 ;
  assign n10076 = n9667 & n31812 ;
  assign n31813 = ~n9657 ;
  assign n10077 = n31813 & n10076 ;
  assign n8160 = n30385 & n8157 ;
  assign n8217 = n30361 & n8195 ;
  assign n9072 = n4811 & n9052 ;
  assign n10078 = n8217 | n9072 ;
  assign n10079 = n740 & n4664 ;
  assign n10080 = n10078 | n10079 ;
  assign n10081 = n8160 | n10080 ;
  assign n10082 = x5 | n10081 ;
  assign n10083 = x5 & n10081 ;
  assign n31814 = ~n10083 ;
  assign n10084 = n10082 & n31814 ;
  assign n31815 = ~n10076 ;
  assign n10085 = n9657 & n31815 ;
  assign n10086 = n10077 | n10085 ;
  assign n31816 = ~n10086 ;
  assign n10087 = n10084 & n31816 ;
  assign n10088 = n10077 | n10087 ;
  assign n10090 = n9655 | n10088 ;
  assign n31817 = ~n9653 ;
  assign n10091 = n31817 & n10090 ;
  assign n31818 = ~n10091 ;
  assign n10093 = n9643 & n31818 ;
  assign n31819 = ~n10093 ;
  assign n10094 = n9641 & n31819 ;
  assign n10096 = n9631 | n10094 ;
  assign n31820 = ~n9630 ;
  assign n10097 = n31820 & n10096 ;
  assign n31821 = ~n10097 ;
  assign n10099 = n9619 & n31821 ;
  assign n31822 = ~n10099 ;
  assign n10100 = n9617 & n31822 ;
  assign n10102 = n9608 | n10100 ;
  assign n31823 = ~n10088 ;
  assign n10089 = n9655 & n31823 ;
  assign n31824 = ~n9655 ;
  assign n10103 = n31824 & n10088 ;
  assign n10104 = n10089 | n10103 ;
  assign n31825 = ~n9561 ;
  assign n10105 = x0 & n31825 ;
  assign n10115 = n30530 & n10105 ;
  assign n31826 = ~x0 ;
  assign n10126 = n31826 & x1 ;
  assign n10138 = n30415 & n10126 ;
  assign n10148 = n10115 | n10138 ;
  assign n10149 = n6411 & n9562 ;
  assign n10150 = n10148 | n10149 ;
  assign n10151 = n30049 & n10150 ;
  assign n5022 = n31643 & n5017 ;
  assign n31827 = ~n5022 ;
  assign n10152 = x2 & n31827 ;
  assign n31828 = ~n10150 ;
  assign n10153 = n31828 & n10152 ;
  assign n10154 = n10151 | n10153 ;
  assign n31829 = ~n10154 ;
  assign n10156 = n10104 & n31829 ;
  assign n31830 = ~n10074 ;
  assign n10157 = n10072 & n31830 ;
  assign n10158 = n10075 | n10157 ;
  assign n10107 = n5017 & n10105 ;
  assign n10145 = n30405 & n10126 ;
  assign n10159 = n10107 | n10145 ;
  assign n10160 = n30512 & n9562 ;
  assign n10161 = n10159 | n10160 ;
  assign n10162 = n30049 & n10161 ;
  assign n4820 = n31643 & n4811 ;
  assign n31831 = ~n4820 ;
  assign n10163 = x2 & n31831 ;
  assign n31832 = ~n10161 ;
  assign n10164 = n31832 & n10163 ;
  assign n10165 = n10162 | n10164 ;
  assign n10166 = n10158 & n10165 ;
  assign n10167 = n10158 | n10165 ;
  assign n10168 = n10068 | n10070 ;
  assign n31833 = ~n10071 ;
  assign n10169 = n31833 & n10168 ;
  assign n10117 = n30405 & n10105 ;
  assign n10134 = n4811 & n10126 ;
  assign n10170 = n10117 | n10134 ;
  assign n10171 = n30578 & n9562 ;
  assign n10172 = n10170 | n10171 ;
  assign n10173 = x2 & n10172 ;
  assign n10174 = n31643 & n4664 ;
  assign n31834 = ~n10174 ;
  assign n10175 = x2 & n31834 ;
  assign n10176 = n10172 | n10175 ;
  assign n31835 = ~n10173 ;
  assign n10177 = n31835 & n10176 ;
  assign n10179 = n10169 & n10177 ;
  assign n10178 = n10169 | n10177 ;
  assign n31836 = ~n9687 ;
  assign n10180 = n31836 & n10063 ;
  assign n10181 = n10064 | n10180 ;
  assign n9555 = n30361 & n9552 ;
  assign n9575 = n30385 & n9562 ;
  assign n10182 = n4811 & n10105 ;
  assign n10183 = n4664 & n10126 ;
  assign n10184 = n10182 | n10183 ;
  assign n10185 = n9575 | n10184 ;
  assign n31837 = ~n10185 ;
  assign n10186 = x2 & n31837 ;
  assign n10187 = n30049 & n10185 ;
  assign n10188 = n10186 | n10187 ;
  assign n31838 = ~n9555 ;
  assign n10189 = n31838 & n10188 ;
  assign n10190 = n10181 & n10189 ;
  assign n10191 = n10181 | n10189 ;
  assign n10192 = n10059 | n10061 ;
  assign n31839 = ~n10062 ;
  assign n10193 = n31839 & n10192 ;
  assign n9564 = n4674 & n9562 ;
  assign n10125 = n4664 & n10105 ;
  assign n10141 = n30361 & n10126 ;
  assign n10194 = n10125 | n10141 ;
  assign n10195 = n9564 | n10194 ;
  assign n10196 = n30049 & n10195 ;
  assign n3943 = n733 | n3938 ;
  assign n10197 = x2 & n3943 ;
  assign n31840 = ~n10195 ;
  assign n10198 = n31840 & n10197 ;
  assign n10199 = n10196 | n10198 ;
  assign n10200 = n10193 & n10199 ;
  assign n10201 = n10193 | n10199 ;
  assign n31841 = ~n9707 ;
  assign n10202 = n9706 & n31841 ;
  assign n31842 = ~n10057 ;
  assign n10203 = n31842 & n10202 ;
  assign n31843 = ~n10202 ;
  assign n10204 = n10057 & n31843 ;
  assign n10205 = n10203 | n10204 ;
  assign n9576 = n5723 & n9562 ;
  assign n10119 = n30361 & n10105 ;
  assign n10139 = n30282 & n10126 ;
  assign n10206 = n10119 | n10139 ;
  assign n10207 = n9576 | n10206 ;
  assign n10208 = x2 & n10207 ;
  assign n10209 = n31643 & n4033 ;
  assign n31844 = ~n10209 ;
  assign n10210 = x2 & n31844 ;
  assign n10211 = n10207 | n10210 ;
  assign n31845 = ~n10208 ;
  assign n10212 = n31845 & n10211 ;
  assign n10213 = n10205 | n10212 ;
  assign n10214 = n10205 & n10212 ;
  assign n31846 = ~n9720 ;
  assign n10055 = n31846 & n10054 ;
  assign n10215 = n10055 | n10056 ;
  assign n10120 = n30282 & n10105 ;
  assign n10131 = n4033 & n10126 ;
  assign n10216 = n10120 | n10131 ;
  assign n10217 = n30286 & n9562 ;
  assign n10218 = n10216 | n10217 ;
  assign n10219 = n30049 & n10218 ;
  assign n4096 = n31643 & n4093 ;
  assign n31847 = ~n4096 ;
  assign n10220 = x2 & n31847 ;
  assign n31848 = ~n10218 ;
  assign n10221 = n31848 & n10220 ;
  assign n10222 = n10219 | n10221 ;
  assign n10223 = n10215 & n10222 ;
  assign n10224 = n10215 | n10222 ;
  assign n31849 = ~n9732 ;
  assign n10225 = n31849 & n10052 ;
  assign n10226 = n10053 | n10225 ;
  assign n10116 = n4033 & n10105 ;
  assign n10144 = n4093 & n10126 ;
  assign n10227 = n10116 | n10144 ;
  assign n10228 = n4442 & n9562 ;
  assign n10229 = n10227 | n10228 ;
  assign n10230 = x2 & n10229 ;
  assign n10231 = n733 | n3863 ;
  assign n10232 = x2 & n10231 ;
  assign n10233 = n10229 | n10232 ;
  assign n31850 = ~n10230 ;
  assign n10234 = n31850 & n10233 ;
  assign n10235 = n10226 & n10234 ;
  assign n10236 = n10226 | n10234 ;
  assign n31851 = ~n9779 ;
  assign n10050 = n31851 & n10049 ;
  assign n10533 = n10050 | n10051 ;
  assign n9566 = n30349 & n9562 ;
  assign n10534 = n4093 & n10105 ;
  assign n10535 = n30264 & n10126 ;
  assign n10536 = n10534 | n10535 ;
  assign n10537 = n9566 | n10536 ;
  assign n10538 = n30049 & n10537 ;
  assign n3703 = n31643 & n3700 ;
  assign n31852 = ~n3703 ;
  assign n10540 = x2 & n31852 ;
  assign n31853 = ~n10537 ;
  assign n10541 = n31853 & n10540 ;
  assign n10542 = n10538 | n10541 ;
  assign n10548 = n10533 | n10542 ;
  assign n31854 = ~n9788 ;
  assign n10237 = n31854 & n10047 ;
  assign n31855 = ~n10046 ;
  assign n10238 = n31855 & n10237 ;
  assign n31856 = ~n10237 ;
  assign n10239 = n10046 & n31856 ;
  assign n10240 = n10238 | n10239 ;
  assign n9572 = n30263 & n9562 ;
  assign n10241 = n30264 & n10105 ;
  assign n10242 = n3700 & n10126 ;
  assign n10243 = n10241 | n10242 ;
  assign n10244 = n9572 | n10243 ;
  assign n10245 = x2 & n10244 ;
  assign n10246 = n31643 & n3764 ;
  assign n31857 = ~n10246 ;
  assign n10247 = x2 & n31857 ;
  assign n10248 = n10244 | n10247 ;
  assign n31858 = ~n10245 ;
  assign n10249 = n31858 & n10248 ;
  assign n10250 = n10240 | n10249 ;
  assign n31859 = ~n9811 ;
  assign n10251 = n31859 & n10041 ;
  assign n31860 = ~n10040 ;
  assign n10252 = n31860 & n10251 ;
  assign n31861 = ~n10251 ;
  assign n10253 = n10040 & n31861 ;
  assign n10254 = n10252 | n10253 ;
  assign n31862 = ~n9823 ;
  assign n10038 = n31862 & n10037 ;
  assign n10255 = n10038 | n10039 ;
  assign n10118 = n1074 & n10105 ;
  assign n10147 = n30074 & n10126 ;
  assign n10257 = n10118 | n10147 ;
  assign n2843 = n1082 & n2841 ;
  assign n31863 = ~n2843 ;
  assign n10256 = n31863 & n3780 ;
  assign n31864 = ~n10256 ;
  assign n10258 = n9562 & n31864 ;
  assign n10259 = n10257 | n10258 ;
  assign n10260 = n30049 & n10259 ;
  assign n1224 = n31643 & n1219 ;
  assign n31865 = ~n1224 ;
  assign n10261 = x2 & n31865 ;
  assign n31866 = ~n10259 ;
  assign n10262 = n31866 & n10261 ;
  assign n10263 = n10260 | n10262 ;
  assign n10264 = n10255 & n10263 ;
  assign n10265 = n10255 | n10263 ;
  assign n31867 = ~n9834 ;
  assign n10266 = n31867 & n10035 ;
  assign n10267 = n10036 | n10266 ;
  assign n10121 = n30074 & n10105 ;
  assign n10142 = n1219 & n10126 ;
  assign n10269 = n10121 | n10142 ;
  assign n3394 = n1226 & n2839 ;
  assign n31868 = ~n3394 ;
  assign n10268 = n2840 & n31868 ;
  assign n31869 = ~n10268 ;
  assign n10270 = n9562 & n31869 ;
  assign n10271 = n10269 | n10270 ;
  assign n10272 = n30049 & n10271 ;
  assign n1341 = n733 | n1336 ;
  assign n10273 = x2 & n1341 ;
  assign n31870 = ~n10271 ;
  assign n10274 = n31870 & n10273 ;
  assign n10275 = n10272 | n10274 ;
  assign n10276 = n10267 & n10275 ;
  assign n10277 = n10267 | n10275 ;
  assign n31871 = ~n9847 ;
  assign n10033 = n31871 & n10032 ;
  assign n10278 = n10033 | n10034 ;
  assign n10122 = n1219 & n10105 ;
  assign n10128 = n30082 & n10126 ;
  assign n10280 = n10122 | n10128 ;
  assign n2837 = n1343 & n2835 ;
  assign n31872 = ~n2837 ;
  assign n10279 = n31872 & n2838 ;
  assign n31873 = ~n10279 ;
  assign n10281 = n9562 & n31873 ;
  assign n10282 = n10280 | n10281 ;
  assign n10283 = n30049 & n10282 ;
  assign n1447 = n31643 & n1445 ;
  assign n31874 = ~n1447 ;
  assign n10284 = x2 & n31874 ;
  assign n31875 = ~n10282 ;
  assign n10285 = n31875 & n10284 ;
  assign n10286 = n10283 | n10285 ;
  assign n10287 = n10278 & n10286 ;
  assign n10288 = n10278 | n10286 ;
  assign n9577 = n30203 & n9562 ;
  assign n9557 = n1556 & n9552 ;
  assign n10123 = n30082 & n10105 ;
  assign n10289 = n9557 | n10123 ;
  assign n10290 = n1445 & n10126 ;
  assign n10291 = n10289 | n10290 ;
  assign n10292 = n9577 | n10291 ;
  assign n31876 = ~n10292 ;
  assign n10293 = x2 & n31876 ;
  assign n10295 = n30049 & n10292 ;
  assign n10296 = n10293 | n10295 ;
  assign n31877 = ~n10030 ;
  assign n10297 = n10029 & n31877 ;
  assign n10298 = n10031 | n10297 ;
  assign n10499 = n10296 & n10298 ;
  assign n31878 = ~n9859 ;
  assign n10299 = n31878 & n10016 ;
  assign n10300 = n10017 | n10299 ;
  assign n10301 = n9872 | n10014 ;
  assign n31879 = ~n10015 ;
  assign n10302 = n31879 & n10301 ;
  assign n10106 = n1556 & n10105 ;
  assign n10143 = n30196 & n10126 ;
  assign n10304 = n10106 | n10143 ;
  assign n31880 = ~n2828 ;
  assign n3305 = n1678 & n31880 ;
  assign n10303 = n2829 | n3305 ;
  assign n10305 = n9562 & n10303 ;
  assign n10306 = n10304 | n10305 ;
  assign n10307 = n30049 & n10306 ;
  assign n1754 = n733 | n1752 ;
  assign n10308 = x2 & n1754 ;
  assign n31881 = ~n10306 ;
  assign n10309 = n31881 & n10308 ;
  assign n10310 = n10307 | n10309 ;
  assign n10311 = n10302 & n10310 ;
  assign n10312 = n10302 | n10310 ;
  assign n31882 = ~n9884 ;
  assign n10313 = n31882 & n10012 ;
  assign n10314 = n10013 | n10313 ;
  assign n10113 = n30196 & n10105 ;
  assign n10132 = n30105 & n10126 ;
  assign n10316 = n10113 | n10132 ;
  assign n2826 = n1757 | n2824 ;
  assign n31883 = ~n2827 ;
  assign n10315 = n2826 & n31883 ;
  assign n31884 = ~n10315 ;
  assign n10317 = n9562 & n31884 ;
  assign n10318 = n10316 | n10317 ;
  assign n10319 = x2 & n10318 ;
  assign n1817 = n31643 & n1812 ;
  assign n31885 = ~n1817 ;
  assign n10320 = x2 & n31885 ;
  assign n10321 = n10318 | n10320 ;
  assign n31886 = ~n10319 ;
  assign n10322 = n31886 & n10321 ;
  assign n10324 = n10314 & n10322 ;
  assign n31887 = ~n9897 ;
  assign n10010 = n31887 & n10009 ;
  assign n10325 = n10010 | n10011 ;
  assign n9563 = n4230 & n9562 ;
  assign n10326 = n30105 & n10105 ;
  assign n10327 = n1812 & n10126 ;
  assign n10328 = n10326 | n10327 ;
  assign n10329 = n9563 | n10328 ;
  assign n10330 = x2 | n10329 ;
  assign n10331 = x2 & n10329 ;
  assign n31888 = ~n10331 ;
  assign n10332 = n10330 & n31888 ;
  assign n10333 = n30108 & n9552 ;
  assign n31889 = ~n10333 ;
  assign n10334 = n10332 & n31889 ;
  assign n10478 = n10325 & n10334 ;
  assign n31890 = ~n9906 ;
  assign n10336 = n31890 & n9907 ;
  assign n31891 = ~n10007 ;
  assign n10337 = n31891 & n10336 ;
  assign n31892 = ~n10336 ;
  assign n10338 = n10007 & n31892 ;
  assign n10339 = n10337 | n10338 ;
  assign n10112 = n1812 & n10105 ;
  assign n10136 = n30108 & n10126 ;
  assign n10341 = n10112 | n10136 ;
  assign n31893 = ~n2818 ;
  assign n2820 = n1891 & n31893 ;
  assign n10340 = n2820 | n2821 ;
  assign n10342 = n9562 & n10340 ;
  assign n10343 = n10341 | n10342 ;
  assign n10344 = x2 & n10343 ;
  assign n1963 = n733 | n1957 ;
  assign n10345 = x2 & n1963 ;
  assign n10346 = n10343 | n10345 ;
  assign n31894 = ~n10344 ;
  assign n10347 = n31894 & n10346 ;
  assign n10348 = n10339 | n10347 ;
  assign n31895 = ~n9920 ;
  assign n10005 = n31895 & n10004 ;
  assign n10349 = n10005 | n10006 ;
  assign n9578 = n30310 & n9562 ;
  assign n9554 = n30123 & n9552 ;
  assign n10135 = n30114 & n10126 ;
  assign n10350 = n9554 | n10135 ;
  assign n10351 = n30108 & n10105 ;
  assign n10352 = n10350 | n10351 ;
  assign n10353 = n9578 | n10352 ;
  assign n31896 = ~n10353 ;
  assign n10354 = x2 & n31896 ;
  assign n10355 = n30049 & n10353 ;
  assign n10356 = n10354 | n10355 ;
  assign n10357 = n10349 | n10356 ;
  assign n31897 = ~n9933 ;
  assign n10358 = n31897 & n10002 ;
  assign n10359 = n10003 | n10358 ;
  assign n9571 = n5251 & n9562 ;
  assign n10360 = n30114 & n10105 ;
  assign n10361 = n30123 & n10126 ;
  assign n10362 = n10360 | n10361 ;
  assign n10363 = n9571 | n10362 ;
  assign n10364 = x2 & n10363 ;
  assign n2107 = n31643 & n2102 ;
  assign n31898 = ~n2107 ;
  assign n10366 = x2 & n31898 ;
  assign n10367 = n10363 | n10366 ;
  assign n31899 = ~n10364 ;
  assign n10368 = n31899 & n10367 ;
  assign n10470 = n10359 & n10368 ;
  assign n31900 = ~n9946 ;
  assign n10369 = n31900 & n9947 ;
  assign n10370 = n10000 & n10369 ;
  assign n10371 = n10000 | n10369 ;
  assign n31901 = ~n10370 ;
  assign n10372 = n31901 & n10371 ;
  assign n9565 = n30440 & n9562 ;
  assign n10373 = n30123 & n10105 ;
  assign n10374 = n2102 & n10126 ;
  assign n10375 = n10373 | n10374 ;
  assign n10376 = n9565 | n10375 ;
  assign n10377 = n30049 & n10376 ;
  assign n2218 = n31643 & n2216 ;
  assign n31902 = ~n2218 ;
  assign n10378 = x2 & n31902 ;
  assign n31903 = ~n10376 ;
  assign n10379 = n31903 & n10378 ;
  assign n10380 = n10377 | n10379 ;
  assign n10381 = n10372 & n10380 ;
  assign n10108 = n2102 & n10105 ;
  assign n10133 = n2216 & n10126 ;
  assign n10382 = n10108 | n10133 ;
  assign n10383 = n4352 & n9562 ;
  assign n10384 = n10382 | n10383 ;
  assign n10385 = x2 & n10384 ;
  assign n9556 = n2295 & n9552 ;
  assign n31904 = ~n9556 ;
  assign n10386 = x2 & n31904 ;
  assign n10387 = n10384 | n10386 ;
  assign n31905 = ~n10385 ;
  assign n10388 = n31905 & n10387 ;
  assign n10389 = n9993 | n9995 ;
  assign n31906 = ~n9996 ;
  assign n10390 = n31906 & n10389 ;
  assign n9568 = n30444 & n9562 ;
  assign n10391 = n2216 & n10105 ;
  assign n10392 = n2295 & n10126 ;
  assign n10393 = n10391 | n10392 ;
  assign n10394 = n9568 | n10393 ;
  assign n10395 = x2 & n10394 ;
  assign n10396 = n30445 & n9552 ;
  assign n31907 = ~n10396 ;
  assign n10397 = x2 & n31907 ;
  assign n10398 = n10394 | n10397 ;
  assign n31908 = ~n10395 ;
  assign n10399 = n31908 & n10398 ;
  assign n10400 = n10390 & n10399 ;
  assign n10401 = n10390 | n10399 ;
  assign n9579 = n30452 & n9562 ;
  assign n9558 = n30453 & n9552 ;
  assign n10137 = n30157 & n10126 ;
  assign n10402 = n9558 | n10137 ;
  assign n10403 = n30445 & n10105 ;
  assign n10404 = n10402 | n10403 ;
  assign n10405 = n9579 | n10404 ;
  assign n31909 = ~n10405 ;
  assign n10406 = x2 & n31909 ;
  assign n10407 = n30049 & n10405 ;
  assign n10408 = n10406 | n10407 ;
  assign n31910 = ~n9974 ;
  assign n9975 = n9970 & n31910 ;
  assign n31911 = ~n9970 ;
  assign n10409 = n31911 & n9974 ;
  assign n10410 = n9975 | n10409 ;
  assign n9553 = n2639 & n9552 ;
  assign n9580 = n30458 & n9562 ;
  assign n10411 = n30157 & n10105 ;
  assign n10412 = n30453 & n10126 ;
  assign n10413 = n10411 | n10412 ;
  assign n10414 = n9580 | n10413 ;
  assign n31912 = ~n10414 ;
  assign n10415 = x2 & n31912 ;
  assign n10416 = n30049 & n10414 ;
  assign n10417 = n10415 | n10416 ;
  assign n31913 = ~n9553 ;
  assign n10418 = n31913 & n10417 ;
  assign n10420 = n10410 & n10418 ;
  assign n10419 = n10410 | n10418 ;
  assign n9570 = n5631 & n9562 ;
  assign n10421 = n30453 & n10105 ;
  assign n10422 = n2639 & n10126 ;
  assign n10423 = n10421 | n10422 ;
  assign n10424 = n9570 | n10423 ;
  assign n2787 = n733 | n2471 ;
  assign n10425 = x2 & n2787 ;
  assign n10426 = n10424 | n10425 ;
  assign n10427 = n738 & n30463 ;
  assign n10428 = x2 & n10424 ;
  assign n31914 = ~n10428 ;
  assign n10429 = n10427 & n31914 ;
  assign n10430 = n10426 & n10429 ;
  assign n10431 = n10419 & n10430 ;
  assign n10432 = n10420 | n10431 ;
  assign n10433 = n10408 | n10432 ;
  assign n10434 = n9977 & n9981 ;
  assign n31915 = ~n10434 ;
  assign n10435 = n9982 & n31915 ;
  assign n10436 = n10433 & n10435 ;
  assign n10437 = n10408 & n10432 ;
  assign n10438 = n10436 | n10437 ;
  assign n31916 = ~n9435 ;
  assign n9984 = n31916 & n9983 ;
  assign n31917 = ~n9983 ;
  assign n10439 = n9435 & n31917 ;
  assign n10440 = n9984 | n10439 ;
  assign n31918 = ~n9992 ;
  assign n10441 = n31918 & n10440 ;
  assign n31919 = ~n10440 ;
  assign n10442 = n9992 & n31919 ;
  assign n10443 = n10441 | n10442 ;
  assign n10444 = n10438 | n10443 ;
  assign n9569 = n5392 & n9562 ;
  assign n10445 = n2295 & n10105 ;
  assign n10446 = n30445 & n10126 ;
  assign n10447 = n10445 | n10446 ;
  assign n10448 = n9569 | n10447 ;
  assign n10449 = x2 & n10448 ;
  assign n2784 = n733 | n2779 ;
  assign n10450 = x2 & n2784 ;
  assign n10451 = n10448 | n10450 ;
  assign n31920 = ~n10449 ;
  assign n10452 = n31920 & n10451 ;
  assign n10453 = n10444 & n10452 ;
  assign n10454 = n10438 & n10443 ;
  assign n10455 = n10453 | n10454 ;
  assign n10456 = n10401 & n10455 ;
  assign n10457 = n10400 | n10456 ;
  assign n10458 = n10388 | n10457 ;
  assign n31921 = ~n9998 ;
  assign n10459 = n9997 & n31921 ;
  assign n10460 = n9999 | n10459 ;
  assign n10461 = n10388 & n10457 ;
  assign n10462 = n10460 | n10461 ;
  assign n10463 = n10458 & n10462 ;
  assign n10464 = n10381 | n10463 ;
  assign n10365 = n30049 & n10363 ;
  assign n31922 = ~n10363 ;
  assign n10465 = n31922 & n10366 ;
  assign n10466 = n10365 | n10465 ;
  assign n10467 = n10359 | n10466 ;
  assign n10468 = n10372 | n10380 ;
  assign n10469 = n10467 & n10468 ;
  assign n10471 = n10464 & n10469 ;
  assign n10472 = n10470 | n10471 ;
  assign n10473 = n10357 & n10472 ;
  assign n10474 = n10339 & n10347 ;
  assign n10475 = n10349 & n10356 ;
  assign n10476 = n10474 | n10475 ;
  assign n10477 = n10473 | n10476 ;
  assign n10479 = n10348 & n10477 ;
  assign n10480 = n10478 | n10479 ;
  assign n10323 = n10314 | n10322 ;
  assign n10335 = n10325 | n10334 ;
  assign n10481 = n10323 & n10335 ;
  assign n10482 = n10480 & n10481 ;
  assign n10483 = n10324 | n10482 ;
  assign n10484 = n10312 & n10483 ;
  assign n10485 = n10311 | n10484 ;
  assign n10486 = n10300 & n10485 ;
  assign n9574 = n30209 & n9562 ;
  assign n10111 = n1445 & n10105 ;
  assign n10130 = n1556 & n10126 ;
  assign n10487 = n10111 | n10130 ;
  assign n10488 = n9574 | n10487 ;
  assign n10489 = n30049 & n10488 ;
  assign n1674 = n733 | n1671 ;
  assign n10490 = x2 & n1674 ;
  assign n31923 = ~n10488 ;
  assign n10491 = n31923 & n10490 ;
  assign n10492 = n10489 | n10491 ;
  assign n10493 = n10486 | n10492 ;
  assign n10294 = x2 | n10292 ;
  assign n10494 = x2 & n10292 ;
  assign n31924 = ~n10494 ;
  assign n10495 = n10294 & n31924 ;
  assign n10496 = n10298 | n10495 ;
  assign n10497 = n10300 | n10485 ;
  assign n10498 = n10496 & n10497 ;
  assign n10500 = n10493 & n10498 ;
  assign n10501 = n10499 | n10500 ;
  assign n10502 = n10288 & n10501 ;
  assign n10503 = n10287 | n10502 ;
  assign n10504 = n10277 & n10503 ;
  assign n10505 = n10276 | n10504 ;
  assign n10506 = n10265 & n10505 ;
  assign n10507 = n10264 | n10506 ;
  assign n10509 = n10254 & n10507 ;
  assign n10508 = n10254 | n10507 ;
  assign n9573 = n4420 & n9562 ;
  assign n10124 = n3764 & n10105 ;
  assign n10140 = n1074 & n10126 ;
  assign n10510 = n10124 | n10140 ;
  assign n10511 = n30074 & n9552 ;
  assign n10512 = n10510 | n10511 ;
  assign n10513 = n9573 | n10512 ;
  assign n31925 = ~n10513 ;
  assign n10514 = x2 & n31925 ;
  assign n10515 = n30049 & n10513 ;
  assign n10516 = n10514 | n10515 ;
  assign n10517 = n10508 & n10516 ;
  assign n10518 = n10509 | n10517 ;
  assign n31926 = ~n9801 ;
  assign n10044 = n31926 & n10043 ;
  assign n10519 = n10044 | n10045 ;
  assign n10520 = n10518 & n10519 ;
  assign n9567 = n3787 & n9562 ;
  assign n10521 = n3700 & n10105 ;
  assign n10522 = n3764 & n10126 ;
  assign n10523 = n10521 | n10522 ;
  assign n10524 = n9567 | n10523 ;
  assign n10525 = n30049 & n10524 ;
  assign n1075 = n31643 & n1074 ;
  assign n31927 = ~n1075 ;
  assign n10526 = x2 & n31927 ;
  assign n31928 = ~n10524 ;
  assign n10527 = n31928 & n10526 ;
  assign n10528 = n10525 | n10527 ;
  assign n10529 = n10518 | n10519 ;
  assign n10530 = n10528 & n10529 ;
  assign n10531 = n10520 | n10530 ;
  assign n10532 = n10250 & n10531 ;
  assign n10545 = n10240 & n10249 ;
  assign n10539 = x2 & n10537 ;
  assign n10543 = n10537 | n10540 ;
  assign n31929 = ~n10539 ;
  assign n10544 = n31929 & n10543 ;
  assign n10546 = n10533 & n10544 ;
  assign n10547 = n10545 | n10546 ;
  assign n10549 = n10532 | n10547 ;
  assign n10550 = n10548 & n10549 ;
  assign n10551 = n10236 & n10550 ;
  assign n10552 = n10235 | n10551 ;
  assign n10553 = n10224 & n10552 ;
  assign n10554 = n10223 | n10553 ;
  assign n10555 = n10214 | n10554 ;
  assign n10556 = n10213 & n10555 ;
  assign n10557 = n10201 & n10556 ;
  assign n10558 = n10200 | n10557 ;
  assign n10559 = n10191 & n10558 ;
  assign n10560 = n10190 | n10559 ;
  assign n10561 = n10178 & n10560 ;
  assign n10562 = n10179 | n10561 ;
  assign n10563 = n10167 & n10562 ;
  assign n10564 = n10166 | n10563 ;
  assign n10114 = n30415 & n10105 ;
  assign n10146 = n5017 & n10126 ;
  assign n10565 = n10114 | n10146 ;
  assign n10566 = n30410 & n9562 ;
  assign n10567 = n10565 | n10566 ;
  assign n10568 = n30049 & n10567 ;
  assign n5111 = n733 | n5105 ;
  assign n10569 = x2 & n5111 ;
  assign n31930 = ~n10567 ;
  assign n10570 = n31930 & n10569 ;
  assign n10571 = n10568 | n10570 ;
  assign n10573 = n10564 | n10571 ;
  assign n10572 = n10564 & n10571 ;
  assign n31931 = ~n10084 ;
  assign n10574 = n31931 & n10086 ;
  assign n10575 = n10087 | n10574 ;
  assign n31932 = ~n10572 ;
  assign n10576 = n31932 & n10575 ;
  assign n31933 = ~n10576 ;
  assign n10577 = n10573 & n31933 ;
  assign n31934 = ~n10104 ;
  assign n10155 = n31934 & n10154 ;
  assign n10578 = n10155 | n10156 ;
  assign n10579 = n10577 | n10578 ;
  assign n31935 = ~n10156 ;
  assign n10580 = n31935 & n10579 ;
  assign n10110 = n30535 & n10105 ;
  assign n10129 = n30530 & n10126 ;
  assign n10581 = n10110 | n10129 ;
  assign n10582 = n30587 & n9562 ;
  assign n10583 = n10581 | n10582 ;
  assign n10584 = n30049 & n10583 ;
  assign n4940 = n733 | n4925 ;
  assign n10585 = x2 & n4940 ;
  assign n31936 = ~n10583 ;
  assign n10586 = n31936 & n10585 ;
  assign n10587 = n10584 | n10586 ;
  assign n10588 = n10580 & n10587 ;
  assign n10092 = n9643 & n10091 ;
  assign n10589 = n9643 | n10091 ;
  assign n31937 = ~n10092 ;
  assign n10590 = n31937 & n10589 ;
  assign n10591 = n10580 | n10587 ;
  assign n31938 = ~n10588 ;
  assign n10592 = n31938 & n10591 ;
  assign n10593 = n10590 & n10592 ;
  assign n10594 = n10588 | n10593 ;
  assign n10109 = n30545 & n10105 ;
  assign n10127 = n30535 & n10126 ;
  assign n10595 = n10109 | n10127 ;
  assign n10596 = n30540 & n9562 ;
  assign n10597 = n10595 | n10596 ;
  assign n10598 = x2 & n10597 ;
  assign n10599 = n733 | n5870 ;
  assign n10600 = x2 & n10599 ;
  assign n10601 = n10597 | n10600 ;
  assign n31939 = ~n10598 ;
  assign n10602 = n31939 & n10601 ;
  assign n10604 = n10594 & n10602 ;
  assign n10603 = n10594 | n10602 ;
  assign n31940 = ~n9631 ;
  assign n10095 = n31940 & n10094 ;
  assign n31941 = ~n10094 ;
  assign n10605 = n9631 & n31941 ;
  assign n10606 = n10095 | n10605 ;
  assign n31942 = ~n10606 ;
  assign n10607 = n10603 & n31942 ;
  assign n10608 = n10604 | n10607 ;
  assign n10609 = n6445 & n9562 ;
  assign n10610 = n30545 & n10126 ;
  assign n10611 = n10609 | n10610 ;
  assign n10612 = x2 & n10611 ;
  assign n10613 = n733 | n5912 ;
  assign n10614 = x2 & n10613 ;
  assign n10615 = n10611 | n10614 ;
  assign n31943 = ~n10612 ;
  assign n10616 = n31943 & n10615 ;
  assign n10618 = n10608 & n10616 ;
  assign n10098 = n9619 & n10097 ;
  assign n10619 = n9619 | n10097 ;
  assign n31944 = ~n10098 ;
  assign n10620 = n31944 & n10619 ;
  assign n10621 = n10608 | n10616 ;
  assign n10622 = n10620 & n10621 ;
  assign n10623 = n10618 | n10622 ;
  assign n10101 = n9608 & n10100 ;
  assign n31945 = ~n10101 ;
  assign n10624 = n31945 & n10102 ;
  assign n31946 = ~n10623 ;
  assign n10626 = n31946 & n10624 ;
  assign n31947 = ~n10626 ;
  assign n10627 = n10102 & n31947 ;
  assign n31948 = ~n10627 ;
  assign n10629 = n9606 & n31948 ;
  assign n31949 = ~n10629 ;
  assign n10630 = n9604 & n31949 ;
  assign n31950 = ~n10630 ;
  assign n10631 = n9549 & n31950 ;
  assign n31951 = ~n10631 ;
  assign n10632 = n9547 & n31951 ;
  assign n10634 = n9047 | n10632 ;
  assign n31952 = ~n9046 ;
  assign n10635 = n31952 & n10634 ;
  assign n31953 = ~n10635 ;
  assign n10636 = n8614 & n31953 ;
  assign n31954 = ~n10636 ;
  assign n10637 = n8612 & n31954 ;
  assign n10640 = n8151 | n10637 ;
  assign n31955 = ~n8149 ;
  assign n10641 = n31955 & n10640 ;
  assign n31956 = ~n10641 ;
  assign n10642 = n7767 & n31956 ;
  assign n31957 = ~n10642 ;
  assign n10643 = n7766 & n31957 ;
  assign n31958 = ~n10643 ;
  assign n10646 = n7416 & n31958 ;
  assign n31959 = ~n10646 ;
  assign n10647 = n7414 & n31959 ;
  assign n31960 = ~n10647 ;
  assign n10649 = n7012 & n31960 ;
  assign n31961 = ~n10649 ;
  assign n10650 = n7010 & n31961 ;
  assign n31962 = ~n10650 ;
  assign n10652 = n6722 & n31962 ;
  assign n31963 = ~n10652 ;
  assign n10653 = n6720 & n31963 ;
  assign n10654 = n6440 & n10653 ;
  assign n10655 = n6440 | n10653 ;
  assign n31964 = ~n10654 ;
  assign n10656 = n31964 & n10655 ;
  assign n10651 = n6722 & n10650 ;
  assign n10678 = n6722 | n10650 ;
  assign n31965 = ~n10651 ;
  assign n10679 = n31965 & n10678 ;
  assign n10648 = n7012 | n10647 ;
  assign n10680 = n7012 & n10647 ;
  assign n31966 = ~n10680 ;
  assign n10681 = n10648 & n31966 ;
  assign n10644 = n7416 & n10643 ;
  assign n10702 = n7416 | n10643 ;
  assign n31967 = ~n10644 ;
  assign n10703 = n31967 & n10702 ;
  assign n31968 = ~n7767 ;
  assign n10726 = n31968 & n10641 ;
  assign n10727 = n10642 | n10726 ;
  assign n31969 = ~n8151 ;
  assign n10638 = n31969 & n10637 ;
  assign n31970 = ~n10637 ;
  assign n10749 = n8151 & n31970 ;
  assign n10750 = n10638 | n10749 ;
  assign n10771 = n8614 & n10635 ;
  assign n10772 = n8614 | n10635 ;
  assign n31971 = ~n10771 ;
  assign n10773 = n31971 & n10772 ;
  assign n31972 = ~n9047 ;
  assign n10633 = n31972 & n10632 ;
  assign n31973 = ~n10632 ;
  assign n10794 = n9047 & n31973 ;
  assign n10795 = n10633 | n10794 ;
  assign n31974 = ~n9549 ;
  assign n10817 = n31974 & n10630 ;
  assign n10818 = n10631 | n10817 ;
  assign n31975 = ~n9606 ;
  assign n10628 = n31975 & n10627 ;
  assign n10841 = n10628 | n10629 ;
  assign n10625 = n10623 & n10624 ;
  assign n10864 = n10623 | n10624 ;
  assign n31976 = ~n10625 ;
  assign n10865 = n31976 & n10864 ;
  assign n31977 = ~n10616 ;
  assign n10617 = n10608 & n31977 ;
  assign n31978 = ~n10608 ;
  assign n10888 = n31978 & n10616 ;
  assign n10889 = n10617 | n10888 ;
  assign n31979 = ~n10620 ;
  assign n10890 = n31979 & n10889 ;
  assign n31980 = ~n10889 ;
  assign n10891 = n10620 & n31980 ;
  assign n10892 = n10890 | n10891 ;
  assign n31981 = ~n10604 ;
  assign n10914 = n10603 & n31981 ;
  assign n10915 = n10606 & n10914 ;
  assign n10916 = n10606 | n10914 ;
  assign n31982 = ~n10915 ;
  assign n10917 = n31982 & n10916 ;
  assign n10939 = n10590 | n10592 ;
  assign n31983 = ~n10593 ;
  assign n10940 = n31983 & n10939 ;
  assign n10973 = n10577 & n10578 ;
  assign n31984 = ~n10973 ;
  assign n10974 = n10579 & n31984 ;
  assign n10989 = n31932 & n10573 ;
  assign n31985 = ~n10575 ;
  assign n10990 = n31985 & n10989 ;
  assign n31986 = ~n10989 ;
  assign n10991 = n10575 & n31986 ;
  assign n10992 = n10990 | n10991 ;
  assign n10994 = n10974 | n10992 ;
  assign n31987 = ~n10940 ;
  assign n10996 = n31987 & n10994 ;
  assign n10998 = n10917 | n10996 ;
  assign n31988 = ~n10892 ;
  assign n10999 = n31988 & n10998 ;
  assign n31989 = ~n10999 ;
  assign n11001 = n10865 & n31989 ;
  assign n11002 = n10841 | n11001 ;
  assign n11004 = n10818 & n11002 ;
  assign n31990 = ~n11004 ;
  assign n11005 = n10795 & n31990 ;
  assign n31991 = ~n11005 ;
  assign n11007 = n10773 & n31991 ;
  assign n31992 = ~n11007 ;
  assign n11008 = n10750 & n31992 ;
  assign n31993 = ~n11008 ;
  assign n11010 = n10727 & n31993 ;
  assign n11011 = n10703 | n11010 ;
  assign n11013 = n10681 & n11011 ;
  assign n31994 = ~n10679 ;
  assign n11014 = n31994 & n11013 ;
  assign n31995 = ~n10974 ;
  assign n10975 = n10940 & n31995 ;
  assign n31996 = ~n10975 ;
  assign n11015 = n10917 & n31996 ;
  assign n31997 = ~n11015 ;
  assign n11016 = n10892 & n31997 ;
  assign n11017 = n10865 | n11016 ;
  assign n11018 = n10841 & n11017 ;
  assign n11019 = n10818 | n11018 ;
  assign n31998 = ~n10795 ;
  assign n11020 = n31998 & n11019 ;
  assign n11021 = n10773 | n11020 ;
  assign n31999 = ~n10750 ;
  assign n11022 = n31999 & n11021 ;
  assign n11023 = n10727 | n11022 ;
  assign n11024 = n10703 & n11023 ;
  assign n11025 = n10681 | n11024 ;
  assign n32000 = ~n11025 ;
  assign n11026 = n10679 & n32000 ;
  assign n11027 = n11014 | n11026 ;
  assign n11028 = n10656 & n11027 ;
  assign n11029 = n10656 | n11027 ;
  assign n32001 = ~n11028 ;
  assign n11030 = n32001 & n11029 ;
  assign n11031 = n889 & n11030 ;
  assign n10689 = n3311 & n10681 ;
  assign n11055 = n3329 & n10679 ;
  assign n11063 = n10689 | n11055 ;
  assign n11064 = n3343 & n10656 ;
  assign n11065 = n11063 | n11064 ;
  assign n11066 = n11031 | n11065 ;
  assign n11068 = n888 & n11066 ;
  assign n32002 = ~n11068 ;
  assign n11069 = n887 & n32002 ;
  assign n731 = n581 & n730 ;
  assign n32003 = ~n731 ;
  assign n11070 = n32003 & n732 ;
  assign n32004 = ~n11069 ;
  assign n11071 = n32004 & n11070 ;
  assign n32005 = ~n11071 ;
  assign n11072 = n732 & n32005 ;
  assign n11073 = n584 & n11072 ;
  assign n11074 = n584 | n11072 ;
  assign n32006 = ~n11073 ;
  assign n11075 = n32006 & n11074 ;
  assign n6167 = n37300 & n30587 ;
  assign n5178 = n30415 & n5166 ;
  assign n5915 = n5191 & n30535 ;
  assign n11076 = n5178 | n5915 ;
  assign n11077 = n5144 & n30530 ;
  assign n11078 = n11076 | n11077 ;
  assign n11079 = n6167 | n11078 ;
  assign n32007 = ~n11079 ;
  assign n11080 = x17 & n32007 ;
  assign n11081 = n30580 & n11079 ;
  assign n11082 = n11080 | n11081 ;
  assign n5747 = n4686 & n30512 ;
  assign n4819 = n4726 & n4811 ;
  assign n5109 = n4706 & n30405 ;
  assign n11083 = n4819 | n5109 ;
  assign n11084 = n4748 & n5017 ;
  assign n11085 = n11083 | n11084 ;
  assign n11086 = n5747 | n11085 ;
  assign n32008 = ~n11086 ;
  assign n11087 = x20 & n32008 ;
  assign n11088 = n30374 & n11086 ;
  assign n11089 = n11087 | n11088 ;
  assign n4445 = n3791 & n4442 ;
  assign n3865 = n209 & n30264 ;
  assign n4095 = n3802 & n4093 ;
  assign n11090 = n3865 | n4095 ;
  assign n11091 = n3818 & n4033 ;
  assign n11092 = n11090 | n11091 ;
  assign n11093 = n4445 | n11092 ;
  assign n11094 = x26 | n11093 ;
  assign n11095 = x26 & n11093 ;
  assign n32009 = ~n11095 ;
  assign n11096 = n11094 & n32009 ;
  assign n11097 = n3367 | n3379 ;
  assign n11098 = n2983 | n3048 ;
  assign n11099 = n492 | n532 ;
  assign n11100 = n662 | n1455 ;
  assign n11101 = n11099 | n11100 ;
  assign n11102 = n759 | n11101 ;
  assign n11103 = n2704 | n11102 ;
  assign n11104 = n282 | n300 ;
  assign n11105 = n670 | n11104 ;
  assign n11106 = n1879 | n11105 ;
  assign n11107 = n2397 | n2917 ;
  assign n11108 = n11106 | n11107 ;
  assign n11109 = n807 | n1200 ;
  assign n11110 = n4526 | n4538 ;
  assign n11111 = n11109 | n11110 ;
  assign n11112 = n5292 | n11111 ;
  assign n11113 = n11108 | n11112 ;
  assign n11114 = n4306 | n11113 ;
  assign n11115 = n11103 | n11114 ;
  assign n11116 = n163 | n253 ;
  assign n11117 = n428 | n11116 ;
  assign n11118 = n621 | n11117 ;
  assign n11119 = n349 | n441 ;
  assign n11120 = n509 | n11119 ;
  assign n11121 = n2500 | n11120 ;
  assign n11122 = n11118 | n11121 ;
  assign n11123 = n2409 | n11122 ;
  assign n11124 = n296 | n1895 ;
  assign n11125 = n3737 | n11124 ;
  assign n11126 = n293 | n647 ;
  assign n11127 = n568 | n11126 ;
  assign n11128 = n721 | n811 ;
  assign n11129 = n1111 | n11128 ;
  assign n11130 = n11127 | n11129 ;
  assign n11131 = n11125 | n11130 ;
  assign n11132 = n4655 | n11131 ;
  assign n11133 = n11123 | n11132 ;
  assign n11134 = n925 | n1091 ;
  assign n11135 = n553 | n698 ;
  assign n11136 = n11134 | n11135 ;
  assign n11137 = n162 | n332 ;
  assign n11138 = n469 | n520 ;
  assign n11139 = n11137 | n11138 ;
  assign n11140 = n104 | n411 ;
  assign n11141 = n11139 | n11140 ;
  assign n11142 = n3272 | n3683 ;
  assign n11143 = n11141 | n11142 ;
  assign n11144 = n11136 | n11143 ;
  assign n11145 = n793 | n2225 ;
  assign n11146 = n451 | n635 ;
  assign n11147 = n2477 | n11146 ;
  assign n11148 = n4791 | n4986 ;
  assign n11149 = n11147 | n11148 ;
  assign n11150 = n420 | n916 ;
  assign n11151 = n11149 | n11150 ;
  assign n11152 = n11145 | n11151 ;
  assign n11153 = n257 | n338 ;
  assign n11154 = n345 | n11153 ;
  assign n11155 = n4020 | n4274 ;
  assign n11156 = n11154 | n11155 ;
  assign n11157 = n3004 | n11156 ;
  assign n11158 = n11152 | n11157 ;
  assign n11159 = n11144 | n11158 ;
  assign n11160 = n11133 | n11159 ;
  assign n11161 = n11115 | n11160 ;
  assign n32010 = ~n11161 ;
  assign n11162 = n11098 & n32010 ;
  assign n32011 = ~n11098 ;
  assign n11163 = n32011 & n11161 ;
  assign n11164 = n11162 | n11163 ;
  assign n3630 = n889 & n30238 ;
  assign n3320 = n1445 & n3311 ;
  assign n3342 = n30082 & n3329 ;
  assign n11165 = n3320 | n3342 ;
  assign n11166 = n1219 & n3343 ;
  assign n11167 = n11165 | n11166 ;
  assign n11168 = n3630 | n11167 ;
  assign n11169 = n11164 | n11168 ;
  assign n11171 = n11164 & n11168 ;
  assign n32012 = ~n11171 ;
  assign n11172 = n11169 & n32012 ;
  assign n11173 = n11097 & n11172 ;
  assign n4422 = n895 & n4420 ;
  assign n2853 = n1074 & n2849 ;
  assign n3770 = n894 & n3764 ;
  assign n11174 = n2853 | n3770 ;
  assign n11175 = n30074 & n2861 ;
  assign n11176 = n11174 | n11175 ;
  assign n11177 = n4422 | n11176 ;
  assign n32013 = ~n11177 ;
  assign n11178 = x29 & n32013 ;
  assign n11179 = n30024 & n11177 ;
  assign n11180 = n11178 | n11179 ;
  assign n11181 = n11097 | n11172 ;
  assign n32014 = ~n11173 ;
  assign n11182 = n32014 & n11181 ;
  assign n32015 = ~n11180 ;
  assign n11183 = n32015 & n11182 ;
  assign n11184 = n11173 | n11183 ;
  assign n11185 = n253 | n312 ;
  assign n11186 = n451 | n512 ;
  assign n11187 = n608 | n11186 ;
  assign n11188 = n11185 | n11187 ;
  assign n11189 = n320 | n432 ;
  assign n11190 = n479 | n11189 ;
  assign n11191 = n276 | n713 ;
  assign n11192 = n756 | n11191 ;
  assign n11193 = n11190 | n11192 ;
  assign n11194 = n2457 | n4635 ;
  assign n11195 = n11193 | n11194 ;
  assign n11196 = n11188 | n11195 ;
  assign n11197 = n359 | n369 ;
  assign n11198 = n195 | n11197 ;
  assign n11199 = n488 | n2768 ;
  assign n11200 = n11198 | n11199 ;
  assign n11201 = n1855 | n11200 ;
  assign n11202 = n4295 | n11201 ;
  assign n11203 = n202 | n410 ;
  assign n11204 = n554 | n679 ;
  assign n11205 = n11203 | n11204 ;
  assign n11206 = n2887 | n11205 ;
  assign n11207 = n1130 | n11206 ;
  assign n11208 = n199 | n750 ;
  assign n11209 = n653 | n4911 ;
  assign n11210 = n11208 | n11209 ;
  assign n11211 = n11207 | n11210 ;
  assign n11212 = n11202 | n11211 ;
  assign n11213 = n11196 | n11212 ;
  assign n11214 = n5000 | n5830 ;
  assign n11215 = n434 | n446 ;
  assign n11216 = n956 | n11215 ;
  assign n11217 = n1892 | n4255 ;
  assign n11218 = n11216 | n11217 ;
  assign n11219 = n834 | n2147 ;
  assign n11220 = n11218 | n11219 ;
  assign n11221 = n11214 | n11220 ;
  assign n11222 = n179 | n314 ;
  assign n11223 = n233 | n2071 ;
  assign n11224 = n11222 | n11223 ;
  assign n11225 = n168 | n1787 ;
  assign n11226 = n788 | n11225 ;
  assign n11227 = n97 | n239 ;
  assign n11228 = n11226 | n11227 ;
  assign n11229 = n11224 | n11228 ;
  assign n11230 = n366 | n469 ;
  assign n11231 = n4978 | n11230 ;
  assign n11232 = n405 | n491 ;
  assign n11233 = n3125 | n11232 ;
  assign n11234 = n570 | n780 ;
  assign n11235 = n11233 | n11234 ;
  assign n11236 = n11231 | n11235 ;
  assign n11237 = n11229 | n11236 ;
  assign n11238 = n11221 | n11237 ;
  assign n11239 = n4340 | n4597 ;
  assign n11240 = n532 | n815 ;
  assign n11241 = n2732 | n11240 ;
  assign n11242 = n3900 | n11241 ;
  assign n11243 = n11239 | n11242 ;
  assign n11244 = n595 | n2394 ;
  assign n11245 = n3753 | n11244 ;
  assign n11246 = n162 | n241 ;
  assign n11247 = n2243 | n3233 ;
  assign n11248 = n11246 | n11247 ;
  assign n11249 = n346 | n368 ;
  assign n11250 = n642 | n11249 ;
  assign n11251 = n849 | n1323 ;
  assign n11252 = n11250 | n11251 ;
  assign n11253 = n11248 | n11252 ;
  assign n11254 = n11245 | n11253 ;
  assign n11255 = n11243 | n11254 ;
  assign n11256 = n11238 | n11255 ;
  assign n11257 = n11213 | n11256 ;
  assign n11258 = n32010 & n11257 ;
  assign n32016 = ~n11257 ;
  assign n11259 = n11161 & n32016 ;
  assign n11260 = n11258 | n11259 ;
  assign n3399 = n889 & n30212 ;
  assign n3313 = n30082 & n3311 ;
  assign n3352 = n30074 & n3343 ;
  assign n11261 = n3313 | n3352 ;
  assign n11262 = n1219 & n3329 ;
  assign n11263 = n11261 | n11262 ;
  assign n11264 = n3399 | n11263 ;
  assign n11265 = n11260 | n11264 ;
  assign n11267 = n11260 & n11264 ;
  assign n32017 = ~n11267 ;
  assign n11268 = n11265 & n32017 ;
  assign n11170 = n11162 | n11168 ;
  assign n32018 = ~n11163 ;
  assign n11269 = n32018 & n11170 ;
  assign n11270 = n11268 & n11269 ;
  assign n11271 = n11268 | n11269 ;
  assign n32019 = ~n11270 ;
  assign n11272 = n32019 & n11271 ;
  assign n32020 = ~n11272 ;
  assign n11273 = n11184 & n32020 ;
  assign n32021 = ~n11184 ;
  assign n11274 = n32021 & n11272 ;
  assign n11275 = n11273 | n11274 ;
  assign n3789 = n895 & n3787 ;
  assign n2874 = n1074 & n2861 ;
  assign n3766 = n2849 & n3764 ;
  assign n11276 = n2874 | n3766 ;
  assign n11277 = n894 & n3700 ;
  assign n11278 = n11276 | n11277 ;
  assign n11279 = n3789 | n11278 ;
  assign n32022 = ~n11279 ;
  assign n11280 = x29 & n32022 ;
  assign n11281 = n30024 & n11279 ;
  assign n11282 = n11280 | n11281 ;
  assign n11283 = n11275 | n11282 ;
  assign n11284 = n11275 & n11282 ;
  assign n32023 = ~n11284 ;
  assign n11285 = n11283 & n32023 ;
  assign n11286 = n11096 & n11285 ;
  assign n11287 = n11096 | n11285 ;
  assign n32024 = ~n11286 ;
  assign n11288 = n32024 & n11287 ;
  assign n32025 = ~n11182 ;
  assign n11289 = n11180 & n32025 ;
  assign n11290 = n11183 | n11289 ;
  assign n11291 = n3381 | n3410 ;
  assign n32026 = ~n3414 ;
  assign n11292 = n32026 & n11291 ;
  assign n11294 = n11290 & n11292 ;
  assign n4509 = n3791 & n30349 ;
  assign n3706 = n209 & n3700 ;
  assign n4094 = n3818 & n4093 ;
  assign n11295 = n3706 | n4094 ;
  assign n11296 = n3802 & n30264 ;
  assign n11297 = n11295 | n11296 ;
  assign n11298 = n4509 | n11297 ;
  assign n32027 = ~n11298 ;
  assign n11299 = x26 & n32027 ;
  assign n11300 = n30019 & n11298 ;
  assign n11301 = n11299 | n11300 ;
  assign n32028 = ~n11290 ;
  assign n11293 = n32028 & n11292 ;
  assign n32029 = ~n11292 ;
  assign n11302 = n11290 & n32029 ;
  assign n11303 = n11293 | n11302 ;
  assign n11305 = n11301 & n11303 ;
  assign n11306 = n11294 | n11305 ;
  assign n32030 = ~n11306 ;
  assign n11307 = n11288 & n32030 ;
  assign n32031 = ~n11288 ;
  assign n11308 = n32031 & n11306 ;
  assign n11309 = n11307 | n11308 ;
  assign n4676 = n4135 & n4674 ;
  assign n4575 = n4148 & n30361 ;
  assign n4667 = n4165 & n4664 ;
  assign n11310 = n4575 | n4667 ;
  assign n11311 = n30282 & n4185 ;
  assign n11312 = n11310 | n11311 ;
  assign n11313 = n4676 | n11312 ;
  assign n32032 = ~n11313 ;
  assign n11314 = x23 & n32032 ;
  assign n11315 = n30030 & n11313 ;
  assign n11316 = n11314 | n11315 ;
  assign n32033 = ~n11316 ;
  assign n11317 = n11309 & n32033 ;
  assign n32034 = ~n11309 ;
  assign n11318 = n32034 & n11316 ;
  assign n11319 = n11317 | n11318 ;
  assign n32035 = ~n11301 ;
  assign n11304 = n32035 & n11303 ;
  assign n32036 = ~n11303 ;
  assign n11320 = n11301 & n32036 ;
  assign n11321 = n11304 | n11320 ;
  assign n32037 = ~n3884 ;
  assign n11322 = n3846 & n32037 ;
  assign n11324 = n11321 | n11322 ;
  assign n32038 = ~n11321 ;
  assign n11323 = n32038 & n11322 ;
  assign n32039 = ~n11322 ;
  assign n11325 = n11321 & n32039 ;
  assign n11326 = n11323 | n11325 ;
  assign n5727 = n4135 & n5723 ;
  assign n4195 = n4033 & n4185 ;
  assign n4571 = n4165 & n30361 ;
  assign n11327 = n4195 | n4571 ;
  assign n11328 = n30282 & n4148 ;
  assign n11329 = n11327 | n11328 ;
  assign n11330 = n5727 | n11329 ;
  assign n32040 = ~n11330 ;
  assign n11331 = x23 & n32040 ;
  assign n11332 = n30030 & n11330 ;
  assign n11333 = n11331 | n11332 ;
  assign n32041 = ~n11333 ;
  assign n11334 = n11326 & n32041 ;
  assign n32042 = ~n11334 ;
  assign n11335 = n11324 & n32042 ;
  assign n32043 = ~n11319 ;
  assign n11336 = n32043 & n11335 ;
  assign n32044 = ~n11335 ;
  assign n11337 = n11319 & n32044 ;
  assign n11338 = n11336 | n11337 ;
  assign n32045 = ~n11089 ;
  assign n11339 = n32045 & n11338 ;
  assign n32046 = ~n11338 ;
  assign n11340 = n11089 & n32046 ;
  assign n11341 = n11339 | n11340 ;
  assign n32047 = ~n11326 ;
  assign n11342 = n32047 & n11333 ;
  assign n11343 = n11334 | n11342 ;
  assign n11344 = n3886 | n4210 ;
  assign n32048 = ~n4457 ;
  assign n11345 = n4213 & n32048 ;
  assign n32049 = ~n11345 ;
  assign n11346 = n11344 & n32049 ;
  assign n11348 = n11343 | n11346 ;
  assign n6144 = n4686 & n30578 ;
  assign n4743 = n4664 & n4726 ;
  assign n4817 = n4706 & n4811 ;
  assign n11349 = n4743 | n4817 ;
  assign n11350 = n4748 & n30405 ;
  assign n11351 = n11349 | n11350 ;
  assign n11352 = n6144 | n11351 ;
  assign n32050 = ~n11352 ;
  assign n11353 = x20 & n32050 ;
  assign n11354 = n30374 & n11352 ;
  assign n11355 = n11353 | n11354 ;
  assign n32051 = ~n11343 ;
  assign n11347 = n32051 & n11346 ;
  assign n32052 = ~n11346 ;
  assign n11356 = n11343 & n32052 ;
  assign n11357 = n11347 | n11356 ;
  assign n32053 = ~n11355 ;
  assign n11358 = n32053 & n11357 ;
  assign n32054 = ~n11358 ;
  assign n11359 = n11348 & n32054 ;
  assign n32055 = ~n11341 ;
  assign n11360 = n32055 & n11359 ;
  assign n32056 = ~n11359 ;
  assign n11361 = n11341 & n32056 ;
  assign n11362 = n11360 | n11361 ;
  assign n32057 = ~n11082 ;
  assign n11363 = n32057 & n11362 ;
  assign n32058 = ~n11362 ;
  assign n11364 = n11082 & n32058 ;
  assign n11365 = n11363 | n11364 ;
  assign n6268 = n5937 & n30597 ;
  assign n11366 = n5994 | n6268 ;
  assign n11367 = n30545 & n11366 ;
  assign n11368 = x14 & n11367 ;
  assign n11369 = x14 | n11367 ;
  assign n32059 = ~n11368 ;
  assign n11370 = n32059 & n11369 ;
  assign n32060 = ~n11357 ;
  assign n11371 = n11355 & n32060 ;
  assign n11372 = n11358 | n11371 ;
  assign n11373 = n4460 | n4777 ;
  assign n32061 = ~n4851 ;
  assign n11374 = n32061 & n11373 ;
  assign n11376 = n11372 | n11374 ;
  assign n6415 = n37300 & n6411 ;
  assign n5162 = n30415 & n5144 ;
  assign n5168 = n5017 & n5166 ;
  assign n11377 = n5162 | n5168 ;
  assign n11378 = n5191 & n30530 ;
  assign n11379 = n11377 | n11378 ;
  assign n11380 = n6415 | n11379 ;
  assign n32062 = ~n11380 ;
  assign n11381 = x17 & n32062 ;
  assign n11382 = n30580 & n11380 ;
  assign n11383 = n11381 | n11382 ;
  assign n32063 = ~n11372 ;
  assign n11375 = n32063 & n11374 ;
  assign n32064 = ~n11374 ;
  assign n11384 = n11372 & n32064 ;
  assign n11385 = n11375 | n11384 ;
  assign n32065 = ~n11383 ;
  assign n11386 = n32065 & n11385 ;
  assign n32066 = ~n11386 ;
  assign n11387 = n11376 & n32066 ;
  assign n11388 = n11370 & n11387 ;
  assign n11389 = n11370 | n11387 ;
  assign n32067 = ~n11388 ;
  assign n11390 = n32067 & n11389 ;
  assign n32068 = ~n11365 ;
  assign n11391 = n32068 & n11390 ;
  assign n32069 = ~n11390 ;
  assign n11392 = n11365 & n32069 ;
  assign n11393 = n11391 | n11392 ;
  assign n6448 = n5937 & n6445 ;
  assign n11394 = n30545 & n5970 ;
  assign n11395 = n30535 & n5994 ;
  assign n11396 = n11394 | n11395 ;
  assign n11397 = n6448 | n11396 ;
  assign n11398 = x14 | n11397 ;
  assign n11399 = x14 & n11397 ;
  assign n32070 = ~n11399 ;
  assign n11400 = n11398 & n32070 ;
  assign n11401 = n4853 | n5219 ;
  assign n32071 = ~n5760 ;
  assign n11402 = n5222 & n32071 ;
  assign n32072 = ~n11402 ;
  assign n11403 = n11401 & n32072 ;
  assign n11404 = n11400 & n11403 ;
  assign n32073 = ~n11385 ;
  assign n11405 = n11383 & n32073 ;
  assign n11406 = n11386 | n11405 ;
  assign n11407 = n11400 | n11403 ;
  assign n32074 = ~n11404 ;
  assign n11408 = n32074 & n11407 ;
  assign n11410 = n11406 & n11408 ;
  assign n11411 = n11404 | n11410 ;
  assign n32075 = ~n11411 ;
  assign n11412 = n11393 & n32075 ;
  assign n32076 = ~n11393 ;
  assign n11413 = n32076 & n11411 ;
  assign n11414 = n11412 | n11413 ;
  assign n32077 = ~n11406 ;
  assign n11409 = n32077 & n11408 ;
  assign n32078 = ~n11408 ;
  assign n11415 = n11406 & n32078 ;
  assign n11416 = n11409 | n11415 ;
  assign n32079 = ~n6182 ;
  assign n11417 = n6050 & n32079 ;
  assign n11419 = n11416 | n11417 ;
  assign n11418 = n11416 & n11417 ;
  assign n32080 = ~n11418 ;
  assign n11420 = n32080 & n11419 ;
  assign n11421 = n6184 | n6437 ;
  assign n32081 = ~n10653 ;
  assign n11422 = n6440 & n32081 ;
  assign n32082 = ~n11422 ;
  assign n11423 = n11421 & n32082 ;
  assign n32083 = ~n11423 ;
  assign n11426 = n11420 & n32083 ;
  assign n32084 = ~n11426 ;
  assign n11427 = n11419 & n32084 ;
  assign n32085 = ~n11427 ;
  assign n11428 = n11414 & n32085 ;
  assign n32086 = ~n11414 ;
  assign n11429 = n32086 & n11427 ;
  assign n11430 = n11428 | n11429 ;
  assign n32087 = ~n11420 ;
  assign n11424 = n32087 & n11423 ;
  assign n11452 = n11424 | n11426 ;
  assign n11453 = n10679 | n11013 ;
  assign n11455 = n10656 & n11453 ;
  assign n32088 = ~n11452 ;
  assign n11456 = n32088 & n11455 ;
  assign n11457 = n10679 & n11025 ;
  assign n11458 = n10656 | n11457 ;
  assign n32089 = ~n11458 ;
  assign n11459 = n11452 & n32089 ;
  assign n11460 = n11456 | n11459 ;
  assign n11461 = n11430 & n11460 ;
  assign n11462 = n11430 | n11460 ;
  assign n32090 = ~n11461 ;
  assign n11463 = n32090 & n11462 ;
  assign n11466 = n889 & n11463 ;
  assign n10667 = n3311 & n10656 ;
  assign n11425 = n11420 & n11423 ;
  assign n11475 = n11420 | n11423 ;
  assign n32091 = ~n11425 ;
  assign n11476 = n32091 & n11475 ;
  assign n11483 = n3329 & n11476 ;
  assign n11498 = n10667 | n11483 ;
  assign n11499 = n3343 & n11430 ;
  assign n11500 = n11498 | n11499 ;
  assign n11501 = n11466 | n11500 ;
  assign n11502 = n11075 | n11501 ;
  assign n11503 = n11075 & n11501 ;
  assign n32092 = ~n11503 ;
  assign n11504 = n11502 & n32092 ;
  assign n32093 = ~n11070 ;
  assign n11505 = n11069 & n32093 ;
  assign n11506 = n11071 | n11505 ;
  assign n32094 = ~n11453 ;
  assign n11454 = n10656 & n32094 ;
  assign n32095 = ~n10656 ;
  assign n11507 = n32095 & n11457 ;
  assign n11508 = n11454 | n11507 ;
  assign n11509 = n11476 & n11508 ;
  assign n11510 = n11476 | n11508 ;
  assign n32096 = ~n11509 ;
  assign n11511 = n32096 & n11510 ;
  assign n11512 = n889 & n11511 ;
  assign n10665 = n3329 & n10656 ;
  assign n11052 = n3311 & n10679 ;
  assign n11523 = n10665 | n11052 ;
  assign n11524 = n3343 & n11452 ;
  assign n11525 = n11523 | n11524 ;
  assign n11526 = n11512 | n11525 ;
  assign n32097 = ~n11526 ;
  assign n11528 = n11506 & n32097 ;
  assign n11067 = n888 | n11066 ;
  assign n11529 = n11067 & n32002 ;
  assign n32098 = ~n745 ;
  assign n746 = n744 & n32098 ;
  assign n883 = n746 & n882 ;
  assign n11530 = n746 | n882 ;
  assign n32099 = ~n883 ;
  assign n11531 = n32099 & n11530 ;
  assign n32100 = ~n11011 ;
  assign n11012 = n10681 & n32100 ;
  assign n32101 = ~n10681 ;
  assign n11532 = n32101 & n11024 ;
  assign n11533 = n11012 | n11532 ;
  assign n11534 = n10679 & n11533 ;
  assign n11535 = n10679 | n11533 ;
  assign n32102 = ~n11534 ;
  assign n11536 = n32102 & n11535 ;
  assign n11537 = n889 & n11536 ;
  assign n10690 = n3329 & n10681 ;
  assign n10709 = n3311 & n10703 ;
  assign n11548 = n10690 | n10709 ;
  assign n11549 = n3343 & n10679 ;
  assign n11550 = n11548 | n11549 ;
  assign n11551 = n11537 | n11550 ;
  assign n32103 = ~n11551 ;
  assign n11552 = n11531 & n32103 ;
  assign n11553 = n130 | n310 ;
  assign n11554 = n4967 | n11553 ;
  assign n11555 = n11134 | n11554 ;
  assign n11556 = n335 | n594 ;
  assign n11557 = n448 | n668 ;
  assign n11558 = n765 | n11557 ;
  assign n11559 = n11556 | n11558 ;
  assign n11560 = n11555 | n11559 ;
  assign n11561 = n2627 | n11560 ;
  assign n11562 = n190 | n331 ;
  assign n11563 = n666 | n11562 ;
  assign n11564 = n3001 | n11563 ;
  assign n11565 = n345 | n349 ;
  assign n11566 = n845 | n11565 ;
  assign n11567 = n4636 | n11566 ;
  assign n11568 = n11564 | n11567 ;
  assign n11569 = n3080 | n11568 ;
  assign n11570 = n11561 | n11569 ;
  assign n11571 = n2950 | n11570 ;
  assign n11572 = n201 | n478 ;
  assign n11573 = n923 | n2514 ;
  assign n11574 = n11572 | n11573 ;
  assign n11575 = n240 | n332 ;
  assign n11576 = n440 | n446 ;
  assign n11577 = n2229 | n11576 ;
  assign n11578 = n11575 | n11577 ;
  assign n11579 = n167 | n269 ;
  assign n11580 = n377 | n528 ;
  assign n11581 = n11579 | n11580 ;
  assign n32104 = ~n11581 ;
  assign n11582 = n835 & n32104 ;
  assign n32105 = ~n11578 ;
  assign n11583 = n32105 & n11582 ;
  assign n32106 = ~n3527 ;
  assign n11584 = n32106 & n11583 ;
  assign n32107 = ~n11574 ;
  assign n11585 = n32107 & n11584 ;
  assign n32108 = ~n4946 ;
  assign n11586 = n32108 & n11585 ;
  assign n32109 = ~n11571 ;
  assign n11587 = n32109 & n11586 ;
  assign n32110 = ~n734 ;
  assign n11589 = n32110 & n11587 ;
  assign n11588 = n734 & n11587 ;
  assign n11590 = n734 | n11587 ;
  assign n32111 = ~n11588 ;
  assign n11591 = n32111 & n11590 ;
  assign n11592 = n677 | n1865 ;
  assign n11593 = n11246 | n11592 ;
  assign n11594 = n319 | n399 ;
  assign n11595 = n684 | n11594 ;
  assign n11596 = n257 | n280 ;
  assign n11597 = n237 | n11596 ;
  assign n11598 = n11595 | n11597 ;
  assign n11599 = n11593 | n11598 ;
  assign n11600 = n282 | n529 ;
  assign n11601 = n679 | n2517 ;
  assign n11602 = n11600 | n11601 ;
  assign n11603 = n1847 | n11602 ;
  assign n11604 = n11599 | n11603 ;
  assign n11605 = n1609 | n4052 ;
  assign n11606 = n224 | n453 ;
  assign n11607 = n920 | n11606 ;
  assign n11608 = n5823 | n11607 ;
  assign n11609 = n11605 | n11608 ;
  assign n11610 = n3059 | n11609 ;
  assign n11611 = n4014 | n11610 ;
  assign n11612 = n11604 | n11611 ;
  assign n11613 = n822 | n11612 ;
  assign n11615 = n734 | n11613 ;
  assign n32112 = ~n11613 ;
  assign n11614 = n734 & n32112 ;
  assign n11616 = n32110 & n11613 ;
  assign n11617 = n11614 | n11616 ;
  assign n11618 = n461 | n473 ;
  assign n11619 = n1129 | n11618 ;
  assign n11620 = n1106 | n11619 ;
  assign n11621 = n2200 | n2920 ;
  assign n11622 = n11620 | n11621 ;
  assign n11623 = n348 | n487 ;
  assign n11624 = n1179 | n11623 ;
  assign n11625 = n428 | n11624 ;
  assign n11626 = n2224 | n2767 ;
  assign n11627 = n5354 | n11626 ;
  assign n11628 = n11625 | n11627 ;
  assign n11629 = n11622 | n11628 ;
  assign n11630 = n187 | n368 ;
  assign n11631 = n634 | n11630 ;
  assign n11632 = n900 | n2037 ;
  assign n11633 = n2182 | n11632 ;
  assign n11634 = n11631 | n11633 ;
  assign n11635 = n1657 | n11634 ;
  assign n11636 = n11629 | n11635 ;
  assign n11637 = n440 | n841 ;
  assign n11638 = n1272 | n11637 ;
  assign n11639 = n1593 | n11638 ;
  assign n11640 = n11636 | n11639 ;
  assign n11641 = n401 | n554 ;
  assign n11642 = n687 | n11641 ;
  assign n11643 = n433 | n1091 ;
  assign n11644 = n273 | n354 ;
  assign n11645 = n11643 | n11644 ;
  assign n11646 = n11642 | n11645 ;
  assign n11647 = n983 | n1041 ;
  assign n11648 = n1123 | n2169 ;
  assign n11649 = n11647 | n11648 ;
  assign n11650 = n11646 | n11649 ;
  assign n11651 = n2397 | n3997 ;
  assign n11652 = n5082 | n11651 ;
  assign n11653 = n1877 | n11652 ;
  assign n11654 = n11650 | n11653 ;
  assign n11655 = n223 | n269 ;
  assign n11656 = n360 | n501 ;
  assign n11657 = n11655 | n11656 ;
  assign n11658 = n80 | n434 ;
  assign n11659 = n2051 | n11658 ;
  assign n11660 = n11657 | n11659 ;
  assign n11661 = n1383 | n11660 ;
  assign n11662 = n1647 | n11661 ;
  assign n11663 = n399 | n865 ;
  assign n11664 = n239 | n11663 ;
  assign n11665 = n400 | n814 ;
  assign n11666 = n1606 | n11665 ;
  assign n11667 = n11664 | n11666 ;
  assign n11668 = n5040 | n11667 ;
  assign n32113 = ~n1200 ;
  assign n11669 = n145 & n32113 ;
  assign n11670 = n749 | n4005 ;
  assign n32114 = ~n11670 ;
  assign n11671 = n11669 & n32114 ;
  assign n32115 = ~n11668 ;
  assign n11672 = n32115 & n11671 ;
  assign n32116 = ~n11662 ;
  assign n11673 = n32116 & n11672 ;
  assign n32117 = ~n11654 ;
  assign n11674 = n32117 & n11673 ;
  assign n32118 = ~n11640 ;
  assign n11675 = n32118 & n11674 ;
  assign n32119 = ~n11675 ;
  assign n11677 = n734 & n32119 ;
  assign n11676 = n734 & n11675 ;
  assign n11678 = n734 | n11675 ;
  assign n32120 = ~n11676 ;
  assign n11679 = n32120 & n11678 ;
  assign n10639 = n8151 & n10637 ;
  assign n32121 = ~n10639 ;
  assign n11680 = n32121 & n10640 ;
  assign n11681 = n11007 & n11680 ;
  assign n11682 = n11021 | n11680 ;
  assign n32122 = ~n11681 ;
  assign n11683 = n32122 & n11682 ;
  assign n32123 = ~n11683 ;
  assign n11684 = n10727 & n32123 ;
  assign n32124 = ~n10727 ;
  assign n11685 = n32124 & n11683 ;
  assign n11686 = n11684 | n11685 ;
  assign n32125 = ~n11686 ;
  assign n11687 = n889 & n32125 ;
  assign n10764 = n3329 & n31999 ;
  assign n10785 = n3311 & n10773 ;
  assign n11698 = n10764 | n10785 ;
  assign n11699 = n3343 & n10727 ;
  assign n11700 = n11698 | n11699 ;
  assign n11701 = n11687 | n11700 ;
  assign n32126 = ~n11679 ;
  assign n11703 = n32126 & n11701 ;
  assign n11704 = n11677 | n11703 ;
  assign n32127 = ~n11704 ;
  assign n11705 = n11617 & n32127 ;
  assign n32128 = ~n11705 ;
  assign n11706 = n11615 & n32128 ;
  assign n11708 = n11591 | n11706 ;
  assign n32129 = ~n11589 ;
  assign n11709 = n32129 & n11708 ;
  assign n32130 = ~n11531 ;
  assign n11710 = n32130 & n11551 ;
  assign n11711 = n11552 | n11710 ;
  assign n11712 = n11709 | n11711 ;
  assign n32131 = ~n11552 ;
  assign n11713 = n32131 & n11712 ;
  assign n11715 = n11529 | n11713 ;
  assign n5139 = n4686 & n30410 ;
  assign n4933 = n4748 & n30415 ;
  assign n5112 = n4726 & n30405 ;
  assign n11716 = n4933 | n5112 ;
  assign n11717 = n4706 & n5017 ;
  assign n11718 = n11716 | n11717 ;
  assign n11719 = n5139 | n11718 ;
  assign n32132 = ~n11719 ;
  assign n11720 = x20 & n32132 ;
  assign n11721 = n30374 & n11719 ;
  assign n11722 = n11720 | n11721 ;
  assign n3875 = n895 & n30263 ;
  assign n3708 = n2849 & n3700 ;
  assign n3771 = n2861 & n3764 ;
  assign n11723 = n3708 | n3771 ;
  assign n11724 = n894 & n30264 ;
  assign n11725 = n11723 | n11724 ;
  assign n11726 = n3875 | n11725 ;
  assign n32133 = ~n11726 ;
  assign n11727 = x29 & n32133 ;
  assign n11728 = n30024 & n11726 ;
  assign n11729 = n11727 | n11728 ;
  assign n32134 = ~n112 ;
  assign n11730 = n32134 & n145 ;
  assign n32135 = ~n280 ;
  assign n11731 = n32135 & n11730 ;
  assign n32136 = ~n1466 ;
  assign n11732 = n32136 & n11731 ;
  assign n32137 = ~n2962 ;
  assign n11733 = n32137 & n11732 ;
  assign n11734 = n1731 | n2287 ;
  assign n11735 = n11665 | n11734 ;
  assign n11736 = n951 | n11735 ;
  assign n32138 = ~n11736 ;
  assign n11737 = n11733 & n32138 ;
  assign n11738 = n2458 | n3728 ;
  assign n11739 = n897 | n1210 ;
  assign n11740 = n5060 | n11739 ;
  assign n11741 = n11738 | n11740 ;
  assign n11742 = n797 | n1927 ;
  assign n11743 = n2906 | n11742 ;
  assign n11744 = n296 | n767 ;
  assign n11745 = n237 | n11744 ;
  assign n11746 = n1634 | n11745 ;
  assign n11747 = n11743 | n11746 ;
  assign n11748 = n11741 | n11747 ;
  assign n11749 = n3255 | n11748 ;
  assign n32139 = ~n11749 ;
  assign n11750 = n11737 & n32139 ;
  assign n32140 = ~n5315 ;
  assign n11751 = n32140 & n11750 ;
  assign n32141 = ~n3516 ;
  assign n11752 = n32141 & n11751 ;
  assign n11753 = n32010 & n11752 ;
  assign n32142 = ~n11752 ;
  assign n11754 = n11161 & n32142 ;
  assign n11755 = n11753 | n11754 ;
  assign n11756 = x14 | n11755 ;
  assign n11757 = x14 & n11755 ;
  assign n32143 = ~n11757 ;
  assign n11758 = n11756 & n32143 ;
  assign n11266 = n11258 | n11264 ;
  assign n32144 = ~n11259 ;
  assign n11759 = n32144 & n11266 ;
  assign n11760 = n11758 & n11759 ;
  assign n11761 = n11758 | n11759 ;
  assign n32145 = ~n11760 ;
  assign n11762 = n32145 & n11761 ;
  assign n2848 = n889 & n30173 ;
  assign n3312 = n1219 & n3311 ;
  assign n3356 = n1074 & n3343 ;
  assign n11763 = n3312 | n3356 ;
  assign n11764 = n30074 & n3329 ;
  assign n11765 = n11763 | n11764 ;
  assign n11766 = n2848 | n11765 ;
  assign n32146 = ~n11766 ;
  assign n11767 = n11762 & n32146 ;
  assign n32147 = ~n11762 ;
  assign n11768 = n32147 & n11766 ;
  assign n11769 = n11767 | n11768 ;
  assign n32148 = ~n11269 ;
  assign n11770 = n11268 & n32148 ;
  assign n11771 = n11273 | n11770 ;
  assign n11772 = n11769 | n11771 ;
  assign n11773 = n11769 & n11771 ;
  assign n32149 = ~n11773 ;
  assign n11774 = n11772 & n32149 ;
  assign n11775 = n11729 | n11774 ;
  assign n11776 = n11729 & n11774 ;
  assign n32150 = ~n11776 ;
  assign n11777 = n11775 & n32150 ;
  assign n4127 = n3791 & n30286 ;
  assign n4036 = n3802 & n4033 ;
  assign n4104 = n209 & n4093 ;
  assign n11778 = n4036 | n4104 ;
  assign n11779 = n3818 & n30282 ;
  assign n11780 = n11778 | n11779 ;
  assign n11781 = n4127 | n11780 ;
  assign n32151 = ~n11781 ;
  assign n11782 = x26 & n32151 ;
  assign n11783 = n30019 & n11781 ;
  assign n11784 = n11782 | n11783 ;
  assign n32152 = ~n11784 ;
  assign n11785 = n11777 & n32152 ;
  assign n32153 = ~n11777 ;
  assign n11786 = n32153 & n11784 ;
  assign n11787 = n11785 | n11786 ;
  assign n11788 = n11284 | n11286 ;
  assign n11789 = n11787 | n11788 ;
  assign n11790 = n11787 & n11788 ;
  assign n32154 = ~n11790 ;
  assign n11791 = n11789 & n32154 ;
  assign n11792 = n11288 | n11306 ;
  assign n32155 = ~n11317 ;
  assign n11793 = n32155 & n11792 ;
  assign n32156 = ~n11791 ;
  assign n11794 = n32156 & n11793 ;
  assign n32157 = ~n11793 ;
  assign n11795 = n11791 & n32157 ;
  assign n11796 = n11794 | n11795 ;
  assign n4843 = n4135 & n30385 ;
  assign n4569 = n4185 & n30361 ;
  assign n4816 = n4165 & n4811 ;
  assign n11797 = n4569 | n4816 ;
  assign n11798 = n4148 & n4664 ;
  assign n11799 = n11797 | n11798 ;
  assign n11800 = n4843 | n11799 ;
  assign n32158 = ~n11800 ;
  assign n11801 = x23 & n32158 ;
  assign n11802 = n30030 & n11800 ;
  assign n11803 = n11801 | n11802 ;
  assign n11804 = n11796 | n11803 ;
  assign n11805 = n11796 & n11803 ;
  assign n32159 = ~n11805 ;
  assign n11806 = n11804 & n32159 ;
  assign n11807 = n11319 | n11335 ;
  assign n32160 = ~n11339 ;
  assign n11808 = n32160 & n11807 ;
  assign n32161 = ~n11806 ;
  assign n11809 = n32161 & n11808 ;
  assign n32162 = ~n11808 ;
  assign n11810 = n11806 & n32162 ;
  assign n11811 = n11809 | n11810 ;
  assign n11812 = n11722 | n11811 ;
  assign n11813 = n11722 & n11811 ;
  assign n32163 = ~n11813 ;
  assign n11814 = n11812 & n32163 ;
  assign n5927 = n37300 & n30540 ;
  assign n5795 = n5191 & n30545 ;
  assign n5913 = n5144 & n30535 ;
  assign n11815 = n5795 | n5913 ;
  assign n11816 = n5166 & n30530 ;
  assign n11817 = n11815 | n11816 ;
  assign n11818 = n5927 | n11817 ;
  assign n11819 = x17 | n11818 ;
  assign n11820 = x17 & n11818 ;
  assign n32164 = ~n11820 ;
  assign n11821 = n11819 & n32164 ;
  assign n11822 = n11341 | n11359 ;
  assign n32165 = ~n11363 ;
  assign n11823 = n32165 & n11822 ;
  assign n11824 = n11821 & n11823 ;
  assign n11825 = n11821 | n11823 ;
  assign n32166 = ~n11824 ;
  assign n11826 = n32166 & n11825 ;
  assign n32167 = ~n11814 ;
  assign n11827 = n32167 & n11826 ;
  assign n32168 = ~n11826 ;
  assign n11829 = n11814 & n32168 ;
  assign n11830 = n11827 | n11829 ;
  assign n11831 = n11365 & n11390 ;
  assign n11832 = n11388 | n11831 ;
  assign n32169 = ~n11832 ;
  assign n11833 = n11830 & n32169 ;
  assign n32170 = ~n11830 ;
  assign n11834 = n32170 & n11832 ;
  assign n11835 = n11833 | n11834 ;
  assign n11836 = n11393 | n11411 ;
  assign n32171 = ~n11428 ;
  assign n11837 = n32171 & n11836 ;
  assign n32172 = ~n11835 ;
  assign n11838 = n32172 & n11837 ;
  assign n32173 = ~n11837 ;
  assign n11839 = n11835 & n32173 ;
  assign n11840 = n11838 | n11839 ;
  assign n11862 = n11455 | n11476 ;
  assign n32174 = ~n11862 ;
  assign n11863 = n11430 & n32174 ;
  assign n11864 = n11458 & n11476 ;
  assign n32175 = ~n11430 ;
  assign n11865 = n32175 & n11864 ;
  assign n11866 = n11863 | n11865 ;
  assign n32176 = ~n11840 ;
  assign n11867 = n32176 & n11866 ;
  assign n32177 = ~n11866 ;
  assign n11868 = n11840 & n32177 ;
  assign n11869 = n11867 | n11868 ;
  assign n32178 = ~n11869 ;
  assign n11870 = n895 & n32178 ;
  assign n11437 = n2849 & n11430 ;
  assign n11489 = n2861 & n11476 ;
  assign n11881 = n11437 | n11489 ;
  assign n11882 = n894 & n32176 ;
  assign n11883 = n11881 | n11882 ;
  assign n11884 = n11870 | n11883 ;
  assign n32179 = ~n11884 ;
  assign n11885 = x29 & n32179 ;
  assign n11886 = n30024 & n11884 ;
  assign n11887 = n11885 | n11886 ;
  assign n11714 = n11529 & n11713 ;
  assign n32180 = ~n11714 ;
  assign n11888 = n32180 & n11715 ;
  assign n32181 = ~n11887 ;
  assign n11889 = n32181 & n11888 ;
  assign n32182 = ~n11889 ;
  assign n11890 = n11715 & n32182 ;
  assign n11527 = n11506 | n11526 ;
  assign n11891 = n11506 & n11526 ;
  assign n32183 = ~n11891 ;
  assign n11892 = n11527 & n32183 ;
  assign n11894 = n11890 | n11892 ;
  assign n32184 = ~n11528 ;
  assign n11895 = n32184 & n11894 ;
  assign n32185 = ~n11504 ;
  assign n11896 = n32185 & n11895 ;
  assign n32186 = ~n11895 ;
  assign n11897 = n11504 & n32186 ;
  assign n11898 = n11896 | n11897 ;
  assign n6416 = n4686 & n6411 ;
  assign n4927 = n4706 & n30415 ;
  assign n5024 = n4726 & n5017 ;
  assign n11899 = n4927 | n5024 ;
  assign n11900 = n4748 & n30530 ;
  assign n11901 = n11899 | n11900 ;
  assign n11902 = n6416 | n11901 ;
  assign n32187 = ~n11902 ;
  assign n11903 = x20 & n32187 ;
  assign n11904 = n30374 & n11902 ;
  assign n11905 = n11903 | n11904 ;
  assign n4507 = n895 & n30349 ;
  assign n3702 = n2861 & n3700 ;
  assign n4105 = n894 & n4093 ;
  assign n11906 = n3702 | n4105 ;
  assign n11907 = n2849 & n30264 ;
  assign n11908 = n11906 | n11907 ;
  assign n11909 = n4507 | n11908 ;
  assign n32188 = ~n11909 ;
  assign n11910 = x29 & n32188 ;
  assign n11911 = n30024 & n11909 ;
  assign n11912 = n11910 | n11911 ;
  assign n32189 = ~n11767 ;
  assign n11913 = n11761 & n32189 ;
  assign n32190 = ~n11754 ;
  assign n11914 = n32190 & n11756 ;
  assign n11915 = n1167 | n2659 ;
  assign n11916 = n2746 | n11915 ;
  assign n11917 = n130 | n535 ;
  assign n11918 = n1726 | n11917 ;
  assign n11919 = n11916 | n11918 ;
  assign n11920 = n2049 | n11919 ;
  assign n11921 = n2973 | n2985 ;
  assign n11922 = n3188 | n11124 ;
  assign n11923 = n11921 | n11922 ;
  assign n11924 = n438 | n11923 ;
  assign n11925 = n11920 | n11924 ;
  assign n11926 = n2199 | n11925 ;
  assign n11927 = n371 | n509 ;
  assign n11928 = n542 | n11927 ;
  assign n11929 = n233 | n590 ;
  assign n11930 = n926 | n1825 ;
  assign n11931 = n11929 | n11930 ;
  assign n11932 = n11928 | n11931 ;
  assign n11933 = n573 | n808 ;
  assign n11934 = n2477 | n5764 ;
  assign n11935 = n11933 | n11934 ;
  assign n11936 = n1930 | n11935 ;
  assign n11937 = n3502 | n11936 ;
  assign n11938 = n11932 | n11937 ;
  assign n11939 = n298 | n1241 ;
  assign n11940 = n4790 | n11939 ;
  assign n11941 = n174 | n486 ;
  assign n11942 = n684 | n11941 ;
  assign n11943 = n769 | n11942 ;
  assign n11944 = n11940 | n11943 ;
  assign n11945 = n2285 | n3986 ;
  assign n11946 = n11944 | n11945 ;
  assign n11947 = n2040 | n2407 ;
  assign n11948 = n2430 | n11947 ;
  assign n11949 = n2393 | n11948 ;
  assign n11950 = n11946 | n11949 ;
  assign n11951 = n11103 | n11950 ;
  assign n11952 = n11938 | n11951 ;
  assign n11953 = n11926 | n11952 ;
  assign n11954 = n11914 | n11953 ;
  assign n11955 = n11914 & n11953 ;
  assign n32191 = ~n11955 ;
  assign n11956 = n11954 & n32191 ;
  assign n4425 = n889 & n4420 ;
  assign n3338 = n1074 & n3329 ;
  assign n3772 = n3343 & n3764 ;
  assign n11957 = n3338 | n3772 ;
  assign n11958 = n30074 & n3311 ;
  assign n11959 = n11957 | n11958 ;
  assign n11960 = n4425 | n11959 ;
  assign n32192 = ~n11960 ;
  assign n11961 = n11956 & n32192 ;
  assign n32193 = ~n11956 ;
  assign n11963 = n32193 & n11960 ;
  assign n11964 = n11961 | n11963 ;
  assign n32194 = ~n11964 ;
  assign n11965 = n11913 & n32194 ;
  assign n32195 = ~n11913 ;
  assign n11966 = n32195 & n11964 ;
  assign n11967 = n11965 | n11966 ;
  assign n32196 = ~n11912 ;
  assign n11968 = n32196 & n11967 ;
  assign n32197 = ~n11967 ;
  assign n11969 = n11912 & n32197 ;
  assign n11970 = n11968 | n11969 ;
  assign n32198 = ~n11769 ;
  assign n11971 = n32198 & n11771 ;
  assign n32199 = ~n11971 ;
  assign n11972 = n11775 & n32199 ;
  assign n11973 = n11970 & n11972 ;
  assign n11974 = n11970 | n11972 ;
  assign n32200 = ~n11973 ;
  assign n11975 = n32200 & n11974 ;
  assign n5725 = n3791 & n5723 ;
  assign n4034 = n209 & n4033 ;
  assign n4567 = n3818 & n30361 ;
  assign n11976 = n4034 | n4567 ;
  assign n11977 = n3802 & n30282 ;
  assign n11978 = n11976 | n11977 ;
  assign n11979 = n5725 | n11978 ;
  assign n32201 = ~n11979 ;
  assign n11980 = x26 & n32201 ;
  assign n11981 = n30019 & n11979 ;
  assign n11982 = n11980 | n11981 ;
  assign n32202 = ~n11982 ;
  assign n11983 = n11975 & n32202 ;
  assign n32203 = ~n11975 ;
  assign n11984 = n32203 & n11982 ;
  assign n11985 = n11983 | n11984 ;
  assign n32204 = ~n11785 ;
  assign n11986 = n32204 & n11789 ;
  assign n11987 = n11985 & n11986 ;
  assign n11988 = n11985 | n11986 ;
  assign n32205 = ~n11987 ;
  assign n11989 = n32205 & n11988 ;
  assign n6145 = n4135 & n30578 ;
  assign n4665 = n4185 & n4664 ;
  assign n4814 = n4148 & n4811 ;
  assign n11990 = n4665 | n4814 ;
  assign n11991 = n4165 & n30405 ;
  assign n11992 = n11990 | n11991 ;
  assign n11993 = n6145 | n11992 ;
  assign n32206 = ~n11993 ;
  assign n11994 = x23 & n32206 ;
  assign n11995 = n30030 & n11993 ;
  assign n11996 = n11994 | n11995 ;
  assign n32207 = ~n11996 ;
  assign n11997 = n11989 & n32207 ;
  assign n32208 = ~n11989 ;
  assign n11998 = n32208 & n11996 ;
  assign n11999 = n11997 | n11998 ;
  assign n32209 = ~n11796 ;
  assign n12000 = n32209 & n11803 ;
  assign n12001 = n11794 | n12000 ;
  assign n12002 = n11999 | n12001 ;
  assign n12003 = n11999 & n12001 ;
  assign n32210 = ~n12003 ;
  assign n12004 = n12002 & n32210 ;
  assign n32211 = ~n11905 ;
  assign n12005 = n32211 & n12004 ;
  assign n32212 = ~n12004 ;
  assign n12006 = n11905 & n32212 ;
  assign n12007 = n12005 | n12006 ;
  assign n6449 = n37300 & n6445 ;
  assign n12008 = n5144 & n30545 ;
  assign n12009 = n5166 & n30535 ;
  assign n12010 = n12008 | n12009 ;
  assign n12011 = n6449 | n12010 ;
  assign n32213 = ~n12011 ;
  assign n12012 = x17 & n32213 ;
  assign n12013 = n30580 & n12011 ;
  assign n12014 = n12012 | n12013 ;
  assign n32214 = ~n11811 ;
  assign n12015 = n11722 & n32214 ;
  assign n12016 = n11809 | n12015 ;
  assign n12017 = n12014 | n12016 ;
  assign n12018 = n12014 & n12016 ;
  assign n32215 = ~n12018 ;
  assign n12019 = n12017 & n32215 ;
  assign n32216 = ~n12007 ;
  assign n12020 = n32216 & n12019 ;
  assign n32217 = ~n12019 ;
  assign n12021 = n12007 & n32217 ;
  assign n12022 = n12020 | n12021 ;
  assign n11828 = n11814 & n11826 ;
  assign n32218 = ~n11828 ;
  assign n12023 = n11825 & n32218 ;
  assign n12025 = n12022 | n12023 ;
  assign n12024 = n12022 & n12023 ;
  assign n12026 = n11835 | n11837 ;
  assign n32219 = ~n11833 ;
  assign n12027 = n32219 & n12026 ;
  assign n12028 = n12024 | n12027 ;
  assign n12029 = n12025 & n12028 ;
  assign n6169 = n4686 & n30587 ;
  assign n4938 = n4726 & n30415 ;
  assign n5873 = n4706 & n30530 ;
  assign n12030 = n4938 | n5873 ;
  assign n12031 = n4748 & n30535 ;
  assign n12032 = n12030 | n12031 ;
  assign n12033 = n6169 | n12032 ;
  assign n32220 = ~n12033 ;
  assign n12034 = x20 & n32220 ;
  assign n12035 = n30374 & n12033 ;
  assign n12036 = n12034 | n12035 ;
  assign n5748 = n4135 & n30512 ;
  assign n4822 = n4185 & n4811 ;
  assign n5113 = n4148 & n30405 ;
  assign n12037 = n4822 | n5113 ;
  assign n12038 = n4165 & n5017 ;
  assign n12039 = n12037 | n12038 ;
  assign n12040 = n5748 | n12039 ;
  assign n32221 = ~n12040 ;
  assign n12041 = x23 & n32221 ;
  assign n12042 = n30030 & n12040 ;
  assign n12043 = n12041 | n12042 ;
  assign n12044 = n11913 & n11964 ;
  assign n12045 = n11912 & n11967 ;
  assign n12046 = n12044 | n12045 ;
  assign n4446 = n895 & n4442 ;
  assign n4035 = n894 & n4033 ;
  assign n4099 = n2849 & n4093 ;
  assign n12047 = n4035 | n4099 ;
  assign n12048 = n2861 & n30264 ;
  assign n12049 = n12047 | n12048 ;
  assign n12050 = n4446 | n12049 ;
  assign n32222 = ~n12050 ;
  assign n12051 = x29 & n32222 ;
  assign n12052 = n30024 & n12050 ;
  assign n12053 = n12051 | n12052 ;
  assign n12054 = n1471 | n1859 ;
  assign n12055 = n2718 | n11246 ;
  assign n12056 = n12054 | n12055 ;
  assign n12057 = n318 | n530 ;
  assign n12058 = n972 | n989 ;
  assign n12059 = n12057 | n12058 ;
  assign n12060 = n12056 | n12059 ;
  assign n12061 = n4558 | n12060 ;
  assign n12062 = n853 | n1665 ;
  assign n12063 = n320 | n365 ;
  assign n12064 = n2114 | n12063 ;
  assign n12065 = n3905 | n12064 ;
  assign n12066 = n12062 | n12065 ;
  assign n12067 = n2188 | n12066 ;
  assign n12068 = n12061 | n12067 ;
  assign n12069 = n2753 | n4869 ;
  assign n12070 = n12068 | n12069 ;
  assign n32223 = ~n12070 ;
  assign n12071 = n5051 & n32223 ;
  assign n32224 = ~n11953 ;
  assign n12072 = n32224 & n12071 ;
  assign n32225 = ~n12071 ;
  assign n12073 = n11953 & n32225 ;
  assign n12074 = n12072 | n12073 ;
  assign n11962 = n11954 & n32192 ;
  assign n12075 = n11955 | n11962 ;
  assign n32226 = ~n12075 ;
  assign n12076 = n12074 & n32226 ;
  assign n32227 = ~n12074 ;
  assign n12077 = n32227 & n12075 ;
  assign n12078 = n12076 | n12077 ;
  assign n3790 = n889 & n3787 ;
  assign n3324 = n1074 & n3311 ;
  assign n3707 = n3343 & n3700 ;
  assign n12079 = n3324 | n3707 ;
  assign n12080 = n3329 & n3764 ;
  assign n12081 = n12079 | n12080 ;
  assign n12082 = n3790 | n12081 ;
  assign n32228 = ~n12082 ;
  assign n12083 = n12078 & n32228 ;
  assign n32229 = ~n12078 ;
  assign n12084 = n32229 & n12082 ;
  assign n12085 = n12083 | n12084 ;
  assign n12086 = n12053 | n12085 ;
  assign n12087 = n12053 & n12085 ;
  assign n32230 = ~n12087 ;
  assign n12088 = n12086 & n32230 ;
  assign n12089 = n12046 | n12088 ;
  assign n12090 = n12046 & n12088 ;
  assign n32231 = ~n12090 ;
  assign n12091 = n12089 & n32231 ;
  assign n4677 = n3791 & n4674 ;
  assign n4566 = n3802 & n30361 ;
  assign n4666 = n3818 & n4664 ;
  assign n12092 = n4566 | n4666 ;
  assign n12093 = n209 & n30282 ;
  assign n12094 = n12092 | n12093 ;
  assign n12095 = n4677 | n12094 ;
  assign n32232 = ~n12095 ;
  assign n12096 = x26 & n32232 ;
  assign n12097 = n30019 & n12095 ;
  assign n12098 = n12096 | n12097 ;
  assign n12099 = n12091 | n12098 ;
  assign n12100 = n12091 & n12098 ;
  assign n32233 = ~n12100 ;
  assign n12101 = n12099 & n32233 ;
  assign n12102 = n11975 & n11982 ;
  assign n12103 = n11973 | n12102 ;
  assign n32234 = ~n12103 ;
  assign n12104 = n12101 & n32234 ;
  assign n32235 = ~n12101 ;
  assign n12105 = n32235 & n12103 ;
  assign n12106 = n12104 | n12105 ;
  assign n12107 = n12043 | n12106 ;
  assign n12108 = n12043 & n12106 ;
  assign n32236 = ~n12108 ;
  assign n12109 = n12107 & n32236 ;
  assign n32237 = ~n11997 ;
  assign n12110 = n11988 & n32237 ;
  assign n12111 = n12109 & n12110 ;
  assign n12112 = n12109 | n12110 ;
  assign n32238 = ~n12111 ;
  assign n12113 = n32238 & n12112 ;
  assign n12114 = n12036 | n12113 ;
  assign n12115 = n12036 & n12113 ;
  assign n32239 = ~n12115 ;
  assign n12116 = n12114 & n32239 ;
  assign n6267 = n37300 & n30597 ;
  assign n12117 = n5166 | n6267 ;
  assign n12118 = n30545 & n12117 ;
  assign n12119 = n30580 & n12118 ;
  assign n32240 = ~n12118 ;
  assign n12120 = x17 & n32240 ;
  assign n12121 = n12119 | n12120 ;
  assign n12122 = n11905 & n12004 ;
  assign n12123 = n12003 | n12122 ;
  assign n12124 = n12121 | n12123 ;
  assign n12125 = n12121 & n12123 ;
  assign n32241 = ~n12125 ;
  assign n12126 = n12124 & n32241 ;
  assign n12127 = n12116 & n12126 ;
  assign n12128 = n12116 | n12126 ;
  assign n32242 = ~n12127 ;
  assign n12129 = n32242 & n12128 ;
  assign n32243 = ~n12020 ;
  assign n12130 = n12017 & n32243 ;
  assign n32244 = ~n12129 ;
  assign n12131 = n32244 & n12130 ;
  assign n32245 = ~n12130 ;
  assign n12132 = n12129 & n32245 ;
  assign n12133 = n12131 | n12132 ;
  assign n32246 = ~n12133 ;
  assign n12134 = n12029 & n32246 ;
  assign n32247 = ~n12029 ;
  assign n12135 = n32247 & n12133 ;
  assign n12136 = n12134 | n12135 ;
  assign n32248 = ~n12024 ;
  assign n12158 = n32248 & n12025 ;
  assign n32249 = ~n12027 ;
  assign n12159 = n32249 & n12158 ;
  assign n32250 = ~n12158 ;
  assign n12160 = n12027 & n32250 ;
  assign n12161 = n12159 | n12160 ;
  assign n12183 = n11430 & n11862 ;
  assign n32251 = ~n12183 ;
  assign n12184 = n11840 & n32251 ;
  assign n12185 = n12161 & n12184 ;
  assign n12186 = n11430 | n11864 ;
  assign n12188 = n32176 & n12186 ;
  assign n32252 = ~n12161 ;
  assign n12189 = n32252 & n12188 ;
  assign n12190 = n12185 | n12189 ;
  assign n32253 = ~n12136 ;
  assign n12191 = n32253 & n12190 ;
  assign n32254 = ~n12190 ;
  assign n12192 = n12136 & n32254 ;
  assign n12193 = n12191 | n12192 ;
  assign n32255 = ~n12193 ;
  assign n12194 = n895 & n32255 ;
  assign n11852 = n2861 & n32176 ;
  assign n12165 = n2849 & n12161 ;
  assign n12205 = n11852 | n12165 ;
  assign n12206 = n894 & n32253 ;
  assign n12207 = n12205 | n12206 ;
  assign n12208 = n12194 | n12207 ;
  assign n32256 = ~n12208 ;
  assign n12209 = x29 & n32256 ;
  assign n12210 = n30024 & n12208 ;
  assign n12211 = n12209 | n12210 ;
  assign n12212 = n11898 | n12211 ;
  assign n12213 = n11898 & n12211 ;
  assign n32257 = ~n12213 ;
  assign n12214 = n12212 & n32257 ;
  assign n6166 = n4135 & n30587 ;
  assign n4937 = n4185 & n30415 ;
  assign n5876 = n4148 & n30530 ;
  assign n12215 = n4937 | n5876 ;
  assign n12216 = n4165 & n30535 ;
  assign n12217 = n12215 | n12216 ;
  assign n12218 = n6166 | n12217 ;
  assign n32258 = ~n12218 ;
  assign n12219 = x23 & n32258 ;
  assign n12220 = n30030 & n12218 ;
  assign n12221 = n12219 | n12220 ;
  assign n5746 = n3791 & n30512 ;
  assign n4825 = n209 & n4811 ;
  assign n5114 = n3802 & n30405 ;
  assign n12222 = n4825 | n5114 ;
  assign n12223 = n3818 & n5017 ;
  assign n12224 = n12222 | n12223 ;
  assign n12225 = n5746 | n12224 ;
  assign n32259 = ~n12225 ;
  assign n12226 = x26 & n32259 ;
  assign n12227 = n30019 & n12225 ;
  assign n12228 = n12226 | n12227 ;
  assign n12229 = n461 | n684 ;
  assign n12230 = n704 | n857 ;
  assign n12231 = n12229 | n12230 ;
  assign n12232 = n103 | n158 ;
  assign n12233 = n698 | n12232 ;
  assign n12234 = n955 | n12233 ;
  assign n12235 = n12231 | n12234 ;
  assign n12236 = n1378 | n1731 ;
  assign n12237 = n2252 | n5465 ;
  assign n12238 = n12236 | n12237 ;
  assign n12239 = n807 | n957 ;
  assign n12240 = n989 | n1277 ;
  assign n12241 = n12239 | n12240 ;
  assign n12242 = n12238 | n12241 ;
  assign n12243 = n3495 | n5070 ;
  assign n12244 = n12242 | n12243 ;
  assign n12245 = n12235 | n12244 ;
  assign n12246 = n5563 | n12245 ;
  assign n12247 = n4616 | n12246 ;
  assign n32260 = ~n12247 ;
  assign n12248 = n12071 & n32260 ;
  assign n12249 = n32225 & n12247 ;
  assign n12250 = n12248 | n12249 ;
  assign n12251 = x17 | n12250 ;
  assign n12252 = x17 & n12250 ;
  assign n32261 = ~n12252 ;
  assign n12253 = n12251 & n32261 ;
  assign n12254 = n11953 | n12071 ;
  assign n12255 = n12074 & n12075 ;
  assign n32262 = ~n12255 ;
  assign n12256 = n12254 & n32262 ;
  assign n12258 = n12253 | n12256 ;
  assign n12257 = n12253 & n12256 ;
  assign n32263 = ~n12257 ;
  assign n12259 = n32263 & n12258 ;
  assign n3876 = n889 & n30263 ;
  assign n3709 = n3329 & n3700 ;
  assign n3769 = n3311 & n3764 ;
  assign n12260 = n3709 | n3769 ;
  assign n12261 = n3343 & n30264 ;
  assign n12262 = n12260 | n12261 ;
  assign n12263 = n3876 | n12262 ;
  assign n32264 = ~n12263 ;
  assign n12264 = n12259 & n32264 ;
  assign n32265 = ~n12264 ;
  assign n12265 = n12258 & n32265 ;
  assign n32266 = ~n12249 ;
  assign n12266 = n32266 & n12251 ;
  assign n12267 = n651 | n4069 ;
  assign n12268 = n298 | n4047 ;
  assign n12269 = n5829 | n12268 ;
  assign n12270 = n218 | n223 ;
  assign n12271 = n539 | n12270 ;
  assign n12272 = n12269 | n12271 ;
  assign n12273 = n12267 | n12272 ;
  assign n12274 = n2169 | n2458 ;
  assign n12275 = n2628 | n12274 ;
  assign n12276 = n1807 | n12275 ;
  assign n12277 = n12273 | n12276 ;
  assign n12278 = n2977 | n12277 ;
  assign n12279 = n2453 | n4985 ;
  assign n12280 = n11145 | n12279 ;
  assign n12281 = n962 | n1105 ;
  assign n12282 = n1879 | n5550 ;
  assign n12283 = n12281 | n12282 ;
  assign n12284 = n250 | n302 ;
  assign n12285 = n833 | n1166 ;
  assign n12286 = n12284 | n12285 ;
  assign n12287 = n468 | n12286 ;
  assign n12288 = n12283 | n12287 ;
  assign n12289 = n12280 | n12288 ;
  assign n12290 = n369 | n543 ;
  assign n12291 = n239 | n12290 ;
  assign n12292 = n2531 | n12291 ;
  assign n12293 = n5839 | n11234 ;
  assign n12294 = n12292 | n12293 ;
  assign n12295 = n711 | n2030 ;
  assign n12296 = n4056 | n5071 ;
  assign n12297 = n12295 | n12296 ;
  assign n12298 = n3248 | n12297 ;
  assign n12299 = n12294 | n12298 ;
  assign n12300 = n1062 | n12299 ;
  assign n12301 = n1351 | n12300 ;
  assign n12302 = n12289 | n12301 ;
  assign n12303 = n12278 | n12302 ;
  assign n12305 = n12266 | n12303 ;
  assign n12306 = n12266 & n12303 ;
  assign n32267 = ~n12306 ;
  assign n12307 = n12305 & n32267 ;
  assign n4510 = n889 & n30349 ;
  assign n3705 = n3311 & n3700 ;
  assign n4106 = n3343 & n4093 ;
  assign n12308 = n3705 | n4106 ;
  assign n12309 = n3329 & n30264 ;
  assign n12310 = n12308 | n12309 ;
  assign n12311 = n4510 | n12310 ;
  assign n32268 = ~n12311 ;
  assign n12312 = n12307 & n32268 ;
  assign n32269 = ~n12307 ;
  assign n12314 = n32269 & n12311 ;
  assign n12315 = n12312 | n12314 ;
  assign n12316 = n12265 | n12315 ;
  assign n5728 = n895 & n5723 ;
  assign n3944 = n2849 & n30282 ;
  assign n4568 = n894 & n30361 ;
  assign n12317 = n3944 | n4568 ;
  assign n12318 = n2861 & n4033 ;
  assign n12319 = n12317 | n12318 ;
  assign n12320 = n5728 | n12319 ;
  assign n12321 = x29 | n12320 ;
  assign n12322 = x29 & n12320 ;
  assign n32270 = ~n12322 ;
  assign n12323 = n12321 & n32270 ;
  assign n12324 = n12265 & n12315 ;
  assign n32271 = ~n12324 ;
  assign n12325 = n12316 & n32271 ;
  assign n32272 = ~n12323 ;
  assign n12327 = n32272 & n12325 ;
  assign n32273 = ~n12327 ;
  assign n12328 = n12316 & n32273 ;
  assign n12329 = n2348 | n3124 ;
  assign n12330 = n3922 | n12329 ;
  assign n12331 = n3199 | n12330 ;
  assign n12332 = n383 | n441 ;
  assign n12333 = n1278 | n12332 ;
  assign n12334 = n3549 | n12333 ;
  assign n12335 = n12331 | n12334 ;
  assign n12336 = n257 | n273 ;
  assign n12337 = n996 | n12336 ;
  assign n12338 = n2241 | n2427 ;
  assign n12339 = n4074 | n12338 ;
  assign n12340 = n12337 | n12339 ;
  assign n12341 = n272 | n767 ;
  assign n12342 = n1179 | n12341 ;
  assign n12343 = n344 | n1694 ;
  assign n12344 = n12342 | n12343 ;
  assign n12345 = n5062 | n12344 ;
  assign n12346 = n3138 | n12345 ;
  assign n12347 = n12340 | n12346 ;
  assign n12348 = n12335 | n12347 ;
  assign n12349 = n353 | n359 ;
  assign n12350 = n381 | n849 ;
  assign n12351 = n12349 | n12350 ;
  assign n32274 = ~n12351 ;
  assign n12352 = n633 & n32274 ;
  assign n32275 = ~n3129 ;
  assign n12353 = n32275 & n12352 ;
  assign n12354 = n162 | n376 ;
  assign n12355 = n233 | n12354 ;
  assign n12356 = n2472 | n12355 ;
  assign n12357 = n5466 | n12356 ;
  assign n12358 = n2145 | n12357 ;
  assign n12359 = n3995 | n12358 ;
  assign n32276 = ~n12359 ;
  assign n12360 = n12353 & n32276 ;
  assign n32277 = ~n3174 ;
  assign n12361 = n32277 & n12360 ;
  assign n32278 = ~n12348 ;
  assign n12362 = n32278 & n12361 ;
  assign n12363 = n12303 | n12362 ;
  assign n12364 = n12303 & n12362 ;
  assign n32279 = ~n12364 ;
  assign n12365 = n12363 & n32279 ;
  assign n4447 = n889 & n4442 ;
  assign n3864 = n3311 & n30264 ;
  assign n4103 = n3329 & n4093 ;
  assign n12366 = n3864 | n4103 ;
  assign n12367 = n3343 & n4033 ;
  assign n12368 = n12366 | n12367 ;
  assign n12369 = n4447 | n12368 ;
  assign n32280 = ~n12369 ;
  assign n12370 = n12365 & n32280 ;
  assign n32281 = ~n12365 ;
  assign n12372 = n32281 & n12369 ;
  assign n12373 = n12370 | n12372 ;
  assign n12313 = n12305 & n32268 ;
  assign n12374 = n12306 | n12313 ;
  assign n12375 = n12373 | n12374 ;
  assign n12376 = n12373 & n12374 ;
  assign n32282 = ~n12376 ;
  assign n12377 = n12375 & n32282 ;
  assign n12378 = n12328 | n12377 ;
  assign n12379 = n12328 & n12377 ;
  assign n32283 = ~n12379 ;
  assign n12380 = n12378 & n32283 ;
  assign n4678 = n895 & n4674 ;
  assign n3940 = n2861 & n30282 ;
  assign n4572 = n2849 & n30361 ;
  assign n12381 = n3940 | n4572 ;
  assign n12382 = n894 & n4664 ;
  assign n12383 = n12381 | n12382 ;
  assign n12384 = n4678 | n12383 ;
  assign n12385 = x29 | n12384 ;
  assign n12386 = x29 & n12384 ;
  assign n32284 = ~n12386 ;
  assign n12387 = n12385 & n32284 ;
  assign n32285 = ~n12380 ;
  assign n12388 = n32285 & n12387 ;
  assign n32286 = ~n12387 ;
  assign n12389 = n12380 & n32286 ;
  assign n12390 = n12388 | n12389 ;
  assign n12391 = n12228 | n12390 ;
  assign n12392 = n12228 & n12390 ;
  assign n32287 = ~n12392 ;
  assign n12393 = n12391 & n32287 ;
  assign n12326 = n12323 & n12325 ;
  assign n12394 = n12323 | n12325 ;
  assign n32288 = ~n12326 ;
  assign n12395 = n32288 & n12394 ;
  assign n32289 = ~n12259 ;
  assign n12396 = n32289 & n12263 ;
  assign n12397 = n12264 | n12396 ;
  assign n4126 = n895 & n30286 ;
  assign n3945 = n894 & n30282 ;
  assign n4098 = n2861 & n4093 ;
  assign n12398 = n3945 | n4098 ;
  assign n12399 = n2849 & n4033 ;
  assign n12400 = n12398 | n12399 ;
  assign n12401 = n4126 | n12400 ;
  assign n32290 = ~n12401 ;
  assign n12402 = x29 & n32290 ;
  assign n12403 = n30024 & n12401 ;
  assign n12404 = n12402 | n12403 ;
  assign n12405 = n12397 | n12404 ;
  assign n12406 = n12397 & n12404 ;
  assign n32291 = ~n12406 ;
  assign n12407 = n12405 & n32291 ;
  assign n32292 = ~n12085 ;
  assign n12408 = n12053 & n32292 ;
  assign n12409 = n12084 | n12408 ;
  assign n32293 = ~n12409 ;
  assign n12410 = n12407 & n32293 ;
  assign n32294 = ~n12410 ;
  assign n12411 = n12405 & n32294 ;
  assign n12412 = n12395 & n12411 ;
  assign n6146 = n3791 & n30578 ;
  assign n4668 = n209 & n4664 ;
  assign n4815 = n3802 & n4811 ;
  assign n12413 = n4668 | n4815 ;
  assign n12414 = n3818 & n30405 ;
  assign n12415 = n12413 | n12414 ;
  assign n12416 = n6146 | n12415 ;
  assign n12417 = x26 | n12416 ;
  assign n12418 = x26 & n12416 ;
  assign n32295 = ~n12418 ;
  assign n12419 = n12417 & n32295 ;
  assign n12420 = n12395 | n12411 ;
  assign n32296 = ~n12412 ;
  assign n12421 = n32296 & n12420 ;
  assign n12422 = n12419 & n12421 ;
  assign n12423 = n12412 | n12422 ;
  assign n32297 = ~n12423 ;
  assign n12424 = n12393 & n32297 ;
  assign n32298 = ~n12393 ;
  assign n12425 = n32298 & n12423 ;
  assign n12426 = n12424 | n12425 ;
  assign n12427 = n12221 | n12426 ;
  assign n12428 = n12221 & n12426 ;
  assign n32299 = ~n12428 ;
  assign n12429 = n12427 & n32299 ;
  assign n6269 = n4686 & n30597 ;
  assign n12430 = n4726 | n6269 ;
  assign n12431 = n30545 & n12430 ;
  assign n12432 = x20 & n12431 ;
  assign n12433 = x20 | n12431 ;
  assign n32300 = ~n12432 ;
  assign n12434 = n32300 & n12433 ;
  assign n12435 = n12419 | n12421 ;
  assign n32301 = ~n12422 ;
  assign n12436 = n32301 & n12435 ;
  assign n32302 = ~n12407 ;
  assign n12437 = n32302 & n12409 ;
  assign n12438 = n12410 | n12437 ;
  assign n32303 = ~n12088 ;
  assign n12439 = n12046 & n32303 ;
  assign n32304 = ~n12091 ;
  assign n12440 = n32304 & n12098 ;
  assign n12441 = n12439 | n12440 ;
  assign n12442 = n12438 | n12441 ;
  assign n12443 = n12438 & n12441 ;
  assign n32305 = ~n12443 ;
  assign n12444 = n12442 & n32305 ;
  assign n4842 = n3791 & n30385 ;
  assign n4578 = n209 & n30361 ;
  assign n4818 = n3818 & n4811 ;
  assign n12445 = n4578 | n4818 ;
  assign n12446 = n3802 & n4664 ;
  assign n12447 = n12445 | n12446 ;
  assign n12448 = n4842 | n12447 ;
  assign n32306 = ~n12448 ;
  assign n12449 = x26 & n32306 ;
  assign n12450 = n30019 & n12448 ;
  assign n12451 = n12449 | n12450 ;
  assign n32307 = ~n12451 ;
  assign n12452 = n12444 & n32307 ;
  assign n32308 = ~n12452 ;
  assign n12453 = n12442 & n32308 ;
  assign n12454 = n12436 & n12453 ;
  assign n6417 = n4135 & n6411 ;
  assign n4931 = n4148 & n30415 ;
  assign n5020 = n4185 & n5017 ;
  assign n12455 = n4931 | n5020 ;
  assign n12456 = n4165 & n30530 ;
  assign n12457 = n12455 | n12456 ;
  assign n12458 = n6417 | n12457 ;
  assign n32309 = ~n12458 ;
  assign n12459 = x23 & n32309 ;
  assign n12460 = n30030 & n12458 ;
  assign n12461 = n12459 | n12460 ;
  assign n12462 = n12436 | n12453 ;
  assign n32310 = ~n12454 ;
  assign n12463 = n32310 & n12462 ;
  assign n12465 = n12461 & n12463 ;
  assign n12466 = n12454 | n12465 ;
  assign n32311 = ~n12466 ;
  assign n12467 = n12434 & n32311 ;
  assign n32312 = ~n12434 ;
  assign n12468 = n32312 & n12466 ;
  assign n12469 = n12467 | n12468 ;
  assign n32313 = ~n12429 ;
  assign n12470 = n32313 & n12469 ;
  assign n32314 = ~n12469 ;
  assign n12471 = n12429 & n32314 ;
  assign n12472 = n12470 | n12471 ;
  assign n6450 = n4686 & n6445 ;
  assign n12473 = n4706 & n30545 ;
  assign n12474 = n4726 & n30535 ;
  assign n12475 = n12473 | n12474 ;
  assign n12476 = n6450 | n12475 ;
  assign n12477 = x20 | n12476 ;
  assign n12478 = x20 & n12476 ;
  assign n32315 = ~n12478 ;
  assign n12479 = n12477 & n32315 ;
  assign n32316 = ~n12444 ;
  assign n12480 = n32316 & n12451 ;
  assign n12481 = n12452 | n12480 ;
  assign n32317 = ~n12104 ;
  assign n12482 = n32317 & n12107 ;
  assign n12484 = n12481 | n12482 ;
  assign n32318 = ~n12481 ;
  assign n12483 = n32318 & n12482 ;
  assign n32319 = ~n12482 ;
  assign n12485 = n12481 & n32319 ;
  assign n12486 = n12483 | n12485 ;
  assign n5138 = n4135 & n30410 ;
  assign n4929 = n4165 & n30415 ;
  assign n5108 = n4185 & n30405 ;
  assign n12487 = n4929 | n5108 ;
  assign n12488 = n4148 & n5017 ;
  assign n12489 = n12487 | n12488 ;
  assign n12490 = n5138 | n12489 ;
  assign n32320 = ~n12490 ;
  assign n12491 = x23 & n32320 ;
  assign n12492 = n30030 & n12490 ;
  assign n12493 = n12491 | n12492 ;
  assign n32321 = ~n12493 ;
  assign n12494 = n12486 & n32321 ;
  assign n32322 = ~n12494 ;
  assign n12495 = n12484 & n32322 ;
  assign n12497 = n12479 | n12495 ;
  assign n32323 = ~n12461 ;
  assign n12464 = n32323 & n12463 ;
  assign n32324 = ~n12463 ;
  assign n12498 = n12461 & n32324 ;
  assign n12499 = n12464 | n12498 ;
  assign n12496 = n12479 & n12495 ;
  assign n32325 = ~n12496 ;
  assign n12500 = n32325 & n12497 ;
  assign n32326 = ~n12499 ;
  assign n12502 = n32326 & n12500 ;
  assign n32327 = ~n12502 ;
  assign n12503 = n12497 & n32327 ;
  assign n12504 = n12472 & n12503 ;
  assign n12505 = n12472 | n12503 ;
  assign n32328 = ~n12504 ;
  assign n12506 = n32328 & n12505 ;
  assign n12501 = n12499 & n12500 ;
  assign n12507 = n12499 | n12500 ;
  assign n32329 = ~n12501 ;
  assign n12508 = n32329 & n12507 ;
  assign n32330 = ~n12486 ;
  assign n12509 = n32330 & n12493 ;
  assign n12510 = n12494 | n12509 ;
  assign n32331 = ~n12109 ;
  assign n12511 = n32331 & n12110 ;
  assign n32332 = ~n12113 ;
  assign n12512 = n12036 & n32332 ;
  assign n12513 = n12511 | n12512 ;
  assign n12514 = n12510 | n12513 ;
  assign n12515 = n12510 & n12513 ;
  assign n32333 = ~n12515 ;
  assign n12516 = n12514 & n32333 ;
  assign n5928 = n4686 & n30540 ;
  assign n5796 = n4748 & n30545 ;
  assign n5874 = n4726 & n30530 ;
  assign n12517 = n5796 | n5874 ;
  assign n12518 = n4706 & n30535 ;
  assign n12519 = n12517 | n12518 ;
  assign n12520 = n5928 | n12519 ;
  assign n32334 = ~n12520 ;
  assign n12521 = x20 & n32334 ;
  assign n12522 = n30374 & n12520 ;
  assign n12523 = n12521 | n12522 ;
  assign n32335 = ~n12523 ;
  assign n12524 = n12516 & n32335 ;
  assign n32336 = ~n12524 ;
  assign n12525 = n12514 & n32336 ;
  assign n12527 = n12508 | n12525 ;
  assign n12526 = n12508 & n12525 ;
  assign n32337 = ~n12516 ;
  assign n12528 = n32337 & n12523 ;
  assign n12529 = n12524 | n12528 ;
  assign n12530 = n12124 & n32242 ;
  assign n12532 = n12529 | n12530 ;
  assign n32338 = ~n12529 ;
  assign n12531 = n32338 & n12530 ;
  assign n32339 = ~n12530 ;
  assign n12533 = n12529 & n32339 ;
  assign n12534 = n12531 | n12533 ;
  assign n12535 = n12029 | n12133 ;
  assign n32340 = ~n12132 ;
  assign n12536 = n32340 & n12535 ;
  assign n32341 = ~n12536 ;
  assign n12538 = n12534 & n32341 ;
  assign n32342 = ~n12538 ;
  assign n12539 = n12532 & n32342 ;
  assign n12540 = n12526 | n12539 ;
  assign n12541 = n12527 & n12540 ;
  assign n32343 = ~n12506 ;
  assign n12542 = n32343 & n12541 ;
  assign n32344 = ~n12541 ;
  assign n12543 = n12506 & n32344 ;
  assign n12544 = n12542 | n12543 ;
  assign n32345 = ~n12526 ;
  assign n12567 = n32345 & n12527 ;
  assign n32346 = ~n12539 ;
  assign n12568 = n32346 & n12567 ;
  assign n32347 = ~n12567 ;
  assign n12569 = n12539 & n32347 ;
  assign n12570 = n12568 | n12569 ;
  assign n12537 = n12534 & n12536 ;
  assign n12594 = n12534 | n12536 ;
  assign n32348 = ~n12537 ;
  assign n12595 = n32348 & n12594 ;
  assign n12622 = n12161 | n12188 ;
  assign n12623 = n32253 & n12622 ;
  assign n12624 = n12595 | n12623 ;
  assign n32349 = ~n12624 ;
  assign n12625 = n12570 & n32349 ;
  assign n32350 = ~n12184 ;
  assign n12617 = n12161 & n32350 ;
  assign n32351 = ~n12617 ;
  assign n12619 = n12136 & n32351 ;
  assign n32352 = ~n12619 ;
  assign n12621 = n12595 & n32352 ;
  assign n32353 = ~n12570 ;
  assign n12626 = n32353 & n12621 ;
  assign n12627 = n12625 | n12626 ;
  assign n32354 = ~n12544 ;
  assign n12628 = n32354 & n12627 ;
  assign n32355 = ~n12627 ;
  assign n12629 = n12544 & n32355 ;
  assign n12630 = n12628 | n12629 ;
  assign n32356 = ~n12630 ;
  assign n12631 = n3791 & n32356 ;
  assign n12586 = n3802 & n12570 ;
  assign n12610 = n209 & n12595 ;
  assign n12641 = n12586 | n12610 ;
  assign n12642 = n3818 & n32354 ;
  assign n12643 = n12641 | n12642 ;
  assign n12644 = n12631 | n12643 ;
  assign n12645 = x26 | n12644 ;
  assign n12646 = x26 & n12644 ;
  assign n32357 = ~n12646 ;
  assign n12647 = n12645 & n32357 ;
  assign n32358 = ~n11892 ;
  assign n11893 = n11890 & n32358 ;
  assign n32359 = ~n11890 ;
  assign n12648 = n32359 & n11892 ;
  assign n12649 = n11893 | n12648 ;
  assign n12187 = n11840 | n12186 ;
  assign n12650 = n11840 & n12183 ;
  assign n32360 = ~n12650 ;
  assign n12651 = n12187 & n32360 ;
  assign n32361 = ~n12651 ;
  assign n12652 = n12161 & n32361 ;
  assign n12653 = n32252 & n12651 ;
  assign n12654 = n12652 | n12653 ;
  assign n32362 = ~n12654 ;
  assign n12655 = n895 & n32362 ;
  assign n11439 = n2861 & n11430 ;
  assign n11842 = n2849 & n32176 ;
  assign n12666 = n11439 | n11842 ;
  assign n12667 = n894 & n12161 ;
  assign n12668 = n12666 | n12667 ;
  assign n12669 = n12655 | n12668 ;
  assign n12670 = x29 | n12669 ;
  assign n12671 = x29 & n12669 ;
  assign n32363 = ~n12671 ;
  assign n12672 = n12670 & n32363 ;
  assign n32364 = ~n12672 ;
  assign n12674 = n12649 & n32364 ;
  assign n12673 = n12649 & n12672 ;
  assign n12675 = n12649 | n12672 ;
  assign n32365 = ~n12673 ;
  assign n12676 = n32365 & n12675 ;
  assign n12620 = n12595 & n12619 ;
  assign n32366 = ~n12595 ;
  assign n12677 = n32366 & n12623 ;
  assign n12678 = n12620 | n12677 ;
  assign n12679 = n12570 & n12678 ;
  assign n12680 = n12570 | n12678 ;
  assign n32367 = ~n12679 ;
  assign n12681 = n32367 & n12680 ;
  assign n12682 = n3791 & n12681 ;
  assign n12138 = n209 & n32253 ;
  assign n12608 = n3802 & n12595 ;
  assign n12692 = n12138 | n12608 ;
  assign n12693 = n3818 & n12570 ;
  assign n12694 = n12692 | n12693 ;
  assign n12695 = n12682 | n12694 ;
  assign n32368 = ~n12695 ;
  assign n12696 = x26 & n32368 ;
  assign n12697 = n30019 & n12695 ;
  assign n12698 = n12696 | n12697 ;
  assign n12699 = n12676 | n12698 ;
  assign n32369 = ~n12674 ;
  assign n12700 = n32369 & n12699 ;
  assign n12701 = n12647 & n12700 ;
  assign n12702 = n12647 | n12700 ;
  assign n32370 = ~n12701 ;
  assign n12703 = n32370 & n12702 ;
  assign n12704 = n12214 & n12703 ;
  assign n12705 = n12214 | n12703 ;
  assign n32371 = ~n12704 ;
  assign n12706 = n32371 & n12705 ;
  assign n6418 = n3791 & n6411 ;
  assign n4930 = n3802 & n30415 ;
  assign n5021 = n209 & n5017 ;
  assign n12707 = n4930 | n5021 ;
  assign n12708 = n3818 & n30530 ;
  assign n12709 = n12707 | n12708 ;
  assign n12710 = n6418 | n12709 ;
  assign n32372 = ~n12710 ;
  assign n12711 = x26 & n32372 ;
  assign n12712 = n30019 & n12710 ;
  assign n12713 = n12711 | n12712 ;
  assign n6147 = n895 & n30578 ;
  assign n4813 = n2849 & n4811 ;
  assign n5115 = n894 & n30405 ;
  assign n12714 = n4813 | n5115 ;
  assign n12715 = n2861 & n4664 ;
  assign n12716 = n12714 | n12715 ;
  assign n12717 = n6147 | n12716 ;
  assign n32373 = ~n12717 ;
  assign n12718 = x29 & n32373 ;
  assign n12719 = n30024 & n12717 ;
  assign n12720 = n12718 | n12719 ;
  assign n32374 = ~n12303 ;
  assign n12304 = x20 & n32374 ;
  assign n12721 = n30374 & n12303 ;
  assign n12722 = n12304 | n12721 ;
  assign n12723 = n113 | n570 ;
  assign n12724 = n2472 | n12723 ;
  assign n12725 = n255 | n636 ;
  assign n12726 = n133 | n474 ;
  assign n12727 = n3016 | n12726 ;
  assign n12728 = n12725 | n12727 ;
  assign n12729 = n12724 | n12728 ;
  assign n12730 = n1050 | n2229 ;
  assign n12731 = n130 | n479 ;
  assign n12732 = n816 | n996 ;
  assign n12733 = n12731 | n12732 ;
  assign n12734 = n12730 | n12733 ;
  assign n12735 = n383 | n509 ;
  assign n12736 = n683 | n12735 ;
  assign n12737 = n367 | n12736 ;
  assign n12738 = n12734 | n12737 ;
  assign n12739 = n332 | n430 ;
  assign n12740 = n550 | n12739 ;
  assign n12741 = n2559 | n3496 ;
  assign n12742 = n12740 | n12741 ;
  assign n12743 = n924 | n4650 ;
  assign n12744 = n12742 | n12743 ;
  assign n12745 = n12738 | n12744 ;
  assign n12746 = n12729 | n12745 ;
  assign n12747 = n124 | n2993 ;
  assign n12748 = n5294 | n12747 ;
  assign n12749 = n292 | n1199 ;
  assign n12750 = n568 | n764 ;
  assign n12751 = n857 | n1010 ;
  assign n12752 = n12750 | n12751 ;
  assign n12753 = n187 | n269 ;
  assign n12754 = n296 | n327 ;
  assign n12755 = n12753 | n12754 ;
  assign n12756 = n12752 | n12755 ;
  assign n12757 = n12749 | n12756 ;
  assign n12758 = n12748 | n12757 ;
  assign n12759 = n171 | n439 ;
  assign n12760 = n610 | n12759 ;
  assign n12761 = n2389 | n2768 ;
  assign n12762 = n12760 | n12761 ;
  assign n12763 = n138 | n334 ;
  assign n12764 = n460 | n12763 ;
  assign n12765 = n595 | n12764 ;
  assign n12766 = n12762 | n12765 ;
  assign n12767 = n221 | n301 ;
  assign n12768 = n376 | n591 ;
  assign n12769 = n12767 | n12768 ;
  assign n12770 = n2277 | n12769 ;
  assign n12771 = n4636 | n12770 ;
  assign n12772 = n225 | n1469 ;
  assign n12773 = n2749 | n12772 ;
  assign n12774 = n5098 | n12773 ;
  assign n12775 = n12771 | n12774 ;
  assign n12776 = n12766 | n12775 ;
  assign n12777 = n12758 | n12776 ;
  assign n12778 = n12746 | n12777 ;
  assign n12779 = n3441 | n12778 ;
  assign n12780 = n12722 | n12779 ;
  assign n12781 = n12722 & n12779 ;
  assign n32375 = ~n12781 ;
  assign n12782 = n12780 & n32375 ;
  assign n4128 = n889 & n30286 ;
  assign n3946 = n3343 & n30282 ;
  assign n4101 = n3311 & n4093 ;
  assign n12783 = n3946 | n4101 ;
  assign n12784 = n3329 & n4033 ;
  assign n12785 = n12783 | n12784 ;
  assign n12786 = n4128 | n12785 ;
  assign n32376 = ~n12786 ;
  assign n12788 = n12782 & n32376 ;
  assign n12787 = n12782 | n12786 ;
  assign n12789 = n12782 & n12786 ;
  assign n32377 = ~n12789 ;
  assign n12790 = n12787 & n32377 ;
  assign n12371 = n12363 & n32280 ;
  assign n12791 = n12364 | n12371 ;
  assign n32378 = ~n12790 ;
  assign n12793 = n32378 & n12791 ;
  assign n12794 = n12788 | n12793 ;
  assign n32379 = ~n12722 ;
  assign n12795 = n32379 & n12779 ;
  assign n12796 = n12721 | n12795 ;
  assign n12797 = n179 | n283 ;
  assign n12798 = n950 | n12797 ;
  assign n12799 = n1104 | n12798 ;
  assign n12800 = n12267 | n12799 ;
  assign n12801 = n263 | n668 ;
  assign n12802 = n814 | n12801 ;
  assign n12803 = n751 | n1248 ;
  assign n12804 = n12802 | n12803 ;
  assign n12805 = n2472 | n4016 ;
  assign n12806 = n12804 | n12805 ;
  assign n12807 = n157 | n477 ;
  assign n12808 = n1047 | n12807 ;
  assign n12809 = n2410 | n12808 ;
  assign n12810 = n1689 | n2900 ;
  assign n32380 = ~n12810 ;
  assign n12811 = n3892 & n32380 ;
  assign n32381 = ~n12809 ;
  assign n12812 = n32381 & n12811 ;
  assign n32382 = ~n12806 ;
  assign n12813 = n32382 & n12812 ;
  assign n32383 = ~n12800 ;
  assign n12814 = n32383 & n12813 ;
  assign n32384 = ~n3681 ;
  assign n12815 = n32384 & n12814 ;
  assign n12816 = n220 | n793 ;
  assign n12817 = n335 | n682 ;
  assign n12818 = n845 | n12817 ;
  assign n12819 = n12816 | n12818 ;
  assign n12820 = n1547 | n12819 ;
  assign n12821 = n2487 | n12820 ;
  assign n12822 = n345 | n767 ;
  assign n12823 = n237 | n12822 ;
  assign n12824 = n766 | n946 ;
  assign n12825 = n1152 | n2887 ;
  assign n12826 = n12824 | n12825 ;
  assign n12827 = n12823 | n12826 ;
  assign n12828 = n301 | n323 ;
  assign n12829 = n199 | n12828 ;
  assign n12830 = n833 | n12829 ;
  assign n12831 = n857 | n996 ;
  assign n12832 = n4859 | n4997 ;
  assign n12833 = n12831 | n12832 ;
  assign n12834 = n12830 | n12833 ;
  assign n12835 = n12827 | n12834 ;
  assign n12836 = n12821 | n12835 ;
  assign n12837 = n459 | n12836 ;
  assign n32385 = ~n12837 ;
  assign n12838 = n12815 & n32385 ;
  assign n12839 = n12796 & n12838 ;
  assign n12840 = n12796 | n12838 ;
  assign n32386 = ~n12839 ;
  assign n12841 = n32386 & n12840 ;
  assign n5729 = n889 & n5723 ;
  assign n3939 = n3329 & n30282 ;
  assign n4576 = n3343 & n30361 ;
  assign n12842 = n3939 | n4576 ;
  assign n12843 = n3311 & n4033 ;
  assign n12844 = n12842 | n12843 ;
  assign n12845 = n5729 | n12844 ;
  assign n32387 = ~n12845 ;
  assign n12846 = n12841 & n32387 ;
  assign n32388 = ~n12841 ;
  assign n12848 = n32388 & n12845 ;
  assign n12849 = n12846 | n12848 ;
  assign n12850 = n12794 | n12849 ;
  assign n12851 = n12794 & n12849 ;
  assign n32389 = ~n12851 ;
  assign n12852 = n12850 & n32389 ;
  assign n12853 = n12720 | n12852 ;
  assign n12854 = n12720 & n12852 ;
  assign n32390 = ~n12854 ;
  assign n12855 = n12853 & n32390 ;
  assign n12792 = n12790 | n12791 ;
  assign n12856 = n12790 & n12791 ;
  assign n32391 = ~n12856 ;
  assign n12857 = n12792 & n32391 ;
  assign n32392 = ~n12373 ;
  assign n12858 = n32392 & n12374 ;
  assign n32393 = ~n12858 ;
  assign n12859 = n12378 & n32393 ;
  assign n12861 = n12857 | n12859 ;
  assign n4841 = n895 & n30385 ;
  assign n4579 = n2861 & n30361 ;
  assign n4812 = n894 & n4811 ;
  assign n12862 = n4579 | n4812 ;
  assign n12863 = n2849 & n4664 ;
  assign n12864 = n12862 | n12863 ;
  assign n12865 = n4841 | n12864 ;
  assign n12866 = x29 | n12865 ;
  assign n12867 = x29 & n12865 ;
  assign n32394 = ~n12867 ;
  assign n12868 = n12866 & n32394 ;
  assign n32395 = ~n12857 ;
  assign n12860 = n32395 & n12859 ;
  assign n32396 = ~n12859 ;
  assign n12869 = n12857 & n32396 ;
  assign n12870 = n12860 | n12869 ;
  assign n32397 = ~n12868 ;
  assign n12872 = n32397 & n12870 ;
  assign n32398 = ~n12872 ;
  assign n12873 = n12861 & n32398 ;
  assign n12874 = n12855 & n12873 ;
  assign n12875 = n12855 | n12873 ;
  assign n32399 = ~n12874 ;
  assign n12876 = n32399 & n12875 ;
  assign n12877 = n12713 | n12876 ;
  assign n12878 = n12713 & n12876 ;
  assign n32400 = ~n12878 ;
  assign n12879 = n12877 & n32400 ;
  assign n6451 = n4135 & n6445 ;
  assign n12880 = n4148 & n30545 ;
  assign n12881 = n4185 & n30535 ;
  assign n12882 = n12880 | n12881 ;
  assign n12883 = n6451 | n12882 ;
  assign n12884 = x23 | n12883 ;
  assign n12885 = x23 & n12883 ;
  assign n32401 = ~n12885 ;
  assign n12886 = n12884 & n32401 ;
  assign n12887 = n12879 & n12886 ;
  assign n12888 = n12879 | n12886 ;
  assign n32402 = ~n12887 ;
  assign n12889 = n32402 & n12888 ;
  assign n12871 = n12868 & n12870 ;
  assign n12890 = n12868 | n12870 ;
  assign n32403 = ~n12871 ;
  assign n12891 = n32403 & n12890 ;
  assign n32404 = ~n12389 ;
  assign n12892 = n32404 & n12391 ;
  assign n12893 = n12891 & n12892 ;
  assign n12894 = n12891 | n12892 ;
  assign n32405 = ~n12893 ;
  assign n12895 = n32405 & n12894 ;
  assign n5140 = n3791 & n30410 ;
  assign n4928 = n3818 & n30415 ;
  assign n5023 = n3802 & n5017 ;
  assign n12896 = n4928 | n5023 ;
  assign n12897 = n209 & n30405 ;
  assign n12898 = n12896 | n12897 ;
  assign n12899 = n5140 | n12898 ;
  assign n32406 = ~n12899 ;
  assign n12900 = x26 & n32406 ;
  assign n12901 = n30019 & n12899 ;
  assign n12902 = n12900 | n12901 ;
  assign n12904 = n12895 & n12902 ;
  assign n12905 = n12893 | n12904 ;
  assign n12906 = n12889 | n12905 ;
  assign n12907 = n12889 & n12905 ;
  assign n32407 = ~n12907 ;
  assign n12908 = n12906 & n32407 ;
  assign n32408 = ~n12902 ;
  assign n12903 = n12895 & n32408 ;
  assign n32409 = ~n12895 ;
  assign n12909 = n32409 & n12902 ;
  assign n12910 = n12903 | n12909 ;
  assign n5929 = n4135 & n30540 ;
  assign n5797 = n4165 & n30545 ;
  assign n5871 = n4185 & n30530 ;
  assign n12911 = n5797 | n5871 ;
  assign n12912 = n4148 & n30535 ;
  assign n12913 = n12911 | n12912 ;
  assign n12914 = n5929 | n12913 ;
  assign n32410 = ~n12914 ;
  assign n12915 = x23 & n32410 ;
  assign n12916 = n30030 & n12914 ;
  assign n12917 = n12915 | n12916 ;
  assign n12919 = n12910 | n12917 ;
  assign n32411 = ~n12917 ;
  assign n12918 = n12910 & n32411 ;
  assign n32412 = ~n12910 ;
  assign n12920 = n32412 & n12917 ;
  assign n12921 = n12918 | n12920 ;
  assign n32413 = ~n12426 ;
  assign n12922 = n12221 & n32413 ;
  assign n12923 = n12425 | n12922 ;
  assign n32414 = ~n12923 ;
  assign n12925 = n12921 & n32414 ;
  assign n32415 = ~n12925 ;
  assign n12926 = n12919 & n32415 ;
  assign n32416 = ~n12926 ;
  assign n12928 = n12908 & n32416 ;
  assign n32417 = ~n12908 ;
  assign n12927 = n32417 & n12926 ;
  assign n12924 = n12921 | n12923 ;
  assign n12929 = n12921 & n12923 ;
  assign n32418 = ~n12929 ;
  assign n12930 = n12924 & n32418 ;
  assign n12931 = n12434 | n12466 ;
  assign n12932 = n12429 & n12469 ;
  assign n32419 = ~n12932 ;
  assign n12933 = n12931 & n32419 ;
  assign n12935 = n12930 | n12933 ;
  assign n12934 = n12930 & n12933 ;
  assign n32420 = ~n12472 ;
  assign n12936 = n32420 & n12503 ;
  assign n12937 = n12542 | n12936 ;
  assign n12938 = n12934 | n12937 ;
  assign n12939 = n12935 & n12938 ;
  assign n12940 = n12927 | n12939 ;
  assign n32421 = ~n12928 ;
  assign n12941 = n32421 & n12940 ;
  assign n6165 = n3791 & n30587 ;
  assign n4926 = n209 & n30415 ;
  assign n5914 = n3818 & n30535 ;
  assign n12942 = n4926 | n5914 ;
  assign n12943 = n3802 & n30530 ;
  assign n12944 = n12942 | n12943 ;
  assign n12945 = n6165 | n12944 ;
  assign n12946 = x26 | n12945 ;
  assign n12947 = x26 & n12945 ;
  assign n32422 = ~n12947 ;
  assign n12948 = n12946 & n32422 ;
  assign n32423 = ~n12849 ;
  assign n12949 = n12794 & n32423 ;
  assign n32424 = ~n12949 ;
  assign n12950 = n12853 & n32424 ;
  assign n12951 = n344 | n474 ;
  assign n12952 = n83 | n542 ;
  assign n12953 = n621 | n12952 ;
  assign n12954 = n12951 | n12953 ;
  assign n12955 = n90 | n176 ;
  assign n12956 = n250 | n12955 ;
  assign n12957 = n1865 | n3736 ;
  assign n12958 = n12956 | n12957 ;
  assign n12959 = n3455 | n12958 ;
  assign n12960 = n12954 | n12959 ;
  assign n12961 = n346 | n355 ;
  assign n12962 = n461 | n543 ;
  assign n12963 = n12961 | n12962 ;
  assign n12964 = n412 | n12963 ;
  assign n12965 = n2265 | n12964 ;
  assign n12966 = n223 | n433 ;
  assign n12967 = n453 | n495 ;
  assign n12968 = n12966 | n12967 ;
  assign n12969 = n1390 | n12968 ;
  assign n12970 = n2315 | n12969 ;
  assign n12971 = n12965 | n12970 ;
  assign n12972 = n12960 | n12971 ;
  assign n12973 = n1090 | n12972 ;
  assign n12974 = n11571 | n12973 ;
  assign n32425 = ~n12974 ;
  assign n12975 = n12838 & n32425 ;
  assign n32426 = ~n12838 ;
  assign n12977 = n32426 & n12974 ;
  assign n12978 = n12975 | n12977 ;
  assign n12847 = n12839 | n12845 ;
  assign n12979 = n12840 & n12847 ;
  assign n32427 = ~n12978 ;
  assign n12980 = n32427 & n12979 ;
  assign n32428 = ~n12979 ;
  assign n12981 = n12978 & n32428 ;
  assign n12982 = n12980 | n12981 ;
  assign n4679 = n889 & n4674 ;
  assign n3947 = n3311 & n30282 ;
  assign n4573 = n3329 & n30361 ;
  assign n12983 = n3947 | n4573 ;
  assign n12984 = n3343 & n4664 ;
  assign n12985 = n12983 | n12984 ;
  assign n12986 = n4679 | n12985 ;
  assign n12987 = n12982 | n12986 ;
  assign n12988 = n12982 & n12986 ;
  assign n32429 = ~n12988 ;
  assign n12989 = n12987 & n32429 ;
  assign n12990 = n12950 & n12989 ;
  assign n12991 = n12950 | n12989 ;
  assign n32430 = ~n12990 ;
  assign n12992 = n32430 & n12991 ;
  assign n5745 = n895 & n30512 ;
  assign n4828 = n2861 & n4811 ;
  assign n5106 = n2849 & n30405 ;
  assign n12993 = n4828 | n5106 ;
  assign n12994 = n894 & n5017 ;
  assign n12995 = n12993 | n12994 ;
  assign n12996 = n5745 | n12995 ;
  assign n12997 = x29 | n12996 ;
  assign n12998 = x29 & n12996 ;
  assign n32431 = ~n12998 ;
  assign n12999 = n12997 & n32431 ;
  assign n13000 = n12992 & n12999 ;
  assign n13001 = n12992 | n12999 ;
  assign n32432 = ~n13000 ;
  assign n13002 = n32432 & n13001 ;
  assign n13003 = n12948 & n13002 ;
  assign n13004 = n12948 | n13002 ;
  assign n32433 = ~n13003 ;
  assign n13005 = n32433 & n13004 ;
  assign n6270 = n4135 & n30597 ;
  assign n13006 = n4185 | n6270 ;
  assign n13007 = n30545 & n13006 ;
  assign n13008 = n30030 & n13007 ;
  assign n32434 = ~n13007 ;
  assign n13009 = x23 & n32434 ;
  assign n13010 = n13008 | n13009 ;
  assign n32435 = ~n12855 ;
  assign n13011 = n32435 & n12873 ;
  assign n32436 = ~n12876 ;
  assign n13012 = n12713 & n32436 ;
  assign n13013 = n13011 | n13012 ;
  assign n13014 = n13010 | n13013 ;
  assign n13015 = n13010 & n13013 ;
  assign n32437 = ~n13015 ;
  assign n13016 = n13014 & n32437 ;
  assign n32438 = ~n13005 ;
  assign n13017 = n32438 & n13016 ;
  assign n32439 = ~n13016 ;
  assign n13018 = n13005 & n32439 ;
  assign n13019 = n13017 | n13018 ;
  assign n32440 = ~n12886 ;
  assign n13020 = n12879 & n32440 ;
  assign n32441 = ~n13020 ;
  assign n13021 = n12906 & n32441 ;
  assign n13022 = n13019 & n13021 ;
  assign n13023 = n13019 | n13021 ;
  assign n32442 = ~n13022 ;
  assign n13024 = n32442 & n13023 ;
  assign n32443 = ~n12941 ;
  assign n13025 = n32443 & n13024 ;
  assign n32444 = ~n13024 ;
  assign n13026 = n12941 & n32444 ;
  assign n13027 = n13025 | n13026 ;
  assign n13049 = n12927 | n12928 ;
  assign n32445 = ~n13049 ;
  assign n13050 = n12939 & n32445 ;
  assign n32446 = ~n12939 ;
  assign n13051 = n32446 & n13049 ;
  assign n13052 = n13050 | n13051 ;
  assign n32447 = ~n12934 ;
  assign n13074 = n32447 & n12935 ;
  assign n32448 = ~n12937 ;
  assign n13075 = n32448 & n13074 ;
  assign n32449 = ~n13074 ;
  assign n13076 = n12937 & n32449 ;
  assign n13077 = n13075 | n13076 ;
  assign n13099 = n12570 | n12621 ;
  assign n13101 = n32354 & n13099 ;
  assign n13102 = n13077 | n13101 ;
  assign n13103 = n13052 | n13102 ;
  assign n13104 = n12570 & n12624 ;
  assign n32450 = ~n13104 ;
  assign n13105 = n12544 & n32450 ;
  assign n32451 = ~n13105 ;
  assign n13107 = n13077 & n32451 ;
  assign n13108 = n13052 & n13107 ;
  assign n32452 = ~n13108 ;
  assign n13109 = n13103 & n32452 ;
  assign n32453 = ~n13109 ;
  assign n13110 = n13027 & n32453 ;
  assign n32454 = ~n13027 ;
  assign n13111 = n32454 & n13109 ;
  assign n13112 = n13110 | n13111 ;
  assign n32455 = ~n13112 ;
  assign n13114 = n4135 & n32455 ;
  assign n32456 = ~n13052 ;
  assign n13057 = n4148 & n32456 ;
  assign n13088 = n4185 & n13077 ;
  assign n13124 = n13057 | n13088 ;
  assign n13125 = n4165 & n13027 ;
  assign n13126 = n13124 | n13125 ;
  assign n13127 = n13114 | n13126 ;
  assign n32457 = ~n13127 ;
  assign n13128 = x23 & n32457 ;
  assign n13129 = n30030 & n13127 ;
  assign n13130 = n13128 | n13129 ;
  assign n32458 = ~n13130 ;
  assign n13131 = n12706 & n32458 ;
  assign n32459 = ~n12706 ;
  assign n13132 = n32459 & n13130 ;
  assign n13133 = n13131 | n13132 ;
  assign n13134 = n12676 & n12698 ;
  assign n32460 = ~n13134 ;
  assign n13135 = n12699 & n32460 ;
  assign n32461 = ~n11888 ;
  assign n13136 = n11887 & n32461 ;
  assign n13137 = n11889 | n13136 ;
  assign n13138 = n11709 & n11711 ;
  assign n32462 = ~n13138 ;
  assign n13139 = n11712 & n32462 ;
  assign n11467 = n895 & n11463 ;
  assign n10660 = n2861 & n10656 ;
  assign n11487 = n2849 & n11476 ;
  assign n13140 = n10660 | n11487 ;
  assign n13141 = n894 & n11430 ;
  assign n13142 = n13140 | n13141 ;
  assign n13143 = n11467 | n13142 ;
  assign n32463 = ~n13143 ;
  assign n13144 = x29 & n32463 ;
  assign n13145 = n30024 & n13143 ;
  assign n13146 = n13144 | n13145 ;
  assign n32464 = ~n13146 ;
  assign n13147 = n13139 & n32464 ;
  assign n32465 = ~n13139 ;
  assign n13148 = n32465 & n13146 ;
  assign n13149 = n13147 | n13148 ;
  assign n11707 = n11591 & n11706 ;
  assign n32466 = ~n11707 ;
  assign n13150 = n32466 & n11708 ;
  assign n32467 = ~n7416 ;
  assign n10645 = n32467 & n10643 ;
  assign n13151 = n10645 | n10646 ;
  assign n32468 = ~n13151 ;
  assign n13152 = n11010 & n32468 ;
  assign n32469 = ~n11023 ;
  assign n13153 = n32469 & n13151 ;
  assign n13154 = n13152 | n13153 ;
  assign n13155 = n10681 & n13154 ;
  assign n13156 = n10681 | n13154 ;
  assign n32470 = ~n13155 ;
  assign n13157 = n32470 & n13156 ;
  assign n13158 = n889 & n13157 ;
  assign n10722 = n3329 & n10703 ;
  assign n10740 = n3311 & n10727 ;
  assign n13169 = n10722 | n10740 ;
  assign n13170 = n3343 & n10681 ;
  assign n13171 = n13169 | n13170 ;
  assign n13172 = n13158 | n13171 ;
  assign n32471 = ~n13172 ;
  assign n13173 = n13150 & n32471 ;
  assign n32472 = ~n13150 ;
  assign n13174 = n32472 & n13172 ;
  assign n13175 = n13173 | n13174 ;
  assign n32473 = ~n11617 ;
  assign n13176 = n32473 & n11704 ;
  assign n13177 = n11705 | n13176 ;
  assign n11009 = n10727 & n11008 ;
  assign n13178 = n32124 & n11022 ;
  assign n13179 = n11009 | n13178 ;
  assign n13180 = n10703 & n13179 ;
  assign n13181 = n10703 | n13179 ;
  assign n32474 = ~n13180 ;
  assign n13182 = n32474 & n13181 ;
  assign n13183 = n889 & n13182 ;
  assign n10738 = n3329 & n10727 ;
  assign n10761 = n3311 & n31999 ;
  assign n13194 = n10738 | n10761 ;
  assign n13195 = n3343 & n13151 ;
  assign n13196 = n13194 | n13195 ;
  assign n13197 = n13183 | n13196 ;
  assign n13199 = n13177 & n13197 ;
  assign n13200 = n1435 | n2030 ;
  assign n13201 = n2558 | n4556 ;
  assign n13202 = n13200 | n13201 ;
  assign n13203 = n327 | n359 ;
  assign n13204 = n507 | n13203 ;
  assign n13205 = n2148 | n13204 ;
  assign n13206 = n13202 | n13205 ;
  assign n13207 = n2516 | n12743 ;
  assign n13208 = n13206 | n13207 ;
  assign n13209 = n540 | n2475 ;
  assign n13210 = n159 | n241 ;
  assign n13211 = n542 | n13210 ;
  assign n13212 = n1367 | n13211 ;
  assign n13213 = n13209 | n13212 ;
  assign n13214 = n289 | n372 ;
  assign n13215 = n512 | n13214 ;
  assign n13216 = n124 | n900 ;
  assign n13217 = n2905 | n13216 ;
  assign n13218 = n13215 | n13217 ;
  assign n13219 = n2173 | n13218 ;
  assign n13220 = n13213 | n13219 ;
  assign n13221 = n13208 | n13220 ;
  assign n13222 = n4091 | n11238 ;
  assign n13223 = n13221 | n13222 ;
  assign n11006 = n10773 & n11005 ;
  assign n32475 = ~n10773 ;
  assign n13224 = n32475 & n11020 ;
  assign n13225 = n11006 | n13224 ;
  assign n13226 = n31999 & n13225 ;
  assign n32476 = ~n13225 ;
  assign n13227 = n10750 & n32476 ;
  assign n13228 = n13226 | n13227 ;
  assign n32477 = ~n13228 ;
  assign n13229 = n889 & n32477 ;
  assign n10782 = n3329 & n10773 ;
  assign n10807 = n3311 & n31998 ;
  assign n13240 = n10782 | n10807 ;
  assign n32478 = ~n11680 ;
  assign n13241 = n3343 & n32478 ;
  assign n13242 = n13240 | n13241 ;
  assign n13243 = n13229 | n13242 ;
  assign n13244 = n13223 | n13243 ;
  assign n13245 = n13223 & n13243 ;
  assign n32479 = ~n13245 ;
  assign n13246 = n13244 & n32479 ;
  assign n13247 = n151 | n978 ;
  assign n13248 = n356 | n13247 ;
  assign n13249 = n2426 | n2559 ;
  assign n13250 = n13248 | n13249 ;
  assign n13251 = n3906 | n13250 ;
  assign n13252 = n497 | n528 ;
  assign n13253 = n12831 | n13252 ;
  assign n13254 = n214 | n495 ;
  assign n13255 = n348 | n721 ;
  assign n13256 = n13254 | n13255 ;
  assign n13257 = n13253 | n13256 ;
  assign n13258 = n2323 | n13257 ;
  assign n13259 = n13251 | n13258 ;
  assign n13260 = n613 | n1044 ;
  assign n13261 = n2749 | n4652 ;
  assign n13262 = n13260 | n13261 ;
  assign n13263 = n679 | n750 ;
  assign n13264 = n816 | n13263 ;
  assign n13265 = n90 | n190 ;
  assign n13266 = n301 | n608 ;
  assign n13267 = n13265 | n13266 ;
  assign n13268 = n13264 | n13267 ;
  assign n13269 = n13262 | n13268 ;
  assign n13270 = n4271 | n13269 ;
  assign n13271 = n13259 | n13270 ;
  assign n13272 = n1780 | n13271 ;
  assign n13273 = n4001 | n13272 ;
  assign n13274 = n10795 & n11004 ;
  assign n13275 = n10795 | n11019 ;
  assign n32480 = ~n13274 ;
  assign n13276 = n32480 & n13275 ;
  assign n32481 = ~n13276 ;
  assign n13277 = n10773 & n32481 ;
  assign n13278 = n32475 & n13276 ;
  assign n13279 = n13277 | n13278 ;
  assign n32482 = ~n13279 ;
  assign n13282 = n889 & n32482 ;
  assign n10806 = n3329 & n31998 ;
  assign n10827 = n3311 & n10818 ;
  assign n13293 = n10806 | n10827 ;
  assign n32483 = ~n8614 ;
  assign n13291 = n32483 & n10635 ;
  assign n13292 = n10636 | n13291 ;
  assign n13294 = n3343 & n13292 ;
  assign n13295 = n13293 | n13294 ;
  assign n13296 = n13282 | n13295 ;
  assign n13297 = n13273 | n13296 ;
  assign n13298 = n13273 & n13296 ;
  assign n32484 = ~n13298 ;
  assign n13299 = n13297 & n32484 ;
  assign n13300 = n643 | n1438 ;
  assign n13301 = n2594 | n11127 ;
  assign n13302 = n13300 | n13301 ;
  assign n13303 = n216 | n464 ;
  assign n13304 = n476 | n795 ;
  assign n13305 = n13303 | n13304 ;
  assign n13306 = n1537 | n1731 ;
  assign n13307 = n13305 | n13306 ;
  assign n13308 = n5807 | n13307 ;
  assign n13309 = n13302 | n13308 ;
  assign n13310 = n2675 | n13309 ;
  assign n13311 = n1640 | n13310 ;
  assign n13312 = n11640 | n13311 ;
  assign n32485 = ~n11002 ;
  assign n11003 = n10818 & n32485 ;
  assign n32486 = ~n10818 ;
  assign n13313 = n32486 & n11018 ;
  assign n13314 = n11003 | n13313 ;
  assign n13315 = n31998 & n13314 ;
  assign n32487 = ~n13314 ;
  assign n13316 = n10795 & n32487 ;
  assign n13317 = n13315 | n13316 ;
  assign n32488 = ~n13317 ;
  assign n13318 = n889 & n32488 ;
  assign n10830 = n3329 & n10818 ;
  assign n10855 = n3311 & n10841 ;
  assign n13329 = n10830 | n10855 ;
  assign n13330 = n3343 & n31998 ;
  assign n13331 = n13329 | n13330 ;
  assign n13332 = n13318 | n13331 ;
  assign n13334 = n13312 & n13332 ;
  assign n13333 = n13312 | n13332 ;
  assign n32489 = ~n13334 ;
  assign n13335 = n13333 & n32489 ;
  assign n13336 = n495 | n1002 ;
  assign n13337 = n3098 | n13336 ;
  assign n13338 = n2122 | n2412 ;
  assign n13339 = n2746 | n13338 ;
  assign n13340 = n3042 | n13339 ;
  assign n13341 = n13337 | n13340 ;
  assign n13342 = n480 | n814 ;
  assign n13343 = n1152 | n13342 ;
  assign n13344 = n12349 | n13343 ;
  assign n13345 = n5805 | n13344 ;
  assign n13346 = n270 | n506 ;
  assign n13347 = n658 | n961 ;
  assign n13348 = n13346 | n13347 ;
  assign n13349 = n278 | n1500 ;
  assign n13350 = n13348 | n13349 ;
  assign n13351 = n433 | n897 ;
  assign n13352 = n3887 | n13351 ;
  assign n13353 = n13350 | n13352 ;
  assign n13354 = n1359 | n13353 ;
  assign n13355 = n13345 | n13354 ;
  assign n13356 = n13341 | n13355 ;
  assign n13357 = n5546 | n13356 ;
  assign n13358 = n181 | n248 ;
  assign n13359 = n293 | n13358 ;
  assign n13360 = n905 | n1422 ;
  assign n13361 = n1859 | n13360 ;
  assign n13362 = n13359 | n13361 ;
  assign n13363 = n564 | n635 ;
  assign n13364 = n839 | n13363 ;
  assign n13365 = n298 | n1174 ;
  assign n13366 = n13364 | n13365 ;
  assign n13367 = n1067 | n1438 ;
  assign n13368 = n13366 | n13367 ;
  assign n13369 = n1513 | n1860 ;
  assign n13370 = n3503 | n13369 ;
  assign n13371 = n5606 | n13370 ;
  assign n13372 = n13368 | n13371 ;
  assign n13373 = n13362 | n13372 ;
  assign n13374 = n5057 | n12758 ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = n13357 | n13375 ;
  assign n32490 = ~n10841 ;
  assign n13377 = n32490 & n11001 ;
  assign n32491 = ~n11017 ;
  assign n13378 = n10841 & n32491 ;
  assign n13379 = n13377 | n13378 ;
  assign n13380 = n10818 & n13379 ;
  assign n13381 = n10818 | n13379 ;
  assign n32492 = ~n13380 ;
  assign n13382 = n32492 & n13381 ;
  assign n13383 = n889 & n13382 ;
  assign n10854 = n3329 & n10841 ;
  assign n10872 = n3311 & n10865 ;
  assign n13394 = n10854 | n10872 ;
  assign n13395 = n3343 & n10818 ;
  assign n13396 = n13394 | n13395 ;
  assign n13397 = n13383 | n13396 ;
  assign n13398 = n13376 | n13397 ;
  assign n13399 = n13376 & n13397 ;
  assign n32493 = ~n13399 ;
  assign n13400 = n13398 & n32493 ;
  assign n13401 = n217 | n461 ;
  assign n13402 = n647 | n13401 ;
  assign n13403 = n240 | n327 ;
  assign n13404 = n516 | n591 ;
  assign n13405 = n13403 | n13404 ;
  assign n13406 = n1285 | n13405 ;
  assign n13407 = n13402 | n13406 ;
  assign n13408 = n1389 | n11246 ;
  assign n13409 = n290 | n4056 ;
  assign n13410 = n4967 | n13409 ;
  assign n13411 = n12742 | n13410 ;
  assign n13412 = n13408 | n13411 ;
  assign n13413 = n13407 | n13412 ;
  assign n13414 = n5413 | n13413 ;
  assign n13415 = n921 | n1681 ;
  assign n13416 = n302 | n560 ;
  assign n13417 = n381 | n13416 ;
  assign n13418 = n875 | n2182 ;
  assign n13419 = n13417 | n13418 ;
  assign n13420 = n5606 | n13419 ;
  assign n13421 = n13415 | n13420 ;
  assign n13422 = n499 | n2628 ;
  assign n13423 = n3234 | n5822 ;
  assign n13424 = n13422 | n13423 ;
  assign n13425 = n5810 | n13424 ;
  assign n13426 = n13421 | n13425 ;
  assign n13427 = n358 | n500 ;
  assign n13428 = n661 | n13427 ;
  assign n13429 = n1718 | n13428 ;
  assign n13430 = n1697 | n2716 ;
  assign n13431 = n3579 | n12727 ;
  assign n13432 = n13430 | n13431 ;
  assign n13433 = n13429 | n13432 ;
  assign n13434 = n400 | n479 ;
  assign n13435 = n5384 | n13434 ;
  assign n13436 = n2474 | n5317 ;
  assign n13437 = n13435 | n13436 ;
  assign n13438 = n1154 | n2394 ;
  assign n13439 = n90 | n788 ;
  assign n13440 = n3078 | n13439 ;
  assign n13441 = n13438 | n13440 ;
  assign n13442 = n337 | n440 ;
  assign n13443 = n538 | n13442 ;
  assign n13444 = n447 | n1865 ;
  assign n13445 = n13443 | n13444 ;
  assign n13446 = n2450 | n13445 ;
  assign n13447 = n13441 | n13446 ;
  assign n13448 = n13437 | n13447 ;
  assign n13449 = n13433 | n13448 ;
  assign n13450 = n13426 | n13449 ;
  assign n13451 = n13414 | n13450 ;
  assign n11000 = n10865 & n10999 ;
  assign n32494 = ~n10865 ;
  assign n13452 = n32494 & n11016 ;
  assign n13453 = n11000 | n13452 ;
  assign n13454 = n10841 & n13453 ;
  assign n13455 = n10841 | n13453 ;
  assign n32495 = ~n13454 ;
  assign n13456 = n32495 & n13455 ;
  assign n13457 = n889 & n13456 ;
  assign n10874 = n3329 & n10865 ;
  assign n10898 = n3311 & n10892 ;
  assign n13467 = n10874 | n10898 ;
  assign n13468 = n3343 & n10841 ;
  assign n13469 = n13467 | n13468 ;
  assign n13470 = n13457 | n13469 ;
  assign n13471 = n13451 | n13470 ;
  assign n13472 = n13451 & n13470 ;
  assign n32496 = ~n13472 ;
  assign n13473 = n13471 & n32496 ;
  assign n13474 = n304 | n367 ;
  assign n13475 = n249 | n289 ;
  assign n13476 = n395 | n13475 ;
  assign n13477 = n982 | n13476 ;
  assign n13478 = n13474 | n13477 ;
  assign n13479 = n912 | n2517 ;
  assign n13480 = n2768 | n13479 ;
  assign n13481 = n469 | n506 ;
  assign n13482 = n554 | n564 ;
  assign n13483 = n13481 | n13482 ;
  assign n13484 = n766 | n846 ;
  assign n13485 = n13483 | n13484 ;
  assign n13486 = n13480 | n13485 ;
  assign n13487 = n13478 | n13486 ;
  assign n32497 = ~n13487 ;
  assign n13488 = n149 & n32497 ;
  assign n32498 = ~n1140 ;
  assign n13489 = n32498 & n13488 ;
  assign n13490 = n402 | n688 ;
  assign n13491 = n1423 | n11576 ;
  assign n13492 = n13490 | n13491 ;
  assign n13493 = n176 | n560 ;
  assign n13494 = n336 | n13493 ;
  assign n13495 = n3573 | n13494 ;
  assign n13496 = n3753 | n4019 ;
  assign n13497 = n13495 | n13496 ;
  assign n13498 = n13492 | n13497 ;
  assign n13499 = n770 | n1100 ;
  assign n13500 = n3247 | n4285 ;
  assign n13501 = n353 | n451 ;
  assign n13502 = n12732 | n13501 ;
  assign n13503 = n13500 | n13502 ;
  assign n13504 = n1686 | n13503 ;
  assign n13505 = n13499 | n13504 ;
  assign n13506 = n157 | n290 ;
  assign n13507 = n3729 | n12231 ;
  assign n13508 = n13506 | n13507 ;
  assign n13509 = n587 | n1142 ;
  assign n13510 = n1415 | n1943 ;
  assign n13511 = n13509 | n13510 ;
  assign n13512 = n164 | n296 ;
  assign n13513 = n471 | n13512 ;
  assign n13514 = n13511 | n13513 ;
  assign n13515 = n13508 | n13514 ;
  assign n13516 = n13505 | n13515 ;
  assign n13517 = n13498 | n13516 ;
  assign n32499 = ~n13517 ;
  assign n13518 = n13489 & n32499 ;
  assign n13519 = n10892 | n10998 ;
  assign n13520 = n10892 & n11015 ;
  assign n32500 = ~n13520 ;
  assign n13521 = n13519 & n32500 ;
  assign n32501 = ~n13521 ;
  assign n13522 = n10865 & n32501 ;
  assign n13523 = n32494 & n13521 ;
  assign n13524 = n13522 | n13523 ;
  assign n32502 = ~n13524 ;
  assign n13525 = n889 & n32502 ;
  assign n10905 = n3329 & n10892 ;
  assign n32503 = ~n10917 ;
  assign n10929 = n3311 & n32503 ;
  assign n13536 = n10905 | n10929 ;
  assign n13537 = n3343 & n10865 ;
  assign n13538 = n13536 | n13537 ;
  assign n13539 = n13525 | n13538 ;
  assign n32504 = ~n13539 ;
  assign n13540 = n13518 & n32504 ;
  assign n32505 = ~n13518 ;
  assign n13541 = n32505 & n13539 ;
  assign n13542 = n13540 | n13541 ;
  assign n32506 = ~n10994 ;
  assign n10995 = n6562 & n32506 ;
  assign n13544 = n31995 & n10992 ;
  assign n13545 = n108 & n13544 ;
  assign n13547 = n10995 | n13545 ;
  assign n10987 = n6561 & n10974 ;
  assign n13543 = n3329 | n10987 ;
  assign n32507 = ~n10992 ;
  assign n13548 = n32507 & n13543 ;
  assign n13549 = n13547 | n13548 ;
  assign n13550 = n360 | n698 ;
  assign n13551 = n3578 | n13550 ;
  assign n13552 = n372 | n445 ;
  assign n13553 = n508 | n13552 ;
  assign n13554 = n5839 | n13553 ;
  assign n13555 = n13551 | n13554 ;
  assign n13556 = n971 | n1423 ;
  assign n13557 = n1922 | n13556 ;
  assign n13558 = n5301 | n13557 ;
  assign n13559 = n13555 | n13558 ;
  assign n13560 = n495 | n651 ;
  assign n13561 = n281 | n13560 ;
  assign n13562 = n97 | n300 ;
  assign n13563 = n466 | n13562 ;
  assign n13564 = n13561 | n13563 ;
  assign n13565 = n1067 | n13564 ;
  assign n13566 = n4892 | n13362 ;
  assign n13567 = n13565 | n13566 ;
  assign n13568 = n13559 | n13567 ;
  assign n13569 = n257 | n278 ;
  assign n13570 = n1293 | n2224 ;
  assign n13571 = n358 | n399 ;
  assign n13572 = n660 | n682 ;
  assign n13573 = n13571 | n13572 ;
  assign n13574 = n13570 | n13573 ;
  assign n13575 = n13569 | n13574 ;
  assign n13576 = n2088 | n4982 ;
  assign n13577 = n13575 | n13576 ;
  assign n13578 = n1993 | n2012 ;
  assign n13579 = n13577 | n13578 ;
  assign n13580 = n5469 | n13579 ;
  assign n32508 = ~n13580 ;
  assign n13581 = n2332 & n32508 ;
  assign n32509 = ~n13568 ;
  assign n13582 = n32509 & n13581 ;
  assign n32510 = ~n13582 ;
  assign n13584 = n13549 & n32510 ;
  assign n13585 = n1101 | n1229 ;
  assign n13586 = n4804 | n13585 ;
  assign n13587 = n157 | n179 ;
  assign n13588 = n508 | n1252 ;
  assign n13589 = n13587 | n13588 ;
  assign n13590 = n823 | n900 ;
  assign n13591 = n13589 | n13590 ;
  assign n13592 = n13586 | n13591 ;
  assign n13593 = n112 | n380 ;
  assign n13594 = n961 | n13593 ;
  assign n13595 = n2204 | n13594 ;
  assign n13596 = n2615 | n13595 ;
  assign n13597 = n13592 | n13596 ;
  assign n13598 = n256 | n429 ;
  assign n13599 = n749 | n1271 ;
  assign n13600 = n13598 | n13599 ;
  assign n13601 = n1837 | n13600 ;
  assign n13602 = n13597 | n13601 ;
  assign n32511 = ~n13602 ;
  assign n13603 = n646 & n32511 ;
  assign n13604 = n301 | n368 ;
  assign n13605 = n434 | n13604 ;
  assign n13606 = n1032 | n2226 ;
  assign n13607 = n13605 | n13606 ;
  assign n13608 = n214 | n695 ;
  assign n13609 = n1293 | n13608 ;
  assign n13610 = n1370 | n1859 ;
  assign n13611 = n13609 | n13610 ;
  assign n13612 = n2135 | n13611 ;
  assign n13613 = n13499 | n13612 ;
  assign n13614 = n13607 | n13613 ;
  assign n13615 = n1160 | n1857 ;
  assign n13616 = n13572 | n13615 ;
  assign n13617 = n151 | n241 ;
  assign n13618 = n474 | n679 ;
  assign n13619 = n13617 | n13618 ;
  assign n13620 = n1853 | n13619 ;
  assign n13621 = n13616 | n13620 ;
  assign n13622 = n5052 | n13621 ;
  assign n13623 = n2920 | n4534 ;
  assign n13624 = n279 | n486 ;
  assign n13625 = n1199 | n13624 ;
  assign n13626 = n4955 | n13625 ;
  assign n13627 = n13623 | n13626 ;
  assign n13628 = n11668 | n13627 ;
  assign n13629 = n13622 | n13628 ;
  assign n13630 = n13614 | n13629 ;
  assign n32512 = ~n13630 ;
  assign n13631 = n13603 & n32512 ;
  assign n32513 = ~n13631 ;
  assign n13633 = n13584 & n32513 ;
  assign n13632 = n13584 & n13631 ;
  assign n13634 = n13584 | n13631 ;
  assign n32514 = ~n13632 ;
  assign n13635 = n32514 & n13634 ;
  assign n13546 = n10940 & n13544 ;
  assign n13636 = n10940 | n13544 ;
  assign n32515 = ~n13546 ;
  assign n13637 = n32515 & n13636 ;
  assign n13638 = n889 & n13637 ;
  assign n13639 = n3343 & n10940 ;
  assign n13640 = n3329 & n31995 ;
  assign n13641 = n3311 & n32507 ;
  assign n13642 = n13640 | n13641 ;
  assign n13643 = n13639 | n13642 ;
  assign n13644 = n13638 | n13643 ;
  assign n32516 = ~n13635 ;
  assign n13646 = n32516 & n13644 ;
  assign n13647 = n13633 | n13646 ;
  assign n13648 = n186 | n434 ;
  assign n13649 = n767 | n13648 ;
  assign n13650 = n1860 | n2113 ;
  assign n13651 = n13649 | n13650 ;
  assign n13652 = n5535 | n12764 ;
  assign n13653 = n13651 | n13652 ;
  assign n13654 = n4886 | n5363 ;
  assign n13655 = n13653 | n13654 ;
  assign n13656 = n2603 | n3190 ;
  assign n13657 = n13655 | n13656 ;
  assign n13658 = n906 | n965 ;
  assign n13659 = n422 | n11191 ;
  assign n13660 = n3151 | n13659 ;
  assign n13661 = n13658 | n13660 ;
  assign n13662 = n1435 | n1731 ;
  assign n13663 = n3281 | n4303 ;
  assign n13664 = n13662 | n13663 ;
  assign n13665 = n103 | n401 ;
  assign n13666 = n1252 | n13665 ;
  assign n13667 = n595 | n13666 ;
  assign n13668 = n13664 | n13667 ;
  assign n13669 = n13661 | n13668 ;
  assign n13670 = n159 | n377 ;
  assign n13671 = n116 | n13670 ;
  assign n13672 = n2477 | n4963 ;
  assign n13673 = n13671 | n13672 ;
  assign n13674 = n534 | n795 ;
  assign n13675 = n978 | n13674 ;
  assign n13676 = n1276 | n13675 ;
  assign n13677 = n3997 | n5905 ;
  assign n13678 = n13676 | n13677 ;
  assign n13679 = n13673 | n13678 ;
  assign n13680 = n13669 | n13679 ;
  assign n13681 = n13657 | n13680 ;
  assign n13682 = n3441 | n13681 ;
  assign n13684 = n13647 & n13682 ;
  assign n13683 = n13647 | n13682 ;
  assign n32517 = ~n13684 ;
  assign n13685 = n13683 & n32517 ;
  assign n10988 = n10940 & n10974 ;
  assign n13686 = n10940 | n10994 ;
  assign n32518 = ~n10988 ;
  assign n13687 = n32518 & n13686 ;
  assign n13688 = n10917 | n13687 ;
  assign n13689 = n10917 & n13687 ;
  assign n32519 = ~n13689 ;
  assign n13690 = n13688 & n32519 ;
  assign n13691 = n889 & n13690 ;
  assign n10962 = n3329 & n10940 ;
  assign n10977 = n3311 & n31995 ;
  assign n13702 = n10962 | n10977 ;
  assign n13703 = n3343 & n32503 ;
  assign n13704 = n13702 | n13703 ;
  assign n13705 = n13691 | n13704 ;
  assign n13707 = n13685 & n13705 ;
  assign n13708 = n13684 | n13707 ;
  assign n13709 = n811 | n839 ;
  assign n13710 = n358 | n1206 ;
  assign n13711 = n13709 | n13710 ;
  assign n13712 = n472 | n5886 ;
  assign n13713 = n13711 | n13712 ;
  assign n13714 = n320 | n12725 ;
  assign n13715 = n418 | n704 ;
  assign n32520 = ~n13715 ;
  assign n13716 = n5047 & n32520 ;
  assign n32521 = ~n13714 ;
  assign n13717 = n32521 & n13716 ;
  assign n13718 = n1050 | n2071 ;
  assign n13719 = n3015 | n4872 ;
  assign n13720 = n13718 | n13719 ;
  assign n13721 = n199 | n500 ;
  assign n13722 = n453 | n991 ;
  assign n13723 = n13721 | n13722 ;
  assign n13724 = n13720 | n13723 ;
  assign n13725 = n273 | n827 ;
  assign n13726 = n1129 | n1766 ;
  assign n13727 = n13725 | n13726 ;
  assign n13728 = n399 | n410 ;
  assign n13729 = n439 | n13728 ;
  assign n13730 = n11556 | n13729 ;
  assign n13731 = n13727 | n13730 ;
  assign n13732 = n13724 | n13731 ;
  assign n32522 = ~n13732 ;
  assign n13733 = n13717 & n32522 ;
  assign n32523 = ~n13713 ;
  assign n13734 = n32523 & n13733 ;
  assign n13735 = n486 | n816 ;
  assign n13736 = n116 | n13735 ;
  assign n13737 = n398 | n13736 ;
  assign n13738 = n477 | n1136 ;
  assign n13739 = n1279 | n13738 ;
  assign n13740 = n13737 | n13739 ;
  assign n13741 = n131 | n344 ;
  assign n13742 = n530 | n13741 ;
  assign n13743 = n3970 | n13742 ;
  assign n13744 = n11188 | n13743 ;
  assign n13745 = n13740 | n13744 ;
  assign n13746 = n2238 | n13745 ;
  assign n13747 = n1400 | n13746 ;
  assign n32524 = ~n13747 ;
  assign n13748 = n13734 & n32524 ;
  assign n32525 = ~n13748 ;
  assign n13750 = n13708 & n32525 ;
  assign n32526 = ~n13708 ;
  assign n13749 = n32526 & n13748 ;
  assign n13751 = n13749 | n13750 ;
  assign n10997 = n32503 & n10996 ;
  assign n13752 = n10917 & n10975 ;
  assign n13753 = n10997 | n13752 ;
  assign n13754 = n10892 & n13753 ;
  assign n13755 = n10892 | n13753 ;
  assign n32527 = ~n13754 ;
  assign n13756 = n32527 & n13755 ;
  assign n13757 = n889 & n13756 ;
  assign n10932 = n3329 & n32503 ;
  assign n10964 = n3311 & n10940 ;
  assign n13768 = n10932 | n10964 ;
  assign n13769 = n3343 & n10892 ;
  assign n13770 = n13768 | n13769 ;
  assign n13771 = n13757 | n13770 ;
  assign n32528 = ~n13751 ;
  assign n13773 = n32528 & n13771 ;
  assign n13774 = n13750 | n13773 ;
  assign n13775 = n13542 | n13774 ;
  assign n32529 = ~n13540 ;
  assign n13776 = n32529 & n13775 ;
  assign n32530 = ~n13776 ;
  assign n13778 = n13473 & n32530 ;
  assign n32531 = ~n13778 ;
  assign n13779 = n13471 & n32531 ;
  assign n32532 = ~n13779 ;
  assign n13781 = n13400 & n32532 ;
  assign n32533 = ~n13781 ;
  assign n13782 = n13398 & n32533 ;
  assign n13783 = n13335 & n13782 ;
  assign n13784 = n13334 | n13783 ;
  assign n32534 = ~n13784 ;
  assign n13785 = n13299 & n32534 ;
  assign n32535 = ~n13785 ;
  assign n13786 = n13297 & n32535 ;
  assign n32536 = ~n13786 ;
  assign n13788 = n13246 & n32536 ;
  assign n32537 = ~n13788 ;
  assign n13789 = n13244 & n32537 ;
  assign n11702 = n11679 | n11701 ;
  assign n13790 = n11679 & n11701 ;
  assign n32538 = ~n13790 ;
  assign n13791 = n11702 & n32538 ;
  assign n32539 = ~n13791 ;
  assign n13792 = n13789 & n32539 ;
  assign n11538 = n895 & n11536 ;
  assign n10687 = n2849 & n10681 ;
  assign n10720 = n2861 & n10703 ;
  assign n13793 = n10687 | n10720 ;
  assign n13794 = n894 & n10679 ;
  assign n13795 = n13793 | n13794 ;
  assign n13796 = n11538 | n13795 ;
  assign n13797 = x29 | n13796 ;
  assign n13798 = x29 & n13796 ;
  assign n32540 = ~n13798 ;
  assign n13799 = n13797 & n32540 ;
  assign n32541 = ~n13789 ;
  assign n13800 = n32541 & n13791 ;
  assign n13801 = n13792 | n13800 ;
  assign n32542 = ~n13801 ;
  assign n13802 = n13799 & n32542 ;
  assign n13803 = n13792 | n13802 ;
  assign n13198 = n13177 | n13197 ;
  assign n32543 = ~n13199 ;
  assign n13804 = n13198 & n32543 ;
  assign n13806 = n13803 & n13804 ;
  assign n13807 = n13199 | n13806 ;
  assign n13808 = n13175 | n13807 ;
  assign n32544 = ~n13173 ;
  assign n13809 = n32544 & n13808 ;
  assign n13811 = n13149 | n13809 ;
  assign n32545 = ~n13147 ;
  assign n13812 = n32545 & n13811 ;
  assign n13814 = n13137 | n13812 ;
  assign n32546 = ~n13137 ;
  assign n13813 = n32546 & n13812 ;
  assign n32547 = ~n13812 ;
  assign n13815 = n13137 & n32547 ;
  assign n13816 = n13813 | n13815 ;
  assign n12618 = n12136 & n12617 ;
  assign n13817 = n12136 | n12622 ;
  assign n32548 = ~n12618 ;
  assign n13818 = n32548 & n13817 ;
  assign n32549 = ~n13818 ;
  assign n13819 = n12595 & n32549 ;
  assign n13820 = n32366 & n13818 ;
  assign n13821 = n13819 | n13820 ;
  assign n32550 = ~n13821 ;
  assign n13822 = n3791 & n32550 ;
  assign n12141 = n3802 & n32253 ;
  assign n12172 = n209 & n12161 ;
  assign n13833 = n12141 | n12172 ;
  assign n13834 = n3818 & n12595 ;
  assign n13835 = n13833 | n13834 ;
  assign n13836 = n13822 | n13835 ;
  assign n32551 = ~n13836 ;
  assign n13837 = x26 & n32551 ;
  assign n13838 = n30019 & n13836 ;
  assign n13839 = n13837 | n13838 ;
  assign n32552 = ~n13839 ;
  assign n13840 = n13816 & n32552 ;
  assign n32553 = ~n13840 ;
  assign n13841 = n13814 & n32553 ;
  assign n32554 = ~n13841 ;
  assign n13843 = n13135 & n32554 ;
  assign n13106 = n13077 & n13105 ;
  assign n32555 = ~n13077 ;
  assign n13844 = n32555 & n13101 ;
  assign n13845 = n13106 | n13844 ;
  assign n13846 = n32456 & n13845 ;
  assign n32556 = ~n13845 ;
  assign n13847 = n13052 & n32556 ;
  assign n13848 = n13846 | n13847 ;
  assign n32557 = ~n13848 ;
  assign n13849 = n4135 & n32557 ;
  assign n12554 = n4185 & n32354 ;
  assign n13083 = n4148 & n13077 ;
  assign n13860 = n12554 | n13083 ;
  assign n13861 = n4165 & n32456 ;
  assign n13862 = n13860 | n13861 ;
  assign n13863 = n13849 | n13862 ;
  assign n32558 = ~n13863 ;
  assign n13864 = x23 & n32558 ;
  assign n13865 = n30030 & n13863 ;
  assign n13866 = n13864 | n13865 ;
  assign n32559 = ~n13135 ;
  assign n13842 = n32559 & n13841 ;
  assign n13867 = n13842 | n13843 ;
  assign n13868 = n13866 | n13867 ;
  assign n32560 = ~n13843 ;
  assign n13869 = n32560 & n13868 ;
  assign n32561 = ~n13133 ;
  assign n13870 = n32561 & n13869 ;
  assign n32562 = ~n13869 ;
  assign n13871 = n13133 & n32562 ;
  assign n13872 = n13870 | n13871 ;
  assign n6452 = n3791 & n6445 ;
  assign n13873 = n3802 & n30545 ;
  assign n13874 = n209 & n30535 ;
  assign n13875 = n13873 | n13874 ;
  assign n13876 = n6452 | n13875 ;
  assign n13877 = x26 | n13876 ;
  assign n13878 = x26 & n13876 ;
  assign n32563 = ~n13878 ;
  assign n13879 = n13877 & n32563 ;
  assign n12976 = x23 & n32425 ;
  assign n13880 = n30030 & n12974 ;
  assign n13881 = n12976 | n13880 ;
  assign n13882 = n520 | n756 ;
  assign n13883 = n2584 | n13882 ;
  assign n13884 = n712 | n13883 ;
  assign n13885 = n1435 | n4943 ;
  assign n13886 = n2208 | n13885 ;
  assign n13887 = n190 | n405 ;
  assign n13888 = n538 | n13887 ;
  assign n13889 = n794 | n13888 ;
  assign n13890 = n13886 | n13889 ;
  assign n13891 = n13884 | n13890 ;
  assign n13892 = n214 | n220 ;
  assign n13893 = n239 | n13892 ;
  assign n13894 = n585 | n1346 ;
  assign n13895 = n13893 | n13894 ;
  assign n13896 = n1046 | n13895 ;
  assign n13897 = n11625 | n13896 ;
  assign n13898 = n224 | n400 ;
  assign n13899 = n996 | n13898 ;
  assign n13900 = n3055 | n13899 ;
  assign n13901 = n3260 | n13900 ;
  assign n13902 = n873 | n13901 ;
  assign n13903 = n13897 | n13902 ;
  assign n13904 = n13891 | n13903 ;
  assign n13905 = n13357 | n13904 ;
  assign n13906 = n13881 | n13905 ;
  assign n13907 = n13881 & n13905 ;
  assign n32564 = ~n13907 ;
  assign n13908 = n13906 & n32564 ;
  assign n13909 = n12838 & n12974 ;
  assign n13910 = n12981 | n13909 ;
  assign n13911 = n13908 | n13910 ;
  assign n13912 = n13908 & n13910 ;
  assign n32565 = ~n13912 ;
  assign n13913 = n13911 & n32565 ;
  assign n4840 = n889 & n30385 ;
  assign n4580 = n3311 & n30361 ;
  assign n4829 = n3343 & n4811 ;
  assign n13914 = n4580 | n4829 ;
  assign n13915 = n3329 & n4664 ;
  assign n13916 = n13914 | n13915 ;
  assign n13917 = n4840 | n13916 ;
  assign n32566 = ~n13917 ;
  assign n13918 = n13913 & n32566 ;
  assign n32567 = ~n13913 ;
  assign n13919 = n32567 & n13917 ;
  assign n13920 = n13918 | n13919 ;
  assign n32568 = ~n12950 ;
  assign n13921 = n32568 & n12989 ;
  assign n32569 = ~n13921 ;
  assign n13922 = n12987 & n32569 ;
  assign n13924 = n13920 | n13922 ;
  assign n13923 = n13920 & n13922 ;
  assign n32570 = ~n13923 ;
  assign n13925 = n32570 & n13924 ;
  assign n5141 = n895 & n30410 ;
  assign n4936 = n894 & n30415 ;
  assign n5116 = n2861 & n30405 ;
  assign n13926 = n4936 | n5116 ;
  assign n13927 = n2849 & n5017 ;
  assign n13928 = n13926 | n13927 ;
  assign n13929 = n5141 | n13928 ;
  assign n32571 = ~n13929 ;
  assign n13930 = x29 & n32571 ;
  assign n13931 = n30024 & n13929 ;
  assign n13932 = n13930 | n13931 ;
  assign n32572 = ~n13932 ;
  assign n13933 = n13925 & n32572 ;
  assign n32573 = ~n13933 ;
  assign n13934 = n13924 & n32573 ;
  assign n13935 = n13879 & n13934 ;
  assign n6419 = n895 & n6411 ;
  assign n4934 = n2849 & n30415 ;
  assign n5018 = n2861 & n5017 ;
  assign n13936 = n4934 | n5018 ;
  assign n13937 = n894 & n30530 ;
  assign n13938 = n13936 | n13937 ;
  assign n13939 = n6419 | n13938 ;
  assign n32574 = ~n13939 ;
  assign n13940 = x29 & n32574 ;
  assign n13941 = n30024 & n13939 ;
  assign n13942 = n13940 | n13941 ;
  assign n13943 = n13913 & n13917 ;
  assign n32575 = ~n13943 ;
  assign n13944 = n13911 & n32575 ;
  assign n32576 = ~n13881 ;
  assign n13945 = n32576 & n13905 ;
  assign n13946 = n13880 | n13945 ;
  assign n13947 = n318 | n476 ;
  assign n13948 = n528 | n554 ;
  assign n13949 = n13947 | n13948 ;
  assign n13950 = n708 | n13949 ;
  assign n13951 = n2070 | n13950 ;
  assign n13952 = n489 | n635 ;
  assign n13953 = n496 | n13952 ;
  assign n13954 = n2430 | n13953 ;
  assign n13955 = n2628 | n3888 ;
  assign n13956 = n13954 | n13955 ;
  assign n13957 = n4255 | n5830 ;
  assign n13958 = n13434 | n13957 ;
  assign n13959 = n507 | n1497 ;
  assign n13960 = n2243 | n3228 ;
  assign n13961 = n13959 | n13960 ;
  assign n13962 = n13958 | n13961 ;
  assign n13963 = n13956 | n13962 ;
  assign n13964 = n13951 | n13963 ;
  assign n13965 = n4293 | n13964 ;
  assign n13966 = n3546 | n13965 ;
  assign n13967 = n1400 | n13966 ;
  assign n32577 = ~n13967 ;
  assign n13968 = n13946 & n32577 ;
  assign n32578 = ~n13946 ;
  assign n13969 = n32578 & n13967 ;
  assign n13970 = n13968 | n13969 ;
  assign n6143 = n889 & n30578 ;
  assign n4826 = n3329 & n4811 ;
  assign n5117 = n3343 & n30405 ;
  assign n13971 = n4826 | n5117 ;
  assign n13972 = n3311 & n4664 ;
  assign n13973 = n13971 | n13972 ;
  assign n13974 = n6143 | n13973 ;
  assign n13975 = n13970 | n13974 ;
  assign n13977 = n13970 & n13974 ;
  assign n32579 = ~n13977 ;
  assign n13978 = n13975 & n32579 ;
  assign n13979 = n13944 & n13978 ;
  assign n13980 = n13944 | n13978 ;
  assign n32580 = ~n13979 ;
  assign n13981 = n32580 & n13980 ;
  assign n32581 = ~n13942 ;
  assign n13982 = n32581 & n13981 ;
  assign n32582 = ~n13981 ;
  assign n13983 = n13942 & n32582 ;
  assign n13984 = n13982 | n13983 ;
  assign n13985 = n13879 | n13934 ;
  assign n32583 = ~n13935 ;
  assign n13986 = n32583 & n13985 ;
  assign n13988 = n13984 & n13986 ;
  assign n13989 = n13935 | n13988 ;
  assign n6271 = n3791 & n30597 ;
  assign n13990 = n209 | n6271 ;
  assign n13991 = n30545 & n13990 ;
  assign n13992 = n30019 & n13991 ;
  assign n32584 = ~n13991 ;
  assign n13993 = x26 & n32584 ;
  assign n13994 = n13992 | n13993 ;
  assign n13995 = n248 | n270 ;
  assign n13996 = n622 | n13995 ;
  assign n13997 = n1161 | n2584 ;
  assign n13998 = n13996 | n13997 ;
  assign n13999 = n1463 | n2628 ;
  assign n14000 = n13625 | n13999 ;
  assign n14001 = n13998 | n14000 ;
  assign n14002 = n4079 | n14001 ;
  assign n14003 = n4273 | n13209 ;
  assign n14004 = n13476 | n14003 ;
  assign n14005 = n369 | n383 ;
  assign n14006 = n550 | n827 ;
  assign n14007 = n14005 | n14006 ;
  assign n14008 = n133 | n236 ;
  assign n14009 = n242 | n14008 ;
  assign n14010 = n14007 | n14009 ;
  assign n14011 = n382 | n1361 ;
  assign n14012 = n14010 | n14011 ;
  assign n14013 = n14004 | n14012 ;
  assign n14014 = n11229 | n14013 ;
  assign n14015 = n2192 | n5764 ;
  assign n14016 = n13254 | n14015 ;
  assign n14017 = n592 | n833 ;
  assign n14018 = n1422 | n1730 ;
  assign n14019 = n14017 | n14018 ;
  assign n14020 = n14016 | n14019 ;
  assign n14021 = n806 | n1381 ;
  assign n14022 = n14020 | n14021 ;
  assign n14023 = n13498 | n14022 ;
  assign n14024 = n14014 | n14023 ;
  assign n14025 = n14002 | n14024 ;
  assign n14026 = n32577 & n14025 ;
  assign n32585 = ~n14025 ;
  assign n14027 = n13967 & n32585 ;
  assign n14028 = n14026 | n14027 ;
  assign n5749 = n889 & n30512 ;
  assign n4830 = n3311 & n4811 ;
  assign n5118 = n3329 & n30405 ;
  assign n14029 = n4830 | n5118 ;
  assign n14030 = n3343 & n5017 ;
  assign n14031 = n14029 | n14030 ;
  assign n14032 = n5749 | n14031 ;
  assign n14033 = n14028 | n14032 ;
  assign n14035 = n14028 & n14032 ;
  assign n32586 = ~n14035 ;
  assign n14036 = n14033 & n32586 ;
  assign n13976 = n13968 | n13974 ;
  assign n32587 = ~n13969 ;
  assign n14037 = n32587 & n13976 ;
  assign n14038 = n14036 & n14037 ;
  assign n14039 = n14036 | n14037 ;
  assign n32588 = ~n14038 ;
  assign n14040 = n32588 & n14039 ;
  assign n14041 = n13979 | n13982 ;
  assign n14042 = n14040 | n14041 ;
  assign n14043 = n14040 & n14041 ;
  assign n32589 = ~n14043 ;
  assign n14044 = n14042 & n32589 ;
  assign n6170 = n895 & n30587 ;
  assign n4939 = n2861 & n30415 ;
  assign n5875 = n2849 & n30530 ;
  assign n14046 = n4939 | n5875 ;
  assign n14047 = n894 & n30535 ;
  assign n14048 = n14046 | n14047 ;
  assign n14049 = n6170 | n14048 ;
  assign n14050 = n14044 | n14049 ;
  assign n14052 = n14044 & n14049 ;
  assign n32590 = ~n14052 ;
  assign n14053 = n14050 & n32590 ;
  assign n14054 = n30024 & n14053 ;
  assign n32591 = ~n14053 ;
  assign n14055 = x29 & n32591 ;
  assign n14056 = n14054 | n14055 ;
  assign n14057 = n13994 | n14056 ;
  assign n14058 = n13994 & n14056 ;
  assign n32592 = ~n14058 ;
  assign n14059 = n14057 & n32592 ;
  assign n32593 = ~n13989 ;
  assign n14060 = n32593 & n14059 ;
  assign n32594 = ~n14059 ;
  assign n14061 = n13989 & n32594 ;
  assign n14062 = n14060 | n14061 ;
  assign n32595 = ~n13984 ;
  assign n13987 = n32595 & n13986 ;
  assign n32596 = ~n13986 ;
  assign n14063 = n13984 & n32596 ;
  assign n14064 = n13987 | n14063 ;
  assign n32597 = ~n13925 ;
  assign n14065 = n32597 & n13932 ;
  assign n14066 = n13933 | n14065 ;
  assign n5930 = n3791 & n30540 ;
  assign n5794 = n3818 & n30545 ;
  assign n5916 = n3802 & n30535 ;
  assign n14067 = n5794 | n5916 ;
  assign n14068 = n209 & n30530 ;
  assign n14069 = n14067 | n14068 ;
  assign n14070 = n5930 | n14069 ;
  assign n32598 = ~n14070 ;
  assign n14071 = x26 & n32598 ;
  assign n14072 = n30019 & n14070 ;
  assign n14073 = n14071 | n14072 ;
  assign n14074 = n14066 | n14073 ;
  assign n14075 = n14066 & n14073 ;
  assign n32599 = ~n14075 ;
  assign n14076 = n14074 & n32599 ;
  assign n14077 = n13000 | n13003 ;
  assign n32600 = ~n14077 ;
  assign n14078 = n14076 & n32600 ;
  assign n32601 = ~n14078 ;
  assign n14079 = n14074 & n32601 ;
  assign n14081 = n14064 | n14079 ;
  assign n14080 = n14064 & n14079 ;
  assign n32602 = ~n14080 ;
  assign n14082 = n32602 & n14081 ;
  assign n32603 = ~n14076 ;
  assign n14083 = n32603 & n14077 ;
  assign n14084 = n14078 | n14083 ;
  assign n32604 = ~n13017 ;
  assign n14085 = n13014 & n32604 ;
  assign n14087 = n14084 | n14085 ;
  assign n32605 = ~n14084 ;
  assign n14086 = n32605 & n14085 ;
  assign n32606 = ~n14085 ;
  assign n14088 = n14084 & n32606 ;
  assign n14089 = n14086 | n14088 ;
  assign n32607 = ~n13025 ;
  assign n14090 = n13023 & n32607 ;
  assign n32608 = ~n14090 ;
  assign n14092 = n14089 & n32608 ;
  assign n32609 = ~n14092 ;
  assign n14093 = n14087 & n32609 ;
  assign n32610 = ~n14093 ;
  assign n14096 = n14082 & n32610 ;
  assign n32611 = ~n14096 ;
  assign n14097 = n14081 & n32611 ;
  assign n14098 = n14062 | n14097 ;
  assign n14100 = n14062 & n14097 ;
  assign n32612 = ~n14100 ;
  assign n14101 = n14098 & n32612 ;
  assign n14094 = n14082 & n14093 ;
  assign n14123 = n14082 | n14093 ;
  assign n32613 = ~n14094 ;
  assign n14124 = n32613 & n14123 ;
  assign n14091 = n14089 & n14090 ;
  assign n14146 = n14089 | n14090 ;
  assign n32614 = ~n14091 ;
  assign n14147 = n32614 & n14146 ;
  assign n32615 = ~n13107 ;
  assign n14175 = n13052 & n32615 ;
  assign n32616 = ~n14175 ;
  assign n14176 = n13027 & n32616 ;
  assign n14177 = n14147 | n14176 ;
  assign n32617 = ~n14177 ;
  assign n14178 = n14124 & n32617 ;
  assign n14170 = n32456 & n13102 ;
  assign n14172 = n13027 | n14170 ;
  assign n14174 = n14147 & n14172 ;
  assign n32618 = ~n14124 ;
  assign n14179 = n32618 & n14174 ;
  assign n14180 = n14178 | n14179 ;
  assign n14181 = n14101 & n14180 ;
  assign n14182 = n14101 | n14180 ;
  assign n32619 = ~n14181 ;
  assign n14183 = n32619 & n14182 ;
  assign n14184 = n4686 & n14183 ;
  assign n14126 = n4706 & n14124 ;
  assign n14160 = n4726 & n14147 ;
  assign n14197 = n14126 | n14160 ;
  assign n32620 = ~n14097 ;
  assign n14099 = n14062 & n32620 ;
  assign n32621 = ~n14062 ;
  assign n14195 = n32621 & n14097 ;
  assign n14196 = n14099 | n14195 ;
  assign n14198 = n4748 & n14196 ;
  assign n14199 = n14197 | n14198 ;
  assign n14200 = n14184 | n14199 ;
  assign n32622 = ~n14200 ;
  assign n14201 = x20 & n32622 ;
  assign n14202 = n30374 & n14200 ;
  assign n14203 = n14201 | n14202 ;
  assign n32623 = ~n14203 ;
  assign n14204 = n13872 & n32623 ;
  assign n32624 = ~n13872 ;
  assign n14205 = n32624 & n14203 ;
  assign n14206 = n14204 | n14205 ;
  assign n14207 = n13866 & n13867 ;
  assign n32625 = ~n14207 ;
  assign n14208 = n13868 & n32625 ;
  assign n32626 = ~n13816 ;
  assign n14209 = n32626 & n13839 ;
  assign n14210 = n13840 | n14209 ;
  assign n32627 = ~n13149 ;
  assign n13810 = n32627 & n13809 ;
  assign n32628 = ~n13809 ;
  assign n14211 = n13149 & n32628 ;
  assign n14212 = n13810 | n14211 ;
  assign n14213 = n13175 & n13807 ;
  assign n32629 = ~n14213 ;
  assign n14214 = n13808 & n32629 ;
  assign n11514 = n895 & n11511 ;
  assign n10659 = n2849 & n10656 ;
  assign n11045 = n2861 & n10679 ;
  assign n14215 = n10659 | n11045 ;
  assign n14216 = n894 & n11452 ;
  assign n14217 = n14215 | n14216 ;
  assign n14218 = n11514 | n14217 ;
  assign n14219 = x29 | n14218 ;
  assign n14220 = x29 & n14218 ;
  assign n32630 = ~n14220 ;
  assign n14221 = n14219 & n32630 ;
  assign n32631 = ~n14221 ;
  assign n14223 = n14214 & n32631 ;
  assign n12656 = n3791 & n32362 ;
  assign n11444 = n209 & n11430 ;
  assign n11845 = n3802 & n32176 ;
  assign n14224 = n11444 | n11845 ;
  assign n14225 = n3818 & n12161 ;
  assign n14226 = n14224 | n14225 ;
  assign n14227 = n12656 | n14226 ;
  assign n32632 = ~n14227 ;
  assign n14228 = x26 & n32632 ;
  assign n14229 = n30019 & n14227 ;
  assign n14230 = n14228 | n14229 ;
  assign n14222 = n14214 & n14221 ;
  assign n14231 = n14214 | n14221 ;
  assign n32633 = ~n14222 ;
  assign n14232 = n32633 & n14231 ;
  assign n14233 = n14230 | n14232 ;
  assign n32634 = ~n14223 ;
  assign n14234 = n32634 & n14233 ;
  assign n32635 = ~n14234 ;
  assign n14236 = n14212 & n32635 ;
  assign n14235 = n14212 & n14234 ;
  assign n14237 = n14212 | n14234 ;
  assign n32636 = ~n14235 ;
  assign n14238 = n32636 & n14237 ;
  assign n12195 = n3791 & n32255 ;
  assign n11853 = n209 & n32176 ;
  assign n12171 = n3802 & n12161 ;
  assign n14239 = n11853 | n12171 ;
  assign n14240 = n3818 & n32253 ;
  assign n14241 = n14239 | n14240 ;
  assign n14242 = n12195 | n14241 ;
  assign n32637 = ~n14242 ;
  assign n14243 = x26 & n32637 ;
  assign n14244 = n30019 & n14242 ;
  assign n14245 = n14243 | n14244 ;
  assign n14246 = n14238 | n14245 ;
  assign n32638 = ~n14236 ;
  assign n14247 = n32638 & n14246 ;
  assign n14249 = n14210 | n14247 ;
  assign n13100 = n12544 | n13099 ;
  assign n14250 = n12544 & n13104 ;
  assign n32639 = ~n14250 ;
  assign n14251 = n13100 & n32639 ;
  assign n32640 = ~n14251 ;
  assign n14252 = n13077 & n32640 ;
  assign n14253 = n32555 & n14251 ;
  assign n14254 = n14252 | n14253 ;
  assign n32641 = ~n14254 ;
  assign n14256 = n4135 & n32641 ;
  assign n12550 = n4148 & n32354 ;
  assign n12580 = n4185 & n12570 ;
  assign n14266 = n12550 | n12580 ;
  assign n14267 = n4165 & n13077 ;
  assign n14268 = n14266 | n14267 ;
  assign n14269 = n14256 | n14268 ;
  assign n32642 = ~n14269 ;
  assign n14270 = x23 & n32642 ;
  assign n14271 = n30030 & n14269 ;
  assign n14272 = n14270 | n14271 ;
  assign n32643 = ~n14210 ;
  assign n14248 = n32643 & n14247 ;
  assign n32644 = ~n14247 ;
  assign n14273 = n14210 & n32644 ;
  assign n14274 = n14248 | n14273 ;
  assign n32645 = ~n14272 ;
  assign n14275 = n32645 & n14274 ;
  assign n32646 = ~n14275 ;
  assign n14276 = n14249 & n32646 ;
  assign n32647 = ~n14208 ;
  assign n14278 = n32647 & n14276 ;
  assign n32648 = ~n14172 ;
  assign n14173 = n14147 & n32648 ;
  assign n32649 = ~n14147 ;
  assign n14279 = n32649 & n14176 ;
  assign n14280 = n14173 | n14279 ;
  assign n14281 = n14124 & n14280 ;
  assign n14282 = n14124 | n14280 ;
  assign n32650 = ~n14281 ;
  assign n14283 = n32650 & n14282 ;
  assign n14284 = n4686 & n14283 ;
  assign n13043 = n4726 & n13027 ;
  assign n14158 = n4706 & n14147 ;
  assign n14296 = n13043 | n14158 ;
  assign n32651 = ~n14082 ;
  assign n14095 = n32651 & n14093 ;
  assign n14295 = n14095 | n14096 ;
  assign n14297 = n4748 & n14295 ;
  assign n14298 = n14296 | n14297 ;
  assign n14299 = n14284 | n14298 ;
  assign n32652 = ~n14299 ;
  assign n14300 = x20 & n32652 ;
  assign n14301 = n30374 & n14299 ;
  assign n14302 = n14300 | n14301 ;
  assign n14277 = n14208 & n14276 ;
  assign n14303 = n14208 | n14276 ;
  assign n32653 = ~n14277 ;
  assign n14304 = n32653 & n14303 ;
  assign n32654 = ~n14304 ;
  assign n14306 = n14302 & n32654 ;
  assign n14307 = n14278 | n14306 ;
  assign n14308 = n14206 | n14307 ;
  assign n14309 = n14206 & n14307 ;
  assign n32655 = ~n14309 ;
  assign n14310 = n14308 & n32655 ;
  assign n14311 = x26 & n30007 ;
  assign n14312 = n30545 & n14311 ;
  assign n14313 = x29 | n14312 ;
  assign n14314 = n376 | n707 ;
  assign n14315 = n13679 | n14314 ;
  assign n14316 = n279 | n289 ;
  assign n14317 = n508 | n610 ;
  assign n14318 = n14316 | n14317 ;
  assign n14319 = n868 | n1860 ;
  assign n14320 = n14318 | n14319 ;
  assign n14321 = n235 | n591 ;
  assign n14322 = n239 | n14321 ;
  assign n14323 = n1541 | n2985 ;
  assign n14324 = n14322 | n14323 ;
  assign n14325 = n14320 | n14324 ;
  assign n14326 = n2490 | n3031 ;
  assign n14327 = n3967 | n4857 ;
  assign n14328 = n14326 | n14327 ;
  assign n14329 = n249 | n509 ;
  assign n14330 = n2325 | n14329 ;
  assign n14331 = n1126 | n14330 ;
  assign n14332 = n14328 | n14331 ;
  assign n14333 = n1043 | n1637 ;
  assign n14334 = n14332 | n14333 ;
  assign n14335 = n1841 | n2407 ;
  assign n14336 = n2920 | n3729 ;
  assign n14337 = n14335 | n14336 ;
  assign n14338 = n3059 | n14337 ;
  assign n14339 = n14334 | n14338 ;
  assign n14340 = n14325 | n14339 ;
  assign n14341 = n14315 | n14340 ;
  assign n32656 = ~n14341 ;
  assign n14342 = n940 & n32656 ;
  assign n14343 = n1729 | n2478 ;
  assign n14344 = n3537 | n14343 ;
  assign n14345 = n4985 | n14344 ;
  assign n14346 = n5606 | n14345 ;
  assign n14347 = n380 | n497 ;
  assign n14348 = n1199 | n14347 ;
  assign n14349 = n216 | n313 ;
  assign n14350 = n621 | n14349 ;
  assign n14351 = n14348 | n14350 ;
  assign n14352 = n1123 | n4009 ;
  assign n14353 = n14351 | n14352 ;
  assign n14354 = n13269 | n14353 ;
  assign n14355 = n14346 | n14354 ;
  assign n32657 = ~n13669 ;
  assign n14356 = n4532 & n32657 ;
  assign n32658 = ~n14355 ;
  assign n14357 = n32658 & n14356 ;
  assign n32659 = ~n11926 ;
  assign n14358 = n32659 & n14357 ;
  assign n14359 = n14342 & n14358 ;
  assign n14360 = n14342 | n14358 ;
  assign n32660 = ~n14359 ;
  assign n14361 = n32660 & n14360 ;
  assign n14362 = n529 | n532 ;
  assign n14363 = n636 | n839 ;
  assign n14364 = n14362 | n14363 ;
  assign n14365 = n623 | n14364 ;
  assign n14366 = n1853 | n11233 ;
  assign n14367 = n14365 | n14366 ;
  assign n14368 = n13337 | n14367 ;
  assign n14369 = n1826 | n3436 ;
  assign n14370 = n3493 | n13553 ;
  assign n14371 = n14369 | n14370 ;
  assign n14372 = n634 | n858 ;
  assign n14373 = n1101 | n2364 ;
  assign n14374 = n14372 | n14373 ;
  assign n14375 = n353 | n400 ;
  assign n14376 = n344 | n14375 ;
  assign n14377 = n784 | n14376 ;
  assign n14378 = n14374 | n14377 ;
  assign n14379 = n4334 | n14378 ;
  assign n14380 = n14371 | n14379 ;
  assign n14381 = n14368 | n14380 ;
  assign n14382 = n308 | n14381 ;
  assign n14383 = n2508 | n14382 ;
  assign n14385 = n13967 & n14383 ;
  assign n14384 = n13967 | n14383 ;
  assign n32661 = ~n14385 ;
  assign n14386 = n14384 & n32661 ;
  assign n14387 = n30019 & n14386 ;
  assign n14388 = n14385 | n14387 ;
  assign n14389 = n14358 | n14388 ;
  assign n14390 = n14358 & n14388 ;
  assign n6413 = n889 & n6411 ;
  assign n4941 = n3329 & n30415 ;
  assign n5019 = n3311 & n5017 ;
  assign n14391 = n4941 | n5019 ;
  assign n14392 = n3343 & n30530 ;
  assign n14393 = n14391 | n14392 ;
  assign n14394 = n6413 | n14393 ;
  assign n14395 = n14390 | n14394 ;
  assign n14396 = n14389 & n14395 ;
  assign n14397 = n14361 & n14396 ;
  assign n14398 = n14361 | n14396 ;
  assign n32662 = ~n14397 ;
  assign n14399 = n32662 & n14398 ;
  assign n6168 = n889 & n30587 ;
  assign n14402 = n3326 & n30530 ;
  assign n85 = x31 | n84 ;
  assign n14400 = n85 & n5870 ;
  assign n14401 = n81 | n14400 ;
  assign n14403 = n30676 & n14401 ;
  assign n14404 = n14402 | n14403 ;
  assign n14405 = n6168 | n14404 ;
  assign n32663 = ~n14405 ;
  assign n14406 = n14399 & n32663 ;
  assign n32664 = ~n14399 ;
  assign n14407 = n32664 & n14405 ;
  assign n14408 = n14406 | n14407 ;
  assign n14409 = n14313 | n14408 ;
  assign n14410 = n14313 & n14408 ;
  assign n32665 = ~n14410 ;
  assign n14411 = n14409 & n32665 ;
  assign n32666 = ~n14390 ;
  assign n14412 = n14389 & n32666 ;
  assign n32667 = ~n14394 ;
  assign n14413 = n32667 & n14412 ;
  assign n32668 = ~n14412 ;
  assign n14414 = n14394 & n32668 ;
  assign n14415 = n14413 | n14414 ;
  assign n32669 = ~n14386 ;
  assign n14416 = x26 & n32669 ;
  assign n14417 = n14387 | n14416 ;
  assign n14034 = n14026 | n14032 ;
  assign n32670 = ~n14027 ;
  assign n14418 = n32670 & n14034 ;
  assign n32671 = ~n14418 ;
  assign n14420 = n14417 & n32671 ;
  assign n32672 = ~n14417 ;
  assign n14419 = n32672 & n14418 ;
  assign n5142 = n889 & n30410 ;
  assign n4942 = n3343 & n30415 ;
  assign n5119 = n3311 & n30405 ;
  assign n14421 = n4942 | n5119 ;
  assign n14422 = n3329 & n5017 ;
  assign n14423 = n14421 | n14422 ;
  assign n14424 = n5142 | n14423 ;
  assign n14425 = n14419 | n14424 ;
  assign n32673 = ~n14420 ;
  assign n14426 = n32673 & n14425 ;
  assign n14428 = n14415 & n14426 ;
  assign n6453 = n895 & n6445 ;
  assign n14429 = n2849 & n30545 ;
  assign n14430 = n2861 & n30535 ;
  assign n14431 = n14429 | n14430 ;
  assign n14432 = n6453 | n14431 ;
  assign n32674 = ~n14432 ;
  assign n14433 = x29 & n32674 ;
  assign n14434 = n30024 & n14432 ;
  assign n14435 = n14433 | n14434 ;
  assign n32675 = ~n14415 ;
  assign n14427 = n32675 & n14426 ;
  assign n32676 = ~n14426 ;
  assign n14436 = n14415 & n32676 ;
  assign n14437 = n14427 | n14436 ;
  assign n14439 = n14435 & n14437 ;
  assign n14440 = n14428 | n14439 ;
  assign n32677 = ~n14440 ;
  assign n14441 = n14411 & n32677 ;
  assign n32678 = ~n14411 ;
  assign n14442 = n32678 & n14440 ;
  assign n14443 = n14441 | n14442 ;
  assign n32679 = ~n14435 ;
  assign n14438 = n32679 & n14437 ;
  assign n32680 = ~n14437 ;
  assign n14444 = n14435 & n32680 ;
  assign n14445 = n14438 | n14444 ;
  assign n5926 = n895 & n30540 ;
  assign n32681 = ~n2861 ;
  assign n5799 = n32681 & n5793 ;
  assign n14446 = n894 | n5793 ;
  assign n32682 = ~n5799 ;
  assign n14447 = n32682 & n14446 ;
  assign n14448 = n2849 & n30535 ;
  assign n14449 = n14447 | n14448 ;
  assign n14450 = n5926 | n14449 ;
  assign n32683 = ~n14450 ;
  assign n14451 = x29 & n32683 ;
  assign n14452 = n30024 & n14450 ;
  assign n14453 = n14451 | n14452 ;
  assign n32684 = ~n14037 ;
  assign n14454 = n14036 & n32684 ;
  assign n32685 = ~n14040 ;
  assign n14455 = n32685 & n14041 ;
  assign n14456 = n14454 | n14455 ;
  assign n32686 = ~n14453 ;
  assign n14458 = n32686 & n14456 ;
  assign n14457 = n14453 | n14456 ;
  assign n14459 = n14453 & n14456 ;
  assign n32687 = ~n14459 ;
  assign n14460 = n14457 & n32687 ;
  assign n14461 = n14419 | n14420 ;
  assign n14462 = n14424 | n14461 ;
  assign n14463 = n14424 & n14461 ;
  assign n32688 = ~n14463 ;
  assign n14464 = n14462 & n32688 ;
  assign n32689 = ~n14460 ;
  assign n14465 = n32689 & n14464 ;
  assign n14466 = n14458 | n14465 ;
  assign n32690 = ~n14445 ;
  assign n14468 = n32690 & n14466 ;
  assign n32691 = ~n14466 ;
  assign n14467 = n14445 & n32691 ;
  assign n14469 = n14467 | n14468 ;
  assign n32692 = ~n14464 ;
  assign n14470 = n14460 & n32692 ;
  assign n14471 = n14465 | n14470 ;
  assign n14045 = n13994 | n14044 ;
  assign n14472 = n13994 & n14044 ;
  assign n32693 = ~n14049 ;
  assign n14051 = x29 & n32693 ;
  assign n14473 = n30024 & n14049 ;
  assign n14474 = n14051 | n14473 ;
  assign n14475 = n14472 | n14474 ;
  assign n14476 = n14045 & n14475 ;
  assign n14478 = n14471 | n14476 ;
  assign n32694 = ~n14471 ;
  assign n14477 = n32694 & n14476 ;
  assign n32695 = ~n14476 ;
  assign n14479 = n14471 & n32695 ;
  assign n14480 = n14477 | n14479 ;
  assign n14481 = n13989 | n14059 ;
  assign n32696 = ~n14099 ;
  assign n14482 = n32696 & n14481 ;
  assign n32697 = ~n14482 ;
  assign n14483 = n14480 & n32697 ;
  assign n32698 = ~n14483 ;
  assign n14484 = n14478 & n32698 ;
  assign n14486 = n14469 | n14484 ;
  assign n32699 = ~n14468 ;
  assign n14487 = n32699 & n14486 ;
  assign n14488 = n14443 | n14487 ;
  assign n14489 = n14443 & n14487 ;
  assign n32700 = ~n14489 ;
  assign n14490 = n14488 & n32700 ;
  assign n32701 = ~n14469 ;
  assign n14485 = n32701 & n14484 ;
  assign n32702 = ~n14484 ;
  assign n14512 = n14469 & n32702 ;
  assign n14513 = n14485 | n14512 ;
  assign n32703 = ~n14480 ;
  assign n14535 = n32703 & n14482 ;
  assign n14536 = n14483 | n14535 ;
  assign n14561 = n14124 & n14177 ;
  assign n14562 = n14196 | n14561 ;
  assign n14564 = n14536 & n14562 ;
  assign n14565 = n14513 & n14564 ;
  assign n14558 = n14124 | n14174 ;
  assign n14559 = n14101 & n14558 ;
  assign n14560 = n14536 | n14559 ;
  assign n14566 = n14513 | n14560 ;
  assign n32704 = ~n14565 ;
  assign n14567 = n32704 & n14566 ;
  assign n14568 = n14490 | n14567 ;
  assign n14569 = n14490 & n14567 ;
  assign n32705 = ~n14569 ;
  assign n14570 = n14568 & n32705 ;
  assign n14571 = n37300 & n14570 ;
  assign n32706 = ~n14513 ;
  assign n14527 = n5144 & n32706 ;
  assign n14544 = n5166 & n14536 ;
  assign n14582 = n14527 | n14544 ;
  assign n32707 = ~n14490 ;
  assign n14583 = n5191 & n32707 ;
  assign n14584 = n14582 | n14583 ;
  assign n14585 = n14571 | n14584 ;
  assign n32708 = ~n14585 ;
  assign n14586 = x17 & n32708 ;
  assign n14587 = n30580 & n14585 ;
  assign n14588 = n14586 | n14587 ;
  assign n14589 = n14310 | n14588 ;
  assign n14590 = n14310 & n14588 ;
  assign n32709 = ~n14590 ;
  assign n14591 = n14589 & n32709 ;
  assign n14305 = n14302 | n14304 ;
  assign n14592 = n14302 & n14304 ;
  assign n32710 = ~n14592 ;
  assign n14593 = n14305 & n32710 ;
  assign n32711 = ~n14274 ;
  assign n14594 = n14272 & n32711 ;
  assign n14595 = n14275 | n14594 ;
  assign n12632 = n4135 & n32356 ;
  assign n12576 = n4148 & n12570 ;
  assign n12604 = n4185 & n12595 ;
  assign n14596 = n12576 | n12604 ;
  assign n14597 = n4165 & n32354 ;
  assign n14598 = n14596 | n14597 ;
  assign n14599 = n12632 | n14598 ;
  assign n32712 = ~n14599 ;
  assign n14600 = x23 & n32712 ;
  assign n14601 = n30030 & n14599 ;
  assign n14602 = n14600 | n14601 ;
  assign n12684 = n4135 & n12681 ;
  assign n12147 = n4185 & n32253 ;
  assign n12603 = n4148 & n12595 ;
  assign n14603 = n12147 | n12603 ;
  assign n14604 = n4165 & n12570 ;
  assign n14605 = n14603 | n14604 ;
  assign n14606 = n12684 | n14605 ;
  assign n14607 = x23 | n14606 ;
  assign n14608 = x23 & n14606 ;
  assign n32713 = ~n14608 ;
  assign n14609 = n14607 & n32713 ;
  assign n11033 = n895 & n11030 ;
  assign n10688 = n2861 & n10681 ;
  assign n11051 = n2849 & n10679 ;
  assign n14610 = n10688 | n11051 ;
  assign n14611 = n894 & n10656 ;
  assign n14612 = n14610 | n14611 ;
  assign n14613 = n11033 | n14612 ;
  assign n14614 = x29 | n14613 ;
  assign n14615 = x29 & n14613 ;
  assign n32714 = ~n14615 ;
  assign n14616 = n14614 & n32714 ;
  assign n11872 = n3791 & n32178 ;
  assign n11441 = n3802 & n11430 ;
  assign n11482 = n209 & n11476 ;
  assign n14617 = n11441 | n11482 ;
  assign n14618 = n3818 & n32176 ;
  assign n14619 = n14617 | n14618 ;
  assign n14620 = n11872 | n14619 ;
  assign n32715 = ~n14620 ;
  assign n14621 = x26 & n32715 ;
  assign n14622 = n30019 & n14620 ;
  assign n14623 = n14621 | n14622 ;
  assign n14625 = n14616 & n14623 ;
  assign n32716 = ~n13803 ;
  assign n13805 = n32716 & n13804 ;
  assign n32717 = ~n13804 ;
  assign n14626 = n13803 & n32717 ;
  assign n14627 = n13805 | n14626 ;
  assign n32718 = ~n14623 ;
  assign n14624 = n14616 & n32718 ;
  assign n32719 = ~n14616 ;
  assign n14628 = n32719 & n14623 ;
  assign n14629 = n14624 | n14628 ;
  assign n14630 = n14627 & n14629 ;
  assign n14631 = n14625 | n14630 ;
  assign n14633 = n14609 & n14631 ;
  assign n14634 = n14230 & n14232 ;
  assign n32720 = ~n14634 ;
  assign n14635 = n14233 & n32720 ;
  assign n32721 = ~n14631 ;
  assign n14632 = n14609 & n32721 ;
  assign n32722 = ~n14609 ;
  assign n14636 = n32722 & n14631 ;
  assign n14637 = n14632 | n14636 ;
  assign n32723 = ~n14635 ;
  assign n14638 = n32723 & n14637 ;
  assign n14639 = n14633 | n14638 ;
  assign n14641 = n14602 & n14639 ;
  assign n14642 = n14238 & n14245 ;
  assign n32724 = ~n14642 ;
  assign n14643 = n14246 & n32724 ;
  assign n14640 = n14602 | n14639 ;
  assign n32725 = ~n14641 ;
  assign n14644 = n14640 & n32725 ;
  assign n32726 = ~n14643 ;
  assign n14646 = n32726 & n14644 ;
  assign n14647 = n14641 | n14646 ;
  assign n14648 = n14595 | n14647 ;
  assign n14649 = n14595 & n14647 ;
  assign n32727 = ~n14649 ;
  assign n14650 = n14648 & n32727 ;
  assign n14171 = n32454 & n14170 ;
  assign n14651 = n13027 & n14175 ;
  assign n14652 = n14171 | n14651 ;
  assign n14653 = n14147 & n14652 ;
  assign n14654 = n14147 | n14652 ;
  assign n32728 = ~n14653 ;
  assign n14655 = n32728 & n14654 ;
  assign n14656 = n4686 & n14655 ;
  assign n13041 = n4706 & n13027 ;
  assign n13060 = n4726 & n32456 ;
  assign n14667 = n13041 | n13060 ;
  assign n14668 = n4748 & n14147 ;
  assign n14669 = n14667 | n14668 ;
  assign n14670 = n14656 | n14669 ;
  assign n32729 = ~n14670 ;
  assign n14671 = x20 & n32729 ;
  assign n14672 = n30374 & n14670 ;
  assign n14673 = n14671 | n14672 ;
  assign n32730 = ~n14673 ;
  assign n14674 = n14650 & n32730 ;
  assign n32731 = ~n14674 ;
  assign n14675 = n14648 & n32731 ;
  assign n32732 = ~n14675 ;
  assign n14677 = n14593 & n32732 ;
  assign n32733 = ~n14564 ;
  assign n14678 = n14560 & n32733 ;
  assign n14679 = n32706 & n14678 ;
  assign n32734 = ~n14678 ;
  assign n14680 = n14513 & n32734 ;
  assign n14681 = n14679 | n14680 ;
  assign n32735 = ~n14681 ;
  assign n14682 = n37300 & n32735 ;
  assign n14112 = n5166 & n14101 ;
  assign n14551 = n5144 & n14536 ;
  assign n14693 = n14112 | n14551 ;
  assign n14694 = n5191 & n32706 ;
  assign n14695 = n14693 | n14694 ;
  assign n14696 = n14682 | n14695 ;
  assign n14697 = x17 | n14696 ;
  assign n14698 = x17 & n14696 ;
  assign n32736 = ~n14698 ;
  assign n14699 = n14697 & n32736 ;
  assign n32737 = ~n14593 ;
  assign n14676 = n32737 & n14675 ;
  assign n14700 = n14676 | n14677 ;
  assign n14702 = n14699 | n14700 ;
  assign n32738 = ~n14677 ;
  assign n14703 = n32738 & n14702 ;
  assign n32739 = ~n14591 ;
  assign n14704 = n32739 & n14703 ;
  assign n32740 = ~n14703 ;
  assign n14705 = n14591 & n32740 ;
  assign n14706 = n14704 | n14705 ;
  assign n32741 = ~n14700 ;
  assign n14701 = n14699 & n32741 ;
  assign n32742 = ~n14699 ;
  assign n14707 = n32742 & n14700 ;
  assign n14708 = n14701 | n14707 ;
  assign n32743 = ~n14650 ;
  assign n14709 = n32743 & n14673 ;
  assign n14710 = n14674 | n14709 ;
  assign n14645 = n14643 & n14644 ;
  assign n14711 = n14643 | n14644 ;
  assign n32744 = ~n14645 ;
  assign n14712 = n32744 & n14711 ;
  assign n32745 = ~n14637 ;
  assign n14713 = n14635 & n32745 ;
  assign n14714 = n14638 | n14713 ;
  assign n14715 = n14627 | n14629 ;
  assign n32746 = ~n14630 ;
  assign n14716 = n32746 & n14715 ;
  assign n13825 = n4135 & n32550 ;
  assign n12145 = n4148 & n32253 ;
  assign n12169 = n4185 & n12161 ;
  assign n14717 = n12145 | n12169 ;
  assign n14718 = n4165 & n12595 ;
  assign n14719 = n14717 | n14718 ;
  assign n14720 = n13825 | n14719 ;
  assign n14721 = x23 | n14720 ;
  assign n14722 = x23 & n14720 ;
  assign n32747 = ~n14722 ;
  assign n14723 = n14721 & n32747 ;
  assign n14725 = n14716 | n14723 ;
  assign n32748 = ~n14716 ;
  assign n14724 = n32748 & n14723 ;
  assign n32749 = ~n14723 ;
  assign n14726 = n14716 & n32749 ;
  assign n14727 = n14724 | n14726 ;
  assign n32750 = ~n13799 ;
  assign n14728 = n32750 & n13801 ;
  assign n14729 = n13802 | n14728 ;
  assign n11468 = n3791 & n11463 ;
  assign n10658 = n209 & n10656 ;
  assign n11486 = n3802 & n11476 ;
  assign n14730 = n10658 | n11486 ;
  assign n14731 = n3818 & n11430 ;
  assign n14732 = n14730 | n14731 ;
  assign n14733 = n11468 | n14732 ;
  assign n14734 = x26 | n14733 ;
  assign n14735 = x26 & n14733 ;
  assign n32751 = ~n14735 ;
  assign n14736 = n14734 & n32751 ;
  assign n32752 = ~n14729 ;
  assign n14737 = n32752 & n14736 ;
  assign n13787 = n13246 & n13786 ;
  assign n14738 = n13246 | n13786 ;
  assign n32753 = ~n13787 ;
  assign n14739 = n32753 & n14738 ;
  assign n13159 = n895 & n13157 ;
  assign n10721 = n2849 & n10703 ;
  assign n10735 = n2861 & n10727 ;
  assign n14740 = n10721 | n10735 ;
  assign n14741 = n894 & n10681 ;
  assign n14742 = n14740 | n14741 ;
  assign n14743 = n13159 | n14742 ;
  assign n14744 = x29 | n14743 ;
  assign n14745 = x29 & n14743 ;
  assign n32754 = ~n14745 ;
  assign n14746 = n14744 & n32754 ;
  assign n14748 = n14739 | n14746 ;
  assign n32755 = ~n14739 ;
  assign n14747 = n32755 & n14746 ;
  assign n32756 = ~n14746 ;
  assign n14749 = n14739 & n32756 ;
  assign n14750 = n14747 | n14749 ;
  assign n32757 = ~n13299 ;
  assign n14751 = n32757 & n13784 ;
  assign n14752 = n13785 | n14751 ;
  assign n13185 = n895 & n13182 ;
  assign n10734 = n2849 & n10727 ;
  assign n10763 = n2861 & n31999 ;
  assign n14753 = n10734 | n10763 ;
  assign n14754 = n894 & n13151 ;
  assign n14755 = n14753 | n14754 ;
  assign n14756 = n13185 | n14755 ;
  assign n14757 = x29 | n14756 ;
  assign n14758 = x29 & n14756 ;
  assign n32758 = ~n14758 ;
  assign n14759 = n14757 & n32758 ;
  assign n14761 = n14752 | n14759 ;
  assign n32759 = ~n14752 ;
  assign n14760 = n32759 & n14759 ;
  assign n32760 = ~n14759 ;
  assign n14762 = n14752 & n32760 ;
  assign n14763 = n14760 | n14762 ;
  assign n14764 = n13335 | n13782 ;
  assign n32761 = ~n13783 ;
  assign n14765 = n32761 & n14764 ;
  assign n11688 = n895 & n32125 ;
  assign n10756 = n2849 & n31999 ;
  assign n10779 = n2861 & n10773 ;
  assign n14766 = n10756 | n10779 ;
  assign n14767 = n894 & n10727 ;
  assign n14768 = n14766 | n14767 ;
  assign n14769 = n11688 | n14768 ;
  assign n14770 = x29 | n14769 ;
  assign n14771 = x29 & n14769 ;
  assign n32762 = ~n14771 ;
  assign n14772 = n14770 & n32762 ;
  assign n14774 = n14765 | n14772 ;
  assign n13780 = n13400 & n13779 ;
  assign n14775 = n13400 | n13779 ;
  assign n32763 = ~n13780 ;
  assign n14776 = n32763 & n14775 ;
  assign n13230 = n895 & n32477 ;
  assign n10778 = n2849 & n10773 ;
  assign n10808 = n2861 & n31998 ;
  assign n14777 = n10778 | n10808 ;
  assign n14778 = n894 & n32478 ;
  assign n14779 = n14777 | n14778 ;
  assign n14780 = n13230 | n14779 ;
  assign n14781 = x29 | n14780 ;
  assign n14782 = x29 & n14780 ;
  assign n32764 = ~n14782 ;
  assign n14783 = n14781 & n32764 ;
  assign n14785 = n14776 | n14783 ;
  assign n32765 = ~n14776 ;
  assign n14784 = n32765 & n14783 ;
  assign n32766 = ~n14783 ;
  assign n14786 = n14776 & n32766 ;
  assign n14787 = n14784 | n14786 ;
  assign n13777 = n13473 & n13776 ;
  assign n14788 = n13473 | n13776 ;
  assign n32767 = ~n13777 ;
  assign n14789 = n32767 & n14788 ;
  assign n13281 = n895 & n32482 ;
  assign n10805 = n2849 & n31998 ;
  assign n10824 = n2861 & n10818 ;
  assign n14790 = n10805 | n10824 ;
  assign n14791 = n894 & n13292 ;
  assign n14792 = n14790 | n14791 ;
  assign n14793 = n13281 | n14792 ;
  assign n14794 = x29 | n14793 ;
  assign n14795 = x29 & n14793 ;
  assign n32768 = ~n14795 ;
  assign n14796 = n14794 & n32768 ;
  assign n14798 = n14789 | n14796 ;
  assign n32769 = ~n14789 ;
  assign n14797 = n32769 & n14796 ;
  assign n32770 = ~n14796 ;
  assign n14799 = n14789 & n32770 ;
  assign n14800 = n14797 | n14799 ;
  assign n14801 = n13542 & n13774 ;
  assign n32771 = ~n14801 ;
  assign n14802 = n13775 & n32771 ;
  assign n13320 = n895 & n32488 ;
  assign n10826 = n2849 & n10818 ;
  assign n10843 = n2861 & n10841 ;
  assign n14803 = n10826 | n10843 ;
  assign n14804 = n894 & n31998 ;
  assign n14805 = n14803 | n14804 ;
  assign n14806 = n13320 | n14805 ;
  assign n14807 = x29 | n14806 ;
  assign n14808 = x29 & n14806 ;
  assign n32772 = ~n14808 ;
  assign n14809 = n14807 & n32772 ;
  assign n32773 = ~n14809 ;
  assign n14811 = n14802 & n32773 ;
  assign n14810 = n14802 & n14809 ;
  assign n14812 = n14802 | n14809 ;
  assign n32774 = ~n14810 ;
  assign n14813 = n32774 & n14812 ;
  assign n13772 = n13751 | n13771 ;
  assign n14814 = n13751 & n13771 ;
  assign n32775 = ~n14814 ;
  assign n14815 = n13772 & n32775 ;
  assign n13384 = n895 & n13382 ;
  assign n10849 = n2849 & n10841 ;
  assign n10875 = n2861 & n10865 ;
  assign n14816 = n10849 | n10875 ;
  assign n14817 = n894 & n10818 ;
  assign n14818 = n14816 | n14817 ;
  assign n14819 = n13384 | n14818 ;
  assign n14820 = x29 | n14819 ;
  assign n14821 = x29 & n14819 ;
  assign n32776 = ~n14821 ;
  assign n14822 = n14820 & n32776 ;
  assign n32777 = ~n14822 ;
  assign n14824 = n14815 & n32777 ;
  assign n32778 = ~n13705 ;
  assign n13706 = n13685 & n32778 ;
  assign n32779 = ~n13685 ;
  assign n14825 = n32779 & n13705 ;
  assign n14826 = n13706 | n14825 ;
  assign n13458 = n895 & n13456 ;
  assign n10871 = n2849 & n10865 ;
  assign n10903 = n2861 & n10892 ;
  assign n14827 = n10871 | n10903 ;
  assign n14828 = n894 & n10841 ;
  assign n14829 = n14827 | n14828 ;
  assign n14830 = n13458 | n14829 ;
  assign n14831 = x29 | n14830 ;
  assign n14832 = x29 & n14830 ;
  assign n32780 = ~n14832 ;
  assign n14833 = n14831 & n32780 ;
  assign n14835 = n14826 | n14833 ;
  assign n14834 = n14826 & n14833 ;
  assign n32781 = ~n14834 ;
  assign n14836 = n32781 & n14835 ;
  assign n13645 = n13635 | n13644 ;
  assign n14837 = n13635 & n13644 ;
  assign n32782 = ~n14837 ;
  assign n14838 = n13645 & n32782 ;
  assign n13527 = n895 & n32502 ;
  assign n10901 = n2849 & n10892 ;
  assign n10928 = n2861 & n32503 ;
  assign n14839 = n10901 | n10928 ;
  assign n14840 = n894 & n10865 ;
  assign n14841 = n14839 | n14840 ;
  assign n14842 = n13527 | n14841 ;
  assign n14843 = x29 | n14842 ;
  assign n14844 = x29 & n14842 ;
  assign n32783 = ~n14844 ;
  assign n14845 = n14843 & n32783 ;
  assign n32784 = ~n14838 ;
  assign n14846 = n32784 & n14845 ;
  assign n13583 = n13549 & n13582 ;
  assign n14847 = n13549 | n13582 ;
  assign n32785 = ~n13583 ;
  assign n14848 = n32785 & n14847 ;
  assign n13759 = n895 & n13756 ;
  assign n10930 = n2849 & n32503 ;
  assign n10965 = n2861 & n10940 ;
  assign n14849 = n10930 | n10965 ;
  assign n14850 = n894 & n10892 ;
  assign n14851 = n14849 | n14850 ;
  assign n14852 = n13759 | n14851 ;
  assign n14853 = x29 | n14852 ;
  assign n14854 = x29 & n14852 ;
  assign n32786 = ~n14854 ;
  assign n14855 = n14853 & n32786 ;
  assign n32787 = ~n14855 ;
  assign n14857 = n14848 & n32787 ;
  assign n14858 = n891 & n32507 ;
  assign n10993 = n10974 & n10992 ;
  assign n32788 = ~n10993 ;
  assign n14859 = n32788 & n10994 ;
  assign n14860 = n895 & n14859 ;
  assign n14869 = n894 & n31995 ;
  assign n14870 = n2849 & n32507 ;
  assign n14871 = n14869 | n14870 ;
  assign n14872 = n14860 | n14871 ;
  assign n14873 = n14858 | n14872 ;
  assign n14874 = x29 & n14873 ;
  assign n10960 = n894 & n10940 ;
  assign n14875 = n2849 & n31995 ;
  assign n14876 = n2861 & n32507 ;
  assign n14877 = n14875 | n14876 ;
  assign n14878 = n10960 | n14877 ;
  assign n14879 = n895 & n13637 ;
  assign n14880 = n14878 | n14879 ;
  assign n14882 = n14874 | n14880 ;
  assign n32789 = ~n14882 ;
  assign n14883 = x29 & n32789 ;
  assign n14884 = n108 & n32507 ;
  assign n14886 = n14883 | n14884 ;
  assign n13693 = n895 & n13690 ;
  assign n10961 = n2849 & n10940 ;
  assign n10978 = n2861 & n31995 ;
  assign n14887 = n10961 | n10978 ;
  assign n14888 = n894 & n32503 ;
  assign n14889 = n14887 | n14888 ;
  assign n14890 = n13693 | n14889 ;
  assign n32790 = ~n14890 ;
  assign n14891 = x29 & n32790 ;
  assign n14892 = n30024 & n14890 ;
  assign n14893 = n14891 | n14892 ;
  assign n14894 = n14886 & n14893 ;
  assign n32791 = ~n14848 ;
  assign n14856 = n32791 & n14855 ;
  assign n14895 = n14856 | n14857 ;
  assign n14896 = n14894 | n14895 ;
  assign n32792 = ~n14857 ;
  assign n14897 = n32792 & n14896 ;
  assign n32793 = ~n14845 ;
  assign n14898 = n14838 & n32793 ;
  assign n14899 = n14846 | n14898 ;
  assign n32794 = ~n14899 ;
  assign n14900 = n14897 & n32794 ;
  assign n14901 = n14846 | n14900 ;
  assign n32795 = ~n14901 ;
  assign n14902 = n14836 & n32795 ;
  assign n32796 = ~n14902 ;
  assign n14903 = n14835 & n32796 ;
  assign n32797 = ~n14815 ;
  assign n14823 = n32797 & n14822 ;
  assign n14904 = n14823 | n14824 ;
  assign n14906 = n14903 | n14904 ;
  assign n32798 = ~n14824 ;
  assign n14907 = n32798 & n14906 ;
  assign n14909 = n14813 | n14907 ;
  assign n32799 = ~n14811 ;
  assign n14910 = n32799 & n14909 ;
  assign n32800 = ~n14910 ;
  assign n14912 = n14800 & n32800 ;
  assign n32801 = ~n14912 ;
  assign n14913 = n14798 & n32801 ;
  assign n32802 = ~n14913 ;
  assign n14915 = n14787 & n32802 ;
  assign n32803 = ~n14915 ;
  assign n14916 = n14785 & n32803 ;
  assign n14773 = n14765 & n14772 ;
  assign n32804 = ~n14773 ;
  assign n14917 = n32804 & n14774 ;
  assign n32805 = ~n14916 ;
  assign n14919 = n32805 & n14917 ;
  assign n32806 = ~n14919 ;
  assign n14920 = n14774 & n32806 ;
  assign n32807 = ~n14920 ;
  assign n14922 = n14763 & n32807 ;
  assign n32808 = ~n14922 ;
  assign n14923 = n14761 & n32808 ;
  assign n32809 = ~n14923 ;
  assign n14925 = n14750 & n32809 ;
  assign n32810 = ~n14925 ;
  assign n14926 = n14748 & n32810 ;
  assign n32811 = ~n14736 ;
  assign n14927 = n14729 & n32811 ;
  assign n14928 = n14737 | n14927 ;
  assign n32812 = ~n14928 ;
  assign n14929 = n14926 & n32812 ;
  assign n14930 = n14737 | n14929 ;
  assign n32813 = ~n14930 ;
  assign n14931 = n14727 & n32813 ;
  assign n32814 = ~n14931 ;
  assign n14932 = n14725 & n32814 ;
  assign n32815 = ~n14932 ;
  assign n14934 = n14714 & n32815 ;
  assign n13850 = n4686 & n32557 ;
  assign n12548 = n4726 & n32354 ;
  assign n13085 = n4706 & n13077 ;
  assign n14935 = n12548 | n13085 ;
  assign n14936 = n4748 & n32456 ;
  assign n14937 = n14935 | n14936 ;
  assign n14938 = n13850 | n14937 ;
  assign n32816 = ~n14938 ;
  assign n14939 = x20 & n32816 ;
  assign n14940 = n30374 & n14938 ;
  assign n14941 = n14939 | n14940 ;
  assign n32817 = ~n14714 ;
  assign n14933 = n32817 & n14932 ;
  assign n14942 = n14933 | n14934 ;
  assign n14943 = n14941 | n14942 ;
  assign n32818 = ~n14934 ;
  assign n14944 = n32818 & n14943 ;
  assign n32819 = ~n14944 ;
  assign n14946 = n14712 & n32819 ;
  assign n14945 = n14712 & n14944 ;
  assign n14947 = n14712 | n14944 ;
  assign n32820 = ~n14945 ;
  assign n14948 = n32820 & n14947 ;
  assign n13117 = n4686 & n32455 ;
  assign n13062 = n4706 & n32456 ;
  assign n13086 = n4726 & n13077 ;
  assign n14949 = n13062 | n13086 ;
  assign n14950 = n4748 & n13027 ;
  assign n14951 = n14949 | n14950 ;
  assign n14952 = n13117 | n14951 ;
  assign n32821 = ~n14952 ;
  assign n14953 = x20 & n32821 ;
  assign n14954 = n30374 & n14952 ;
  assign n14955 = n14953 | n14954 ;
  assign n14956 = n14948 | n14955 ;
  assign n32822 = ~n14946 ;
  assign n14957 = n32822 & n14956 ;
  assign n14959 = n14710 | n14957 ;
  assign n32823 = ~n14536 ;
  assign n14563 = n14101 & n32823 ;
  assign n32824 = ~n14101 ;
  assign n14960 = n32824 & n14536 ;
  assign n14961 = n14563 | n14960 ;
  assign n14962 = n14559 | n14561 ;
  assign n14963 = n14961 | n14962 ;
  assign n14964 = n14961 & n14962 ;
  assign n32825 = ~n14964 ;
  assign n14965 = n14963 & n32825 ;
  assign n14966 = n37300 & n14965 ;
  assign n14111 = n5144 & n14101 ;
  assign n14136 = n5166 & n14124 ;
  assign n14977 = n14111 | n14136 ;
  assign n14978 = n5191 & n14536 ;
  assign n14979 = n14977 | n14978 ;
  assign n14980 = n14966 | n14979 ;
  assign n32826 = ~n14980 ;
  assign n14981 = x17 & n32826 ;
  assign n14982 = n30580 & n14980 ;
  assign n14983 = n14981 | n14982 ;
  assign n32827 = ~n14710 ;
  assign n14958 = n32827 & n14957 ;
  assign n32828 = ~n14957 ;
  assign n14984 = n14710 & n32828 ;
  assign n14985 = n14958 | n14984 ;
  assign n32829 = ~n14983 ;
  assign n14986 = n32829 & n14985 ;
  assign n32830 = ~n14986 ;
  assign n14987 = n14959 & n32830 ;
  assign n32831 = ~n14708 ;
  assign n14988 = n32831 & n14987 ;
  assign n5798 = n3329 & n30545 ;
  assign n6447 = n889 & n6445 ;
  assign n14989 = n5798 | n6447 ;
  assign n14990 = n368 | n4916 ;
  assign n14991 = n5836 | n14990 ;
  assign n14992 = n2905 | n5604 ;
  assign n14993 = n4895 | n14992 ;
  assign n14994 = n497 | n5860 ;
  assign n14995 = n3197 | n14994 ;
  assign n14996 = n5906 | n14995 ;
  assign n14997 = n1229 | n1625 ;
  assign n14998 = n3736 | n14997 ;
  assign n14999 = n416 | n1049 ;
  assign n15000 = n770 | n1146 ;
  assign n15001 = n14999 | n15000 ;
  assign n15002 = n14998 | n15001 ;
  assign n15003 = n4907 | n15002 ;
  assign n15004 = n14996 | n15003 ;
  assign n15005 = n5820 | n15004 ;
  assign n15006 = n14993 | n15005 ;
  assign n15007 = n14991 | n15006 ;
  assign n32832 = ~n14342 ;
  assign n15009 = n32832 & n15007 ;
  assign n32833 = ~n15007 ;
  assign n15008 = n14342 & n32833 ;
  assign n15010 = n15008 | n15009 ;
  assign n15011 = x29 | n15010 ;
  assign n32834 = ~n15009 ;
  assign n15012 = n32834 & n15011 ;
  assign n15013 = n212 | n2161 ;
  assign n15014 = n2394 | n15013 ;
  assign n15015 = n4879 | n4896 ;
  assign n15016 = n15014 | n15015 ;
  assign n15017 = n3219 | n15016 ;
  assign n15018 = n4253 | n5776 ;
  assign n15019 = n5894 | n15018 ;
  assign n15020 = n15017 | n15019 ;
  assign n32835 = ~n15020 ;
  assign n15021 = n5828 & n32835 ;
  assign n32836 = ~n14991 ;
  assign n15022 = n32836 & n15021 ;
  assign n15023 = n15012 & n15022 ;
  assign n15024 = n15012 | n15022 ;
  assign n32837 = ~n15023 ;
  assign n15025 = n32837 & n15024 ;
  assign n15026 = n14989 | n15025 ;
  assign n15027 = n14989 & n15025 ;
  assign n32838 = ~n15027 ;
  assign n15028 = n15026 & n32838 ;
  assign n15029 = x29 & n15010 ;
  assign n32839 = ~n15029 ;
  assign n15030 = n15011 & n32839 ;
  assign n15031 = n32832 & n14358 ;
  assign n32840 = ~n15031 ;
  assign n15032 = n14398 & n32840 ;
  assign n15033 = n15030 & n15032 ;
  assign n15034 = n15030 | n15032 ;
  assign n32841 = ~n15033 ;
  assign n15035 = n32841 & n15034 ;
  assign n5931 = n889 & n30540 ;
  assign n15036 = n3311 & n30530 ;
  assign n15037 = n3329 & n30535 ;
  assign n15038 = n15036 | n15037 ;
  assign n15039 = n5931 | n15038 ;
  assign n15041 = n15035 & n15039 ;
  assign n15042 = n15033 | n15041 ;
  assign n15043 = n15028 | n15042 ;
  assign n15044 = n15028 & n15042 ;
  assign n32842 = ~n15044 ;
  assign n15045 = n15043 & n32842 ;
  assign n32843 = ~n15039 ;
  assign n15040 = n15035 & n32843 ;
  assign n32844 = ~n15035 ;
  assign n15046 = n32844 & n15039 ;
  assign n15047 = n15040 | n15046 ;
  assign n32845 = ~n14406 ;
  assign n15048 = n32845 & n14409 ;
  assign n15050 = n15047 | n15048 ;
  assign n15049 = n15047 & n15048 ;
  assign n32846 = ~n15049 ;
  assign n15051 = n32846 & n15050 ;
  assign n32847 = ~n14441 ;
  assign n15052 = n32847 & n14488 ;
  assign n32848 = ~n15052 ;
  assign n15054 = n15051 & n32848 ;
  assign n32849 = ~n15054 ;
  assign n15055 = n15050 & n32849 ;
  assign n15056 = n15045 | n15055 ;
  assign n15057 = n15045 & n15055 ;
  assign n32850 = ~n15057 ;
  assign n15058 = n15056 & n32850 ;
  assign n15078 = n32706 & n14560 ;
  assign n32851 = ~n15078 ;
  assign n15079 = n14490 & n32851 ;
  assign n15053 = n15051 & n15052 ;
  assign n15080 = n15051 | n15052 ;
  assign n32852 = ~n15053 ;
  assign n15081 = n32852 & n15080 ;
  assign n32853 = ~n15079 ;
  assign n15083 = n32853 & n15081 ;
  assign n15105 = n14513 & n32733 ;
  assign n15106 = n14490 | n15105 ;
  assign n32854 = ~n15081 ;
  assign n15107 = n32854 & n15106 ;
  assign n15108 = n15083 | n15107 ;
  assign n15109 = n15058 | n15108 ;
  assign n15110 = n15058 & n15108 ;
  assign n32855 = ~n15110 ;
  assign n15111 = n15109 & n32855 ;
  assign n15112 = n5937 & n15111 ;
  assign n14505 = n5994 & n32707 ;
  assign n15101 = n5970 & n15081 ;
  assign n15124 = n14505 | n15101 ;
  assign n32856 = ~n15058 ;
  assign n15125 = n6018 & n32856 ;
  assign n15126 = n15124 | n15125 ;
  assign n15127 = n15112 | n15126 ;
  assign n15128 = x14 | n15127 ;
  assign n15129 = x14 & n15127 ;
  assign n32857 = ~n15129 ;
  assign n15130 = n15128 & n32857 ;
  assign n32858 = ~n14987 ;
  assign n15131 = n14708 & n32858 ;
  assign n15132 = n14988 | n15131 ;
  assign n32859 = ~n15132 ;
  assign n15133 = n15130 & n32859 ;
  assign n15134 = n14988 | n15133 ;
  assign n32860 = ~n14706 ;
  assign n15136 = n32860 & n15134 ;
  assign n15137 = n249 | n560 ;
  assign n15138 = n721 | n15137 ;
  assign n15139 = n1050 | n1662 ;
  assign n15140 = n15138 | n15139 ;
  assign n32861 = ~n15140 ;
  assign n15141 = n4917 & n32861 ;
  assign n32862 = ~n5779 ;
  assign n15142 = n32862 & n15141 ;
  assign n32863 = ~n14996 ;
  assign n15143 = n32863 & n15142 ;
  assign n32864 = ~n5898 ;
  assign n15144 = n32864 & n15143 ;
  assign n15145 = n15022 & n15144 ;
  assign n15146 = n15022 | n15144 ;
  assign n32865 = ~n15145 ;
  assign n15147 = n32865 & n15146 ;
  assign n32866 = ~n15012 ;
  assign n15148 = n32866 & n15022 ;
  assign n32867 = ~n15025 ;
  assign n15149 = n14989 & n32867 ;
  assign n15150 = n15148 | n15149 ;
  assign n32868 = ~n15150 ;
  assign n15151 = n15147 & n32868 ;
  assign n32869 = ~n15147 ;
  assign n15152 = n32869 & n15150 ;
  assign n15153 = n15151 | n15152 ;
  assign n32870 = ~n15042 ;
  assign n15154 = n15028 & n32870 ;
  assign n32871 = ~n15154 ;
  assign n15155 = n15056 & n32871 ;
  assign n32872 = ~n15153 ;
  assign n15156 = n32872 & n15155 ;
  assign n32873 = ~n15155 ;
  assign n15157 = n15153 & n32873 ;
  assign n15158 = n15156 | n15157 ;
  assign n15123 = n15058 & n15083 ;
  assign n15180 = n32856 & n15107 ;
  assign n15181 = n15123 | n15180 ;
  assign n15182 = n15158 & n15181 ;
  assign n15183 = n15158 | n15181 ;
  assign n32874 = ~n15182 ;
  assign n15184 = n32874 & n15183 ;
  assign n32875 = ~n15184 ;
  assign n15185 = n5937 & n32875 ;
  assign n15064 = n5970 & n32856 ;
  assign n15099 = n5994 & n15081 ;
  assign n15196 = n15064 | n15099 ;
  assign n32876 = ~n15158 ;
  assign n15197 = n6018 & n32876 ;
  assign n15198 = n15196 | n15197 ;
  assign n15199 = n15185 | n15198 ;
  assign n15200 = x14 | n15199 ;
  assign n15201 = x14 & n15199 ;
  assign n32877 = ~n15201 ;
  assign n15202 = n15200 & n32877 ;
  assign n15135 = n14706 | n15134 ;
  assign n15203 = n14706 & n15134 ;
  assign n32878 = ~n15203 ;
  assign n15204 = n15135 & n32878 ;
  assign n32879 = ~n15204 ;
  assign n15205 = n15202 & n32879 ;
  assign n15206 = n15136 | n15205 ;
  assign n6214 = x11 & n6213 ;
  assign n15207 = n15153 | n15155 ;
  assign n32880 = ~n15151 ;
  assign n15208 = n32880 & n15207 ;
  assign n15209 = n4251 | n4879 ;
  assign n15210 = n679 | n1049 ;
  assign n15211 = n185 | n15210 ;
  assign n15212 = n5860 | n15211 ;
  assign n15213 = n5904 | n15212 ;
  assign n15214 = n15209 | n15213 ;
  assign n32881 = ~n15214 ;
  assign n15215 = n5849 & n32881 ;
  assign n32882 = ~n15215 ;
  assign n15216 = n15022 & n32882 ;
  assign n15217 = n32865 & n15215 ;
  assign n15218 = n15216 | n15217 ;
  assign n15220 = n15208 | n15218 ;
  assign n15221 = x30 | n15220 ;
  assign n15224 = x10 & n15221 ;
  assign n32883 = ~n15221 ;
  assign n15233 = x11 & n32883 ;
  assign n15247 = n6213 | n15233 ;
  assign n15248 = n15224 | n15247 ;
  assign n32884 = ~n6214 ;
  assign n15249 = n32884 & n15248 ;
  assign n15251 = n15206 & n15249 ;
  assign n15219 = n15208 & n15218 ;
  assign n32885 = ~n15219 ;
  assign n15252 = n32885 & n15220 ;
  assign n15258 = n15058 | n15107 ;
  assign n32886 = ~n15258 ;
  assign n15259 = n15158 & n32886 ;
  assign n32887 = ~n15083 ;
  assign n15257 = n15058 & n32887 ;
  assign n15260 = n32876 & n15257 ;
  assign n15261 = n15259 | n15260 ;
  assign n15262 = n15252 & n15261 ;
  assign n15263 = n15252 | n15261 ;
  assign n32888 = ~n15262 ;
  assign n15264 = n32888 & n15263 ;
  assign n32889 = ~n15264 ;
  assign n15265 = n5937 & n32889 ;
  assign n15069 = n5994 & n32856 ;
  assign n15171 = n5970 & n32876 ;
  assign n15276 = n15069 | n15171 ;
  assign n32890 = ~n15252 ;
  assign n15277 = n6018 & n32890 ;
  assign n15278 = n15276 | n15277 ;
  assign n15279 = n15265 | n15278 ;
  assign n32891 = ~n15279 ;
  assign n15280 = x14 & n32891 ;
  assign n15281 = n30547 & n15279 ;
  assign n15282 = n15280 | n15281 ;
  assign n15283 = n32707 & n14567 ;
  assign n15082 = n15078 | n15081 ;
  assign n15284 = n15078 & n15081 ;
  assign n32892 = ~n15284 ;
  assign n15285 = n15082 & n32892 ;
  assign n15286 = n15283 & n15285 ;
  assign n15287 = n15283 | n15285 ;
  assign n32893 = ~n15286 ;
  assign n15288 = n32893 & n15287 ;
  assign n15289 = n37300 & n15288 ;
  assign n14504 = n5144 & n32707 ;
  assign n14526 = n5166 & n32706 ;
  assign n15300 = n14504 | n14526 ;
  assign n15301 = n5191 & n15081 ;
  assign n15302 = n15300 | n15301 ;
  assign n15303 = n15289 | n15302 ;
  assign n32894 = ~n15303 ;
  assign n15304 = x17 & n32894 ;
  assign n15305 = n30580 & n15303 ;
  assign n15306 = n15304 | n15305 ;
  assign n14968 = n4686 & n14965 ;
  assign n14110 = n4706 & n14101 ;
  assign n14130 = n4726 & n14124 ;
  assign n15307 = n14110 | n14130 ;
  assign n15308 = n4748 & n14536 ;
  assign n15309 = n15307 | n15308 ;
  assign n15310 = n14968 | n15309 ;
  assign n32895 = ~n15310 ;
  assign n15311 = x20 & n32895 ;
  assign n15312 = n30374 & n15310 ;
  assign n15313 = n15311 | n15312 ;
  assign n14658 = n4135 & n14655 ;
  assign n13040 = n4148 & n13027 ;
  assign n13056 = n4185 & n32456 ;
  assign n15314 = n13040 | n13056 ;
  assign n15315 = n4165 & n14147 ;
  assign n15316 = n15314 | n15315 ;
  assign n15317 = n14658 | n15316 ;
  assign n32896 = ~n15317 ;
  assign n15318 = x23 & n32896 ;
  assign n15319 = n30030 & n15317 ;
  assign n15320 = n15318 | n15319 ;
  assign n14257 = n3791 & n32641 ;
  assign n12556 = n3802 & n32354 ;
  assign n12579 = n209 & n12570 ;
  assign n15321 = n12556 | n12579 ;
  assign n15322 = n3818 & n13077 ;
  assign n15323 = n15321 | n15322 ;
  assign n15324 = n14257 | n15323 ;
  assign n32897 = ~n15324 ;
  assign n15325 = x26 & n32897 ;
  assign n15326 = n30019 & n15324 ;
  assign n15327 = n15325 | n15326 ;
  assign n13827 = n895 & n32550 ;
  assign n12149 = n2849 & n32253 ;
  assign n12167 = n2861 & n12161 ;
  assign n15328 = n12149 | n12167 ;
  assign n15329 = n894 & n12595 ;
  assign n15330 = n15328 | n15329 ;
  assign n15331 = n13827 | n15330 ;
  assign n32898 = ~n15331 ;
  assign n15332 = x29 & n32898 ;
  assign n15333 = n30024 & n15331 ;
  assign n15334 = n15332 | n15333 ;
  assign n32899 = ~n11072 ;
  assign n15335 = n584 & n32899 ;
  assign n32900 = ~n11075 ;
  assign n15336 = n32900 & n11501 ;
  assign n15337 = n15335 | n15336 ;
  assign n15338 = n72 | n391 ;
  assign n15339 = n30042 & n15338 ;
  assign n15340 = n1311 | n2512 ;
  assign n15341 = n11126 | n15340 ;
  assign n15342 = n83 | n187 ;
  assign n15343 = n464 | n479 ;
  assign n15344 = n15342 | n15343 ;
  assign n15345 = n1901 | n15344 ;
  assign n15346 = n15341 | n15345 ;
  assign n15347 = n5552 | n15346 ;
  assign n15348 = n815 | n1943 ;
  assign n15349 = n2394 | n14322 ;
  assign n15350 = n15348 | n15349 ;
  assign n15351 = n13218 | n15350 ;
  assign n15352 = n15347 | n15351 ;
  assign n32901 = ~n15352 ;
  assign n15353 = n838 & n32901 ;
  assign n32902 = ~n4333 ;
  assign n15354 = n32902 & n15353 ;
  assign n15355 = n30148 & n15354 ;
  assign n15356 = n15339 & n15355 ;
  assign n15357 = n15339 | n15355 ;
  assign n32903 = ~n15356 ;
  assign n15358 = n32903 & n15357 ;
  assign n11873 = n889 & n32178 ;
  assign n11442 = n3329 & n11430 ;
  assign n11481 = n3311 & n11476 ;
  assign n15359 = n11442 | n11481 ;
  assign n15360 = n3343 & n32176 ;
  assign n15361 = n15359 | n15360 ;
  assign n15362 = n11873 | n15361 ;
  assign n32904 = ~n15362 ;
  assign n15363 = n15358 & n32904 ;
  assign n32905 = ~n15358 ;
  assign n15364 = n32905 & n15362 ;
  assign n15365 = n15363 | n15364 ;
  assign n15366 = n15337 | n15365 ;
  assign n15367 = n15337 & n15365 ;
  assign n32906 = ~n15367 ;
  assign n15368 = n15366 & n32906 ;
  assign n15369 = n15334 | n15368 ;
  assign n15370 = n15334 & n15368 ;
  assign n32907 = ~n15370 ;
  assign n15371 = n15369 & n32907 ;
  assign n32908 = ~n11898 ;
  assign n15372 = n32908 & n12211 ;
  assign n15373 = n11896 | n15372 ;
  assign n32909 = ~n15373 ;
  assign n15374 = n15371 & n32909 ;
  assign n32910 = ~n15371 ;
  assign n15375 = n32910 & n15373 ;
  assign n15376 = n15374 | n15375 ;
  assign n15377 = n15327 | n15376 ;
  assign n15378 = n15327 & n15376 ;
  assign n32911 = ~n15378 ;
  assign n15379 = n15377 & n32911 ;
  assign n15380 = n12702 & n32371 ;
  assign n15381 = n15379 & n15380 ;
  assign n15382 = n15379 | n15380 ;
  assign n32912 = ~n15381 ;
  assign n15383 = n32912 & n15382 ;
  assign n15384 = n15320 | n15383 ;
  assign n15385 = n15320 & n15383 ;
  assign n32913 = ~n15385 ;
  assign n15386 = n15384 & n32913 ;
  assign n15387 = n13133 | n13869 ;
  assign n32914 = ~n13131 ;
  assign n15388 = n32914 & n15387 ;
  assign n15389 = n15386 & n15388 ;
  assign n15390 = n15386 | n15388 ;
  assign n32915 = ~n15389 ;
  assign n15391 = n32915 & n15390 ;
  assign n15392 = n15313 | n15391 ;
  assign n15393 = n15313 & n15391 ;
  assign n32916 = ~n15393 ;
  assign n15394 = n15392 & n32916 ;
  assign n32917 = ~n14206 ;
  assign n15395 = n32917 & n14307 ;
  assign n15396 = n14205 | n15395 ;
  assign n32918 = ~n15396 ;
  assign n15397 = n15394 & n32918 ;
  assign n32919 = ~n15394 ;
  assign n15398 = n32919 & n15396 ;
  assign n15399 = n15397 | n15398 ;
  assign n15400 = n15306 | n15399 ;
  assign n15401 = n15306 & n15399 ;
  assign n32920 = ~n15401 ;
  assign n15402 = n15400 & n32920 ;
  assign n32921 = ~n14310 ;
  assign n15403 = n32921 & n14588 ;
  assign n15404 = n14704 | n15403 ;
  assign n32922 = ~n15404 ;
  assign n15405 = n15402 & n32922 ;
  assign n32923 = ~n15402 ;
  assign n15406 = n32923 & n15404 ;
  assign n15407 = n15405 | n15406 ;
  assign n15408 = n15282 | n15407 ;
  assign n15409 = n15282 & n15407 ;
  assign n32924 = ~n15409 ;
  assign n15410 = n15408 & n32924 ;
  assign n32925 = ~n15206 ;
  assign n15250 = n32925 & n15249 ;
  assign n32926 = ~n15249 ;
  assign n15411 = n15206 & n32926 ;
  assign n15412 = n15250 | n15411 ;
  assign n32927 = ~n15410 ;
  assign n15413 = n32927 & n15412 ;
  assign n15415 = n15251 | n15413 ;
  assign n15114 = n37300 & n15111 ;
  assign n14503 = n5166 & n32707 ;
  assign n15100 = n5144 & n15081 ;
  assign n15416 = n14503 | n15100 ;
  assign n15417 = n5191 & n32856 ;
  assign n15418 = n15416 | n15417 ;
  assign n15419 = n15114 | n15418 ;
  assign n32928 = ~n15419 ;
  assign n15420 = x17 & n32928 ;
  assign n15421 = n30580 & n15419 ;
  assign n15422 = n15420 | n15421 ;
  assign n14685 = n4686 & n32735 ;
  assign n14105 = n4726 & n14101 ;
  assign n14543 = n4706 & n14536 ;
  assign n15423 = n14105 | n14543 ;
  assign n15424 = n4748 & n32706 ;
  assign n15425 = n15423 | n15424 ;
  assign n15426 = n14685 | n15425 ;
  assign n32929 = ~n15426 ;
  assign n15427 = x20 & n32929 ;
  assign n15428 = n30374 & n15426 ;
  assign n15429 = n15427 | n15428 ;
  assign n14286 = n4135 & n14283 ;
  assign n13039 = n4185 & n13027 ;
  assign n14157 = n4148 & n14147 ;
  assign n15430 = n13039 | n14157 ;
  assign n15431 = n4165 & n14295 ;
  assign n15432 = n15430 | n15431 ;
  assign n15433 = n14286 | n15432 ;
  assign n32930 = ~n15433 ;
  assign n15434 = x23 & n32930 ;
  assign n15435 = n30030 & n15433 ;
  assign n15436 = n15434 | n15435 ;
  assign n13851 = n3791 & n32557 ;
  assign n12555 = n209 & n32354 ;
  assign n13082 = n3802 & n13077 ;
  assign n15437 = n12555 | n13082 ;
  assign n15438 = n3818 & n32456 ;
  assign n15439 = n15437 | n15438 ;
  assign n15440 = n13851 | n15439 ;
  assign n32931 = ~n15440 ;
  assign n15441 = x26 & n32931 ;
  assign n15442 = n30019 & n15440 ;
  assign n15443 = n15441 | n15442 ;
  assign n12685 = n895 & n12681 ;
  assign n12142 = n2861 & n32253 ;
  assign n12602 = n2849 & n12595 ;
  assign n15444 = n12142 | n12602 ;
  assign n15445 = n894 & n12570 ;
  assign n15446 = n15444 | n15445 ;
  assign n15447 = n12685 | n15446 ;
  assign n15448 = x29 | n15447 ;
  assign n15449 = x29 & n15447 ;
  assign n32932 = ~n15449 ;
  assign n15450 = n15448 & n32932 ;
  assign n15451 = n507 | n4086 ;
  assign n15452 = n5816 | n15451 ;
  assign n15453 = n1467 | n15452 ;
  assign n15454 = n4072 | n15453 ;
  assign n15455 = n224 | n232 ;
  assign n15456 = n359 | n15455 ;
  assign n15457 = n904 | n15456 ;
  assign n15458 = n124 | n412 ;
  assign n15459 = n1830 | n15458 ;
  assign n15460 = n15457 | n15459 ;
  assign n15461 = n13724 | n15460 ;
  assign n15462 = n15454 | n15461 ;
  assign n15463 = n11938 | n15462 ;
  assign n32933 = ~n15463 ;
  assign n15464 = n13603 & n32933 ;
  assign n32934 = ~n15464 ;
  assign n15465 = n15355 & n32934 ;
  assign n32935 = ~n15355 ;
  assign n15466 = n32935 & n15464 ;
  assign n15467 = n15465 | n15466 ;
  assign n32936 = ~n15339 ;
  assign n15468 = n32936 & n15355 ;
  assign n15469 = n15364 | n15468 ;
  assign n15470 = n15467 | n15469 ;
  assign n15471 = n15467 & n15469 ;
  assign n32937 = ~n15471 ;
  assign n15472 = n15470 & n32937 ;
  assign n12657 = n889 & n32362 ;
  assign n11438 = n3311 & n11430 ;
  assign n11848 = n3329 & n32176 ;
  assign n15473 = n11438 | n11848 ;
  assign n15474 = n3343 & n12161 ;
  assign n15475 = n15473 | n15474 ;
  assign n15476 = n12657 | n15475 ;
  assign n32938 = ~n15476 ;
  assign n15477 = n15472 & n32938 ;
  assign n32939 = ~n15472 ;
  assign n15478 = n32939 & n15476 ;
  assign n15479 = n15477 | n15478 ;
  assign n32940 = ~n15479 ;
  assign n15480 = n15450 & n32940 ;
  assign n32941 = ~n15450 ;
  assign n15481 = n32941 & n15479 ;
  assign n15482 = n15480 | n15481 ;
  assign n32942 = ~n15337 ;
  assign n15483 = n32942 & n15365 ;
  assign n32943 = ~n15483 ;
  assign n15484 = n15369 & n32943 ;
  assign n32944 = ~n15482 ;
  assign n15485 = n32944 & n15484 ;
  assign n32945 = ~n15484 ;
  assign n15486 = n15482 & n32945 ;
  assign n15487 = n15485 | n15486 ;
  assign n15488 = n15443 | n15487 ;
  assign n15489 = n15443 & n15487 ;
  assign n32946 = ~n15489 ;
  assign n15490 = n15488 & n32946 ;
  assign n32947 = ~n15374 ;
  assign n15491 = n32947 & n15377 ;
  assign n15492 = n15490 & n15491 ;
  assign n15493 = n15490 | n15491 ;
  assign n32948 = ~n15492 ;
  assign n15494 = n32948 & n15493 ;
  assign n15495 = n15436 | n15494 ;
  assign n15496 = n15436 & n15494 ;
  assign n32949 = ~n15496 ;
  assign n15497 = n15495 & n32949 ;
  assign n32950 = ~n15380 ;
  assign n15498 = n15379 & n32950 ;
  assign n32951 = ~n15498 ;
  assign n15499 = n15384 & n32951 ;
  assign n32952 = ~n15497 ;
  assign n15500 = n32952 & n15499 ;
  assign n32953 = ~n15499 ;
  assign n15501 = n15497 & n32953 ;
  assign n15502 = n15500 | n15501 ;
  assign n15503 = n15429 | n15502 ;
  assign n15504 = n15429 & n15502 ;
  assign n32954 = ~n15504 ;
  assign n15505 = n15503 & n32954 ;
  assign n32955 = ~n15388 ;
  assign n15506 = n15386 & n32955 ;
  assign n32956 = ~n15506 ;
  assign n15507 = n15392 & n32956 ;
  assign n15508 = n15505 & n15507 ;
  assign n15509 = n15505 | n15507 ;
  assign n32957 = ~n15508 ;
  assign n15510 = n32957 & n15509 ;
  assign n15511 = n15422 | n15510 ;
  assign n15512 = n15422 & n15510 ;
  assign n32958 = ~n15512 ;
  assign n15513 = n15511 & n32958 ;
  assign n15514 = n15158 | n15257 ;
  assign n15515 = n15252 & n15514 ;
  assign n32959 = ~n15515 ;
  assign n15516 = n15221 & n32959 ;
  assign n32960 = ~n15516 ;
  assign n15525 = n15158 & n32960 ;
  assign n15526 = n15261 | n15525 ;
  assign n15527 = n5937 & n15526 ;
  assign n15172 = n5994 & n32876 ;
  assign n15230 = n6018 & n15221 ;
  assign n15537 = n15172 | n15230 ;
  assign n15538 = n5970 & n32890 ;
  assign n15539 = n15537 | n15538 ;
  assign n15540 = n15527 | n15539 ;
  assign n15541 = x14 | n15540 ;
  assign n15542 = x14 & n15540 ;
  assign n32961 = ~n15542 ;
  assign n15543 = n15541 & n32961 ;
  assign n32962 = ~n15397 ;
  assign n15544 = n32962 & n15400 ;
  assign n15545 = n15543 & n15544 ;
  assign n15546 = n15543 | n15544 ;
  assign n32963 = ~n15545 ;
  assign n15547 = n32963 & n15546 ;
  assign n15548 = n15513 & n15547 ;
  assign n15549 = n15513 | n15547 ;
  assign n32964 = ~n15548 ;
  assign n15550 = n32964 & n15549 ;
  assign n6187 = x10 | n6185 ;
  assign n15551 = n6187 & n32884 ;
  assign n32965 = ~n15405 ;
  assign n15552 = n32965 & n15408 ;
  assign n15553 = n15551 & n15552 ;
  assign n15554 = n15551 | n15552 ;
  assign n32966 = ~n15553 ;
  assign n15555 = n32966 & n15554 ;
  assign n32967 = ~n15550 ;
  assign n15556 = n32967 & n15555 ;
  assign n32968 = ~n15555 ;
  assign n15557 = n15550 & n32968 ;
  assign n15558 = n15556 | n15557 ;
  assign n32969 = ~n15415 ;
  assign n15559 = n32969 & n15558 ;
  assign n32970 = ~n15558 ;
  assign n15560 = n15415 & n32970 ;
  assign n15561 = n15559 | n15560 ;
  assign n15414 = n15410 & n15412 ;
  assign n15562 = n15410 | n15412 ;
  assign n32971 = ~n15414 ;
  assign n15563 = n32971 & n15562 ;
  assign n32972 = ~n15202 ;
  assign n15564 = n32972 & n15204 ;
  assign n15565 = n15205 | n15564 ;
  assign n15528 = n6272 & n15526 ;
  assign n15169 = n6244 & n32876 ;
  assign n15223 = n6217 & n15221 ;
  assign n15566 = n15169 | n15223 ;
  assign n15567 = n6190 & n32890 ;
  assign n15568 = n15566 | n15567 ;
  assign n15569 = n15528 | n15568 ;
  assign n15570 = x11 | n15569 ;
  assign n15571 = x11 & n15569 ;
  assign n32973 = ~n15571 ;
  assign n15572 = n15570 & n32973 ;
  assign n32974 = ~n14985 ;
  assign n15573 = n14983 & n32974 ;
  assign n15574 = n14986 | n15573 ;
  assign n15575 = n14948 & n14955 ;
  assign n32975 = ~n15575 ;
  assign n15576 = n14956 & n32975 ;
  assign n14185 = n37300 & n14183 ;
  assign n14135 = n5144 & n14124 ;
  assign n14155 = n5166 & n14147 ;
  assign n15577 = n14135 | n14155 ;
  assign n15578 = n5191 & n14196 ;
  assign n15579 = n15577 | n15578 ;
  assign n15580 = n14185 | n15579 ;
  assign n15581 = x17 | n15580 ;
  assign n15582 = x17 & n15580 ;
  assign n32976 = ~n15582 ;
  assign n15583 = n15581 & n32976 ;
  assign n32977 = ~n15583 ;
  assign n15585 = n15576 & n32977 ;
  assign n15584 = n15576 & n15583 ;
  assign n15586 = n15576 | n15583 ;
  assign n32978 = ~n15584 ;
  assign n15587 = n32978 & n15586 ;
  assign n15588 = n14941 & n14942 ;
  assign n32979 = ~n15588 ;
  assign n15589 = n14943 & n32979 ;
  assign n14287 = n37300 & n14283 ;
  assign n13035 = n5166 & n13027 ;
  assign n14156 = n5144 & n14147 ;
  assign n15590 = n13035 | n14156 ;
  assign n15591 = n5191 & n14295 ;
  assign n15592 = n15590 | n15591 ;
  assign n15593 = n14287 | n15592 ;
  assign n15594 = x17 | n15593 ;
  assign n15595 = x17 & n15593 ;
  assign n32980 = ~n15595 ;
  assign n15596 = n15594 & n32980 ;
  assign n32981 = ~n15596 ;
  assign n15598 = n15589 & n32981 ;
  assign n32982 = ~n15589 ;
  assign n15597 = n32982 & n15596 ;
  assign n15599 = n15597 | n15598 ;
  assign n32983 = ~n14727 ;
  assign n15600 = n32983 & n14930 ;
  assign n15601 = n14931 | n15600 ;
  assign n14259 = n4686 & n32641 ;
  assign n12546 = n4706 & n32354 ;
  assign n12582 = n4726 & n12570 ;
  assign n15602 = n12546 | n12582 ;
  assign n15603 = n4748 & n13077 ;
  assign n15604 = n15602 | n15603 ;
  assign n15605 = n14259 | n15604 ;
  assign n15606 = x20 | n15605 ;
  assign n15607 = x20 & n15605 ;
  assign n32984 = ~n15607 ;
  assign n15608 = n15606 & n32984 ;
  assign n15610 = n15601 | n15608 ;
  assign n32985 = ~n14926 ;
  assign n15611 = n32985 & n14928 ;
  assign n15612 = n14929 | n15611 ;
  assign n12196 = n4135 & n32255 ;
  assign n11843 = n4185 & n32176 ;
  assign n12166 = n4148 & n12161 ;
  assign n15613 = n11843 | n12166 ;
  assign n15614 = n4165 & n32253 ;
  assign n15615 = n15613 | n15614 ;
  assign n15616 = n12196 | n15615 ;
  assign n15617 = x23 | n15616 ;
  assign n15618 = x23 & n15616 ;
  assign n32986 = ~n15618 ;
  assign n15619 = n15617 & n32986 ;
  assign n32987 = ~n15619 ;
  assign n15621 = n15612 & n32987 ;
  assign n32988 = ~n15612 ;
  assign n15620 = n32988 & n15619 ;
  assign n15622 = n15620 | n15621 ;
  assign n14924 = n14750 & n14923 ;
  assign n15623 = n14750 | n14923 ;
  assign n32989 = ~n14924 ;
  assign n15624 = n32989 & n15623 ;
  assign n11515 = n3791 & n11511 ;
  assign n10668 = n3802 & n10656 ;
  assign n11048 = n209 & n10679 ;
  assign n15625 = n10668 | n11048 ;
  assign n15626 = n3818 & n11452 ;
  assign n15627 = n15625 | n15626 ;
  assign n15628 = n11515 | n15627 ;
  assign n15629 = x26 | n15628 ;
  assign n15630 = x26 & n15628 ;
  assign n32990 = ~n15630 ;
  assign n15631 = n15629 & n32990 ;
  assign n15633 = n15624 | n15631 ;
  assign n32991 = ~n15624 ;
  assign n15632 = n32991 & n15631 ;
  assign n32992 = ~n15631 ;
  assign n15634 = n15624 & n32992 ;
  assign n15635 = n15632 | n15634 ;
  assign n14921 = n14763 & n14920 ;
  assign n15636 = n14763 | n14920 ;
  assign n32993 = ~n14921 ;
  assign n15637 = n32993 & n15636 ;
  assign n11032 = n3791 & n11030 ;
  assign n10691 = n209 & n10681 ;
  assign n11050 = n3802 & n10679 ;
  assign n15638 = n10691 | n11050 ;
  assign n15639 = n3818 & n10656 ;
  assign n15640 = n15638 | n15639 ;
  assign n15641 = n11032 | n15640 ;
  assign n15642 = x26 | n15641 ;
  assign n15643 = x26 & n15641 ;
  assign n32994 = ~n15643 ;
  assign n15644 = n15642 & n32994 ;
  assign n15646 = n15637 | n15644 ;
  assign n32995 = ~n15637 ;
  assign n15645 = n32995 & n15644 ;
  assign n32996 = ~n15644 ;
  assign n15647 = n15637 & n32996 ;
  assign n15648 = n15645 | n15647 ;
  assign n14918 = n14916 & n14917 ;
  assign n15649 = n14916 | n14917 ;
  assign n32997 = ~n14918 ;
  assign n15650 = n32997 & n15649 ;
  assign n11539 = n3791 & n11536 ;
  assign n10683 = n3802 & n10681 ;
  assign n10719 = n209 & n10703 ;
  assign n15651 = n10683 | n10719 ;
  assign n15652 = n3818 & n10679 ;
  assign n15653 = n15651 | n15652 ;
  assign n15654 = n11539 | n15653 ;
  assign n15655 = x26 | n15654 ;
  assign n15656 = x26 & n15654 ;
  assign n32998 = ~n15656 ;
  assign n15657 = n15655 & n32998 ;
  assign n15659 = n15650 & n15657 ;
  assign n32999 = ~n15650 ;
  assign n15658 = n32999 & n15657 ;
  assign n33000 = ~n15657 ;
  assign n15660 = n15650 & n33000 ;
  assign n15661 = n15658 | n15660 ;
  assign n14914 = n14787 & n14913 ;
  assign n15662 = n14787 | n14913 ;
  assign n33001 = ~n14914 ;
  assign n15663 = n33001 & n15662 ;
  assign n13161 = n3791 & n13157 ;
  assign n10716 = n3802 & n10703 ;
  assign n10730 = n209 & n10727 ;
  assign n15664 = n10716 | n10730 ;
  assign n15665 = n3818 & n10681 ;
  assign n15666 = n15664 | n15665 ;
  assign n15667 = n13161 | n15666 ;
  assign n15668 = x26 | n15667 ;
  assign n15669 = x26 & n15667 ;
  assign n33002 = ~n15669 ;
  assign n15670 = n15668 & n33002 ;
  assign n15672 = n15663 | n15670 ;
  assign n14911 = n14800 & n14910 ;
  assign n15673 = n14800 | n14910 ;
  assign n33003 = ~n14911 ;
  assign n15674 = n33003 & n15673 ;
  assign n13188 = n3791 & n13182 ;
  assign n10733 = n3802 & n10727 ;
  assign n10760 = n209 & n31999 ;
  assign n15675 = n10733 | n10760 ;
  assign n15676 = n3818 & n13151 ;
  assign n15677 = n15675 | n15676 ;
  assign n15678 = n13188 | n15677 ;
  assign n15679 = x26 | n15678 ;
  assign n15680 = x26 & n15678 ;
  assign n33004 = ~n15680 ;
  assign n15681 = n15679 & n33004 ;
  assign n15683 = n15674 | n15681 ;
  assign n33005 = ~n15674 ;
  assign n15682 = n33005 & n15681 ;
  assign n33006 = ~n15681 ;
  assign n15684 = n15674 & n33006 ;
  assign n15685 = n15682 | n15684 ;
  assign n33007 = ~n14813 ;
  assign n14908 = n33007 & n14907 ;
  assign n33008 = ~n14907 ;
  assign n15686 = n14813 & n33008 ;
  assign n15687 = n14908 | n15686 ;
  assign n11689 = n3791 & n32125 ;
  assign n10754 = n3802 & n31999 ;
  assign n10776 = n209 & n10773 ;
  assign n15688 = n10754 | n10776 ;
  assign n15689 = n3818 & n10727 ;
  assign n15690 = n15688 | n15689 ;
  assign n15691 = n11689 | n15690 ;
  assign n15692 = x26 | n15691 ;
  assign n15693 = x26 & n15691 ;
  assign n33009 = ~n15693 ;
  assign n15694 = n15692 & n33009 ;
  assign n33010 = ~n15687 ;
  assign n15696 = n33010 & n15694 ;
  assign n15695 = n15687 & n15694 ;
  assign n15697 = n15687 | n15694 ;
  assign n33011 = ~n15695 ;
  assign n15698 = n33011 & n15697 ;
  assign n33012 = ~n14904 ;
  assign n14905 = n14903 & n33012 ;
  assign n33013 = ~n14903 ;
  assign n15699 = n33013 & n14904 ;
  assign n15700 = n14905 | n15699 ;
  assign n13232 = n3791 & n32477 ;
  assign n10786 = n3802 & n10773 ;
  assign n10800 = n209 & n31998 ;
  assign n15701 = n10786 | n10800 ;
  assign n15702 = n3818 & n32478 ;
  assign n15703 = n15701 | n15702 ;
  assign n15704 = n13232 | n15703 ;
  assign n15705 = x26 | n15704 ;
  assign n15706 = x26 & n15704 ;
  assign n33014 = ~n15706 ;
  assign n15707 = n15705 & n33014 ;
  assign n33015 = ~n15707 ;
  assign n15709 = n15700 & n33015 ;
  assign n33016 = ~n15700 ;
  assign n15708 = n33016 & n15707 ;
  assign n15710 = n15708 | n15709 ;
  assign n33017 = ~n14836 ;
  assign n15711 = n33017 & n14901 ;
  assign n15712 = n14902 | n15711 ;
  assign n13283 = n3791 & n32482 ;
  assign n10804 = n3802 & n31998 ;
  assign n10825 = n209 & n10818 ;
  assign n15713 = n10804 | n10825 ;
  assign n15714 = n3818 & n13292 ;
  assign n15715 = n15713 | n15714 ;
  assign n15716 = n13283 | n15715 ;
  assign n15717 = x26 | n15716 ;
  assign n15718 = x26 & n15716 ;
  assign n33018 = ~n15718 ;
  assign n15719 = n15717 & n33018 ;
  assign n15721 = n15712 | n15719 ;
  assign n15720 = n15712 & n15719 ;
  assign n33019 = ~n15720 ;
  assign n15722 = n33019 & n15721 ;
  assign n13321 = n3791 & n32488 ;
  assign n10822 = n3802 & n10818 ;
  assign n10850 = n209 & n10841 ;
  assign n15723 = n10822 | n10850 ;
  assign n15724 = n3818 & n31998 ;
  assign n15725 = n15723 | n15724 ;
  assign n15726 = n13321 | n15725 ;
  assign n15727 = x26 | n15726 ;
  assign n15728 = x26 & n15726 ;
  assign n33020 = ~n15728 ;
  assign n15729 = n15727 & n33020 ;
  assign n33021 = ~n14897 ;
  assign n15730 = n33021 & n14899 ;
  assign n15731 = n14900 | n15730 ;
  assign n33022 = ~n15729 ;
  assign n15733 = n33022 & n15731 ;
  assign n33023 = ~n15731 ;
  assign n15732 = n15729 & n33023 ;
  assign n15734 = n15732 | n15733 ;
  assign n15735 = n14894 & n14895 ;
  assign n33024 = ~n15735 ;
  assign n15736 = n14896 & n33024 ;
  assign n13385 = n3791 & n13382 ;
  assign n10848 = n3802 & n10841 ;
  assign n10873 = n209 & n10865 ;
  assign n15737 = n10848 | n10873 ;
  assign n15738 = n3818 & n10818 ;
  assign n15739 = n15737 | n15738 ;
  assign n15740 = n13385 | n15739 ;
  assign n15741 = x26 | n15740 ;
  assign n15742 = x26 & n15740 ;
  assign n33025 = ~n15742 ;
  assign n15743 = n15741 & n33025 ;
  assign n33026 = ~n15743 ;
  assign n15745 = n15736 & n33026 ;
  assign n33027 = ~n15736 ;
  assign n15744 = n33027 & n15743 ;
  assign n15746 = n15744 | n15745 ;
  assign n14885 = n14883 & n14884 ;
  assign n33028 = ~n14885 ;
  assign n15747 = n33028 & n14886 ;
  assign n33029 = ~n14893 ;
  assign n15748 = n33029 & n15747 ;
  assign n33030 = ~n15747 ;
  assign n15749 = n14893 & n33030 ;
  assign n15750 = n15748 | n15749 ;
  assign n13460 = n3791 & n13456 ;
  assign n10870 = n3802 & n10865 ;
  assign n10897 = n209 & n10892 ;
  assign n15751 = n10870 | n10897 ;
  assign n15752 = n3818 & n10841 ;
  assign n15753 = n15751 | n15752 ;
  assign n15754 = n13460 | n15753 ;
  assign n15755 = x26 | n15754 ;
  assign n15756 = x26 & n15754 ;
  assign n33031 = ~n15756 ;
  assign n15757 = n15755 & n33031 ;
  assign n15759 = n15750 | n15757 ;
  assign n33032 = ~n15750 ;
  assign n15758 = n33032 & n15757 ;
  assign n33033 = ~n15757 ;
  assign n15760 = n15750 & n33033 ;
  assign n15761 = n15758 | n15760 ;
  assign n14881 = n14874 & n14880 ;
  assign n33034 = ~n14881 ;
  assign n15762 = n33034 & n14882 ;
  assign n13529 = n3791 & n32502 ;
  assign n10907 = n3802 & n10892 ;
  assign n10924 = n209 & n32503 ;
  assign n15763 = n10907 | n10924 ;
  assign n15764 = n3818 & n10865 ;
  assign n15765 = n15763 | n15764 ;
  assign n15766 = n13529 | n15765 ;
  assign n15767 = x26 | n15766 ;
  assign n15768 = x26 & n15766 ;
  assign n33035 = ~n15768 ;
  assign n15769 = n15767 & n33035 ;
  assign n15770 = n15762 & n15769 ;
  assign n15771 = x29 & n14858 ;
  assign n33036 = ~n14872 ;
  assign n15772 = n33036 & n15771 ;
  assign n33037 = ~n15771 ;
  assign n15773 = n14872 & n33037 ;
  assign n15774 = n15772 | n15773 ;
  assign n13760 = n3791 & n13756 ;
  assign n10926 = n3802 & n32503 ;
  assign n10967 = n209 & n10940 ;
  assign n15775 = n10926 | n10967 ;
  assign n15776 = n3818 & n10892 ;
  assign n15777 = n15775 | n15776 ;
  assign n15778 = n13760 | n15777 ;
  assign n15779 = x26 | n15778 ;
  assign n15780 = x26 & n15778 ;
  assign n33038 = ~n15780 ;
  assign n15781 = n15779 & n33038 ;
  assign n15783 = n15774 | n15781 ;
  assign n15784 = n260 & n32507 ;
  assign n15785 = x26 & n15784 ;
  assign n14862 = n3791 & n14859 ;
  assign n15786 = n3818 & n31995 ;
  assign n15787 = n3802 & n32507 ;
  assign n15788 = n15786 | n15787 ;
  assign n15789 = n14862 | n15788 ;
  assign n15791 = n15785 | n15789 ;
  assign n15792 = x26 & n15791 ;
  assign n10966 = n3818 & n10940 ;
  assign n15793 = n3802 & n31995 ;
  assign n15794 = n209 & n32507 ;
  assign n15795 = n15793 | n15794 ;
  assign n15796 = n10966 | n15795 ;
  assign n15797 = n3791 & n13637 ;
  assign n15798 = n15796 | n15797 ;
  assign n15800 = n15792 | n15798 ;
  assign n33039 = ~n15800 ;
  assign n15801 = x26 & n33039 ;
  assign n15803 = n14858 | n15801 ;
  assign n13695 = n3791 & n13690 ;
  assign n10944 = n3802 & n10940 ;
  assign n10979 = n209 & n31995 ;
  assign n15804 = n10944 | n10979 ;
  assign n15805 = n3818 & n32503 ;
  assign n15806 = n15804 | n15805 ;
  assign n15807 = n13695 | n15806 ;
  assign n33040 = ~n15807 ;
  assign n15808 = x26 & n33040 ;
  assign n15809 = n30019 & n15807 ;
  assign n15810 = n15808 | n15809 ;
  assign n15811 = n15803 & n15810 ;
  assign n15782 = n15774 & n15781 ;
  assign n33041 = ~n15782 ;
  assign n15812 = n33041 & n15783 ;
  assign n33042 = ~n15811 ;
  assign n15813 = n33042 & n15812 ;
  assign n33043 = ~n15813 ;
  assign n15814 = n15783 & n33043 ;
  assign n15815 = n15762 | n15769 ;
  assign n33044 = ~n15770 ;
  assign n15816 = n33044 & n15815 ;
  assign n15817 = n15814 & n15816 ;
  assign n15818 = n15770 | n15817 ;
  assign n33045 = ~n15818 ;
  assign n15819 = n15761 & n33045 ;
  assign n33046 = ~n15819 ;
  assign n15820 = n15759 & n33046 ;
  assign n15822 = n15746 | n15820 ;
  assign n33047 = ~n15745 ;
  assign n15823 = n33047 & n15822 ;
  assign n15825 = n15734 | n15823 ;
  assign n33048 = ~n15733 ;
  assign n15826 = n33048 & n15825 ;
  assign n33049 = ~n15826 ;
  assign n15828 = n15722 & n33049 ;
  assign n33050 = ~n15828 ;
  assign n15829 = n15721 & n33050 ;
  assign n15831 = n15710 | n15829 ;
  assign n33051 = ~n15709 ;
  assign n15832 = n33051 & n15831 ;
  assign n33052 = ~n15698 ;
  assign n15833 = n33052 & n15832 ;
  assign n15834 = n15696 | n15833 ;
  assign n33053 = ~n15834 ;
  assign n15835 = n15685 & n33053 ;
  assign n33054 = ~n15835 ;
  assign n15836 = n15683 & n33054 ;
  assign n15671 = n15663 & n15670 ;
  assign n33055 = ~n15671 ;
  assign n15837 = n33055 & n15672 ;
  assign n33056 = ~n15836 ;
  assign n15839 = n33056 & n15837 ;
  assign n33057 = ~n15839 ;
  assign n15840 = n15672 & n33057 ;
  assign n15841 = n15661 & n15840 ;
  assign n15842 = n15659 | n15841 ;
  assign n33058 = ~n15842 ;
  assign n15843 = n15648 & n33058 ;
  assign n33059 = ~n15843 ;
  assign n15844 = n15646 & n33059 ;
  assign n33060 = ~n15844 ;
  assign n15846 = n15635 & n33060 ;
  assign n33061 = ~n15846 ;
  assign n15847 = n15633 & n33061 ;
  assign n15849 = n15622 | n15847 ;
  assign n33062 = ~n15621 ;
  assign n15850 = n33062 & n15849 ;
  assign n15609 = n15601 & n15608 ;
  assign n33063 = ~n15609 ;
  assign n15851 = n33063 & n15610 ;
  assign n33064 = ~n15850 ;
  assign n15852 = n33064 & n15851 ;
  assign n33065 = ~n15852 ;
  assign n15853 = n15610 & n33065 ;
  assign n15855 = n15599 | n15853 ;
  assign n33066 = ~n15598 ;
  assign n15856 = n33066 & n15855 ;
  assign n15858 = n15587 | n15856 ;
  assign n33067 = ~n15585 ;
  assign n15859 = n33067 & n15858 ;
  assign n15861 = n15574 | n15859 ;
  assign n15291 = n5937 & n15288 ;
  assign n14499 = n5970 & n32707 ;
  assign n14524 = n5994 & n32706 ;
  assign n15862 = n14499 | n14524 ;
  assign n15863 = n6018 & n15081 ;
  assign n15864 = n15862 | n15863 ;
  assign n15865 = n15291 | n15864 ;
  assign n33068 = ~n15865 ;
  assign n15866 = x14 & n33068 ;
  assign n15867 = n30547 & n15865 ;
  assign n15868 = n15866 | n15867 ;
  assign n33069 = ~n15574 ;
  assign n15860 = n33069 & n15859 ;
  assign n33070 = ~n15859 ;
  assign n15869 = n15574 & n33070 ;
  assign n15870 = n15860 | n15869 ;
  assign n33071 = ~n15868 ;
  assign n15871 = n33071 & n15870 ;
  assign n33072 = ~n15871 ;
  assign n15872 = n15861 & n33072 ;
  assign n15874 = n15572 | n15872 ;
  assign n33073 = ~n15130 ;
  assign n15875 = n33073 & n15132 ;
  assign n15876 = n15133 | n15875 ;
  assign n15873 = n15572 & n15872 ;
  assign n33074 = ~n15873 ;
  assign n15877 = n33074 & n15874 ;
  assign n15878 = n15876 & n15877 ;
  assign n33075 = ~n15878 ;
  assign n15879 = n15874 & n33075 ;
  assign n33076 = ~n15879 ;
  assign n15881 = n15565 & n33076 ;
  assign n15517 = n6188 & n15516 ;
  assign n15228 = n6190 & n15221 ;
  assign n15882 = n6217 | n15228 ;
  assign n15883 = n6244 & n32890 ;
  assign n15884 = n15882 | n15883 ;
  assign n15885 = n15517 | n15884 ;
  assign n33077 = ~n15885 ;
  assign n15886 = x11 & n33077 ;
  assign n15887 = n30180 & n15885 ;
  assign n15888 = n15886 | n15887 ;
  assign n33078 = ~n15565 ;
  assign n15880 = n33078 & n15879 ;
  assign n15889 = n15880 | n15881 ;
  assign n15890 = n15888 | n15889 ;
  assign n33079 = ~n15881 ;
  assign n15891 = n33079 & n15890 ;
  assign n33080 = ~n15891 ;
  assign n15893 = n15563 & n33080 ;
  assign n33081 = ~n15563 ;
  assign n15892 = n33081 & n15891 ;
  assign n15894 = n15892 | n15893 ;
  assign n15895 = n15888 & n15889 ;
  assign n33082 = ~n15895 ;
  assign n15896 = n15890 & n33082 ;
  assign n15267 = n6272 & n32889 ;
  assign n15061 = n6244 & n32856 ;
  assign n15173 = n6190 & n32876 ;
  assign n15897 = n15061 | n15173 ;
  assign n15898 = n6217 & n32890 ;
  assign n15899 = n15897 | n15898 ;
  assign n15900 = n15267 | n15899 ;
  assign n15901 = x11 | n15900 ;
  assign n15902 = x11 & n15900 ;
  assign n33083 = ~n15902 ;
  assign n15903 = n15901 & n33083 ;
  assign n33084 = ~n15870 ;
  assign n15904 = n15868 & n33084 ;
  assign n15905 = n15871 | n15904 ;
  assign n15907 = n15903 | n15905 ;
  assign n33085 = ~n15587 ;
  assign n15857 = n33085 & n15856 ;
  assign n33086 = ~n15856 ;
  assign n15908 = n15587 & n33086 ;
  assign n15909 = n15857 | n15908 ;
  assign n14573 = n5937 & n14570 ;
  assign n14521 = n5970 & n32706 ;
  assign n14550 = n5994 & n14536 ;
  assign n15910 = n14521 | n14550 ;
  assign n15911 = n6018 & n32707 ;
  assign n15912 = n15910 | n15911 ;
  assign n15913 = n14573 | n15912 ;
  assign n15914 = x14 | n15913 ;
  assign n15915 = x14 & n15913 ;
  assign n33087 = ~n15915 ;
  assign n15916 = n15914 & n33087 ;
  assign n33088 = ~n15916 ;
  assign n15918 = n15909 & n33088 ;
  assign n15917 = n15909 & n15916 ;
  assign n15919 = n15909 | n15916 ;
  assign n33089 = ~n15917 ;
  assign n15920 = n33089 & n15919 ;
  assign n33090 = ~n15599 ;
  assign n15854 = n33090 & n15853 ;
  assign n33091 = ~n15853 ;
  assign n15921 = n15599 & n33091 ;
  assign n15922 = n15854 | n15921 ;
  assign n14687 = n5937 & n32735 ;
  assign n14107 = n5994 & n14101 ;
  assign n14548 = n5970 & n14536 ;
  assign n15923 = n14107 | n14548 ;
  assign n15924 = n6018 & n32706 ;
  assign n15925 = n15923 | n15924 ;
  assign n15926 = n14687 | n15925 ;
  assign n15927 = x14 | n15926 ;
  assign n15928 = x14 & n15926 ;
  assign n33092 = ~n15928 ;
  assign n15929 = n15927 & n33092 ;
  assign n33093 = ~n15929 ;
  assign n15931 = n15922 & n33093 ;
  assign n33094 = ~n15851 ;
  assign n15932 = n15850 & n33094 ;
  assign n15933 = n15852 | n15932 ;
  assign n14660 = n37300 & n14655 ;
  assign n13034 = n5144 & n13027 ;
  assign n13066 = n5166 & n32456 ;
  assign n15934 = n13034 | n13066 ;
  assign n15935 = n5191 & n14147 ;
  assign n15936 = n15934 | n15935 ;
  assign n15937 = n14660 | n15936 ;
  assign n15938 = x17 | n15937 ;
  assign n15939 = x17 & n15937 ;
  assign n33095 = ~n15939 ;
  assign n15940 = n15938 & n33095 ;
  assign n15942 = n15933 | n15940 ;
  assign n33096 = ~n15622 ;
  assign n15848 = n33096 & n15847 ;
  assign n33097 = ~n15847 ;
  assign n15943 = n15622 & n33097 ;
  assign n15944 = n15848 | n15943 ;
  assign n12633 = n4686 & n32356 ;
  assign n12572 = n4706 & n12570 ;
  assign n12601 = n4726 & n12595 ;
  assign n15945 = n12572 | n12601 ;
  assign n15946 = n4748 & n32354 ;
  assign n15947 = n15945 | n15946 ;
  assign n15948 = n12633 | n15947 ;
  assign n15949 = x20 | n15948 ;
  assign n15950 = x20 & n15948 ;
  assign n33098 = ~n15950 ;
  assign n15951 = n15949 & n33098 ;
  assign n33099 = ~n15951 ;
  assign n15953 = n15944 & n33099 ;
  assign n15952 = n15944 & n15951 ;
  assign n15954 = n15944 | n15951 ;
  assign n33100 = ~n15952 ;
  assign n15955 = n33100 & n15954 ;
  assign n15845 = n15635 & n15844 ;
  assign n15956 = n15635 | n15844 ;
  assign n33101 = ~n15845 ;
  assign n15957 = n33101 & n15956 ;
  assign n12659 = n4135 & n32362 ;
  assign n11436 = n4185 & n11430 ;
  assign n11844 = n4148 & n32176 ;
  assign n15958 = n11436 | n11844 ;
  assign n15959 = n4165 & n12161 ;
  assign n15960 = n15958 | n15959 ;
  assign n15961 = n12659 | n15960 ;
  assign n15962 = x23 | n15961 ;
  assign n15963 = x23 & n15961 ;
  assign n33102 = ~n15963 ;
  assign n15964 = n15962 & n33102 ;
  assign n15966 = n15957 | n15964 ;
  assign n33103 = ~n15957 ;
  assign n15965 = n33103 & n15964 ;
  assign n33104 = ~n15964 ;
  assign n15967 = n15957 & n33104 ;
  assign n15968 = n15965 | n15967 ;
  assign n33105 = ~n15648 ;
  assign n15969 = n33105 & n15842 ;
  assign n15970 = n15843 | n15969 ;
  assign n11875 = n4135 & n32178 ;
  assign n11432 = n4148 & n11430 ;
  assign n11479 = n4185 & n11476 ;
  assign n15971 = n11432 | n11479 ;
  assign n15972 = n4165 & n32176 ;
  assign n15973 = n15971 | n15972 ;
  assign n15974 = n11875 | n15973 ;
  assign n15975 = x23 | n15974 ;
  assign n15976 = x23 & n15974 ;
  assign n33106 = ~n15976 ;
  assign n15977 = n15975 & n33106 ;
  assign n15979 = n15970 | n15977 ;
  assign n33107 = ~n15970 ;
  assign n15978 = n33107 & n15977 ;
  assign n33108 = ~n15977 ;
  assign n15980 = n15970 & n33108 ;
  assign n15981 = n15978 | n15980 ;
  assign n15982 = n15661 | n15840 ;
  assign n33109 = ~n15841 ;
  assign n15983 = n33109 & n15982 ;
  assign n11470 = n4135 & n11463 ;
  assign n10663 = n4185 & n10656 ;
  assign n11480 = n4148 & n11476 ;
  assign n15984 = n10663 | n11480 ;
  assign n15985 = n4165 & n11430 ;
  assign n15986 = n15984 | n15985 ;
  assign n15987 = n11470 | n15986 ;
  assign n15988 = x23 | n15987 ;
  assign n15989 = x23 & n15987 ;
  assign n33110 = ~n15989 ;
  assign n15990 = n15988 & n33110 ;
  assign n15992 = n15983 | n15990 ;
  assign n15991 = n15983 & n15990 ;
  assign n33111 = ~n15991 ;
  assign n15993 = n33111 & n15992 ;
  assign n15838 = n15836 & n15837 ;
  assign n15994 = n15836 | n15837 ;
  assign n33112 = ~n15838 ;
  assign n15995 = n33112 & n15994 ;
  assign n11516 = n4135 & n11511 ;
  assign n10661 = n4148 & n10656 ;
  assign n11049 = n4185 & n10679 ;
  assign n15996 = n10661 | n11049 ;
  assign n15997 = n4165 & n11452 ;
  assign n15998 = n15996 | n15997 ;
  assign n15999 = n11516 | n15998 ;
  assign n16000 = x23 | n15999 ;
  assign n16001 = x23 & n15999 ;
  assign n33113 = ~n16001 ;
  assign n16002 = n16000 & n33113 ;
  assign n16004 = n15995 | n16002 ;
  assign n33114 = ~n15995 ;
  assign n16003 = n33114 & n16002 ;
  assign n33115 = ~n16002 ;
  assign n16005 = n15995 & n33115 ;
  assign n16006 = n16003 | n16005 ;
  assign n33116 = ~n15685 ;
  assign n16007 = n33116 & n15834 ;
  assign n16008 = n15835 | n16007 ;
  assign n11034 = n4135 & n11030 ;
  assign n10685 = n4185 & n10681 ;
  assign n11047 = n4148 & n10679 ;
  assign n16009 = n10685 | n11047 ;
  assign n16010 = n4165 & n10656 ;
  assign n16011 = n16009 | n16010 ;
  assign n16012 = n11034 | n16011 ;
  assign n16013 = x23 | n16012 ;
  assign n16014 = x23 & n16012 ;
  assign n33117 = ~n16014 ;
  assign n16015 = n16013 & n33117 ;
  assign n16017 = n16008 | n16015 ;
  assign n33118 = ~n16008 ;
  assign n16016 = n33118 & n16015 ;
  assign n33119 = ~n16015 ;
  assign n16018 = n16008 & n33119 ;
  assign n16019 = n16016 | n16018 ;
  assign n33120 = ~n15832 ;
  assign n16020 = n15698 & n33120 ;
  assign n16021 = n15833 | n16020 ;
  assign n11540 = n4135 & n11536 ;
  assign n10682 = n4148 & n10681 ;
  assign n10712 = n4185 & n10703 ;
  assign n16022 = n10682 | n10712 ;
  assign n16023 = n4165 & n10679 ;
  assign n16024 = n16022 | n16023 ;
  assign n16025 = n11540 | n16024 ;
  assign n16026 = x23 | n16025 ;
  assign n16027 = x23 & n16025 ;
  assign n33121 = ~n16027 ;
  assign n16028 = n16026 & n33121 ;
  assign n33122 = ~n16028 ;
  assign n16030 = n16021 & n33122 ;
  assign n33123 = ~n16021 ;
  assign n16029 = n33123 & n16028 ;
  assign n16031 = n16029 | n16030 ;
  assign n33124 = ~n15710 ;
  assign n15830 = n33124 & n15829 ;
  assign n33125 = ~n15829 ;
  assign n16032 = n15710 & n33125 ;
  assign n16033 = n15830 | n16032 ;
  assign n13162 = n4135 & n13157 ;
  assign n10710 = n4148 & n10703 ;
  assign n10729 = n4185 & n10727 ;
  assign n16034 = n10710 | n10729 ;
  assign n16035 = n4165 & n10681 ;
  assign n16036 = n16034 | n16035 ;
  assign n16037 = n13162 | n16036 ;
  assign n16038 = x23 | n16037 ;
  assign n16039 = x23 & n16037 ;
  assign n33126 = ~n16039 ;
  assign n16040 = n16038 & n33126 ;
  assign n33127 = ~n16040 ;
  assign n16042 = n16033 & n33127 ;
  assign n16041 = n16033 & n16040 ;
  assign n16043 = n16033 | n16040 ;
  assign n33128 = ~n16041 ;
  assign n16044 = n33128 & n16043 ;
  assign n15827 = n15722 & n15826 ;
  assign n16045 = n15722 | n15826 ;
  assign n33129 = ~n15827 ;
  assign n16046 = n33129 & n16045 ;
  assign n13190 = n4135 & n13182 ;
  assign n10731 = n4148 & n10727 ;
  assign n10757 = n4185 & n31999 ;
  assign n16047 = n10731 | n10757 ;
  assign n16048 = n4165 & n13151 ;
  assign n16049 = n16047 | n16048 ;
  assign n16050 = n13190 | n16049 ;
  assign n33130 = ~n16050 ;
  assign n16051 = x23 & n33130 ;
  assign n16052 = n30030 & n16050 ;
  assign n16053 = n16051 | n16052 ;
  assign n16054 = n16046 | n16053 ;
  assign n16055 = n16046 & n16053 ;
  assign n33131 = ~n16055 ;
  assign n16056 = n16054 & n33131 ;
  assign n33132 = ~n15734 ;
  assign n15824 = n33132 & n15823 ;
  assign n33133 = ~n15823 ;
  assign n16057 = n15734 & n33133 ;
  assign n16058 = n15824 | n16057 ;
  assign n11690 = n4135 & n32125 ;
  assign n10758 = n4148 & n31999 ;
  assign n10777 = n4185 & n10773 ;
  assign n16059 = n10758 | n10777 ;
  assign n16060 = n4165 & n10727 ;
  assign n16061 = n16059 | n16060 ;
  assign n16062 = n11690 | n16061 ;
  assign n16063 = x23 | n16062 ;
  assign n16064 = x23 & n16062 ;
  assign n33134 = ~n16064 ;
  assign n16065 = n16063 & n33134 ;
  assign n33135 = ~n16065 ;
  assign n16067 = n16058 & n33135 ;
  assign n33136 = ~n16058 ;
  assign n16066 = n33136 & n16065 ;
  assign n16068 = n16066 | n16067 ;
  assign n33137 = ~n15746 ;
  assign n15821 = n33137 & n15820 ;
  assign n33138 = ~n15820 ;
  assign n16069 = n15746 & n33138 ;
  assign n16070 = n15821 | n16069 ;
  assign n13234 = n4135 & n32477 ;
  assign n10774 = n4148 & n10773 ;
  assign n10802 = n4185 & n31998 ;
  assign n16071 = n10774 | n10802 ;
  assign n16072 = n4165 & n32478 ;
  assign n16073 = n16071 | n16072 ;
  assign n16074 = n13234 | n16073 ;
  assign n16075 = x23 | n16074 ;
  assign n16076 = x23 & n16074 ;
  assign n33139 = ~n16076 ;
  assign n16077 = n16075 & n33139 ;
  assign n33140 = ~n16077 ;
  assign n16079 = n16070 & n33140 ;
  assign n33141 = ~n16070 ;
  assign n16078 = n33141 & n16077 ;
  assign n16080 = n16078 | n16079 ;
  assign n33142 = ~n15761 ;
  assign n16081 = n33142 & n15818 ;
  assign n16082 = n15819 | n16081 ;
  assign n13284 = n4135 & n32482 ;
  assign n10803 = n4148 & n31998 ;
  assign n10821 = n4185 & n10818 ;
  assign n16083 = n10803 | n10821 ;
  assign n16084 = n4165 & n13292 ;
  assign n16085 = n16083 | n16084 ;
  assign n16086 = n13284 | n16085 ;
  assign n16087 = x23 | n16086 ;
  assign n16088 = x23 & n16086 ;
  assign n33143 = ~n16088 ;
  assign n16089 = n16087 & n33143 ;
  assign n16091 = n16082 | n16089 ;
  assign n16090 = n16082 & n16089 ;
  assign n33144 = ~n16090 ;
  assign n16092 = n33144 & n16091 ;
  assign n13322 = n4135 & n32488 ;
  assign n10829 = n4148 & n10818 ;
  assign n10852 = n4185 & n10841 ;
  assign n16093 = n10829 | n10852 ;
  assign n16094 = n4165 & n31998 ;
  assign n16095 = n16093 | n16094 ;
  assign n16096 = n13322 | n16095 ;
  assign n16097 = x23 | n16096 ;
  assign n16098 = x23 & n16096 ;
  assign n33145 = ~n16098 ;
  assign n16099 = n16097 & n33145 ;
  assign n16100 = n15814 | n15816 ;
  assign n33146 = ~n15817 ;
  assign n16101 = n33146 & n16100 ;
  assign n16103 = n16099 | n16101 ;
  assign n16102 = n16099 & n16101 ;
  assign n33147 = ~n16102 ;
  assign n16104 = n33147 & n16103 ;
  assign n13388 = n4135 & n13382 ;
  assign n10846 = n4148 & n10841 ;
  assign n10869 = n4185 & n10865 ;
  assign n16105 = n10846 | n10869 ;
  assign n16106 = n4165 & n10818 ;
  assign n16107 = n16105 | n16106 ;
  assign n16108 = n13388 | n16107 ;
  assign n16109 = x23 | n16108 ;
  assign n16110 = x23 & n16108 ;
  assign n33148 = ~n16110 ;
  assign n16111 = n16109 & n33148 ;
  assign n33149 = ~n15812 ;
  assign n16112 = n15811 & n33149 ;
  assign n16113 = n15813 | n16112 ;
  assign n16115 = n16111 | n16113 ;
  assign n33150 = ~n16113 ;
  assign n16114 = n16111 & n33150 ;
  assign n33151 = ~n16111 ;
  assign n16116 = n33151 & n16113 ;
  assign n16117 = n16114 | n16116 ;
  assign n33152 = ~n14858 ;
  assign n15802 = n33152 & n15801 ;
  assign n33153 = ~n15801 ;
  assign n16118 = n14858 & n33153 ;
  assign n16119 = n15802 | n16118 ;
  assign n33154 = ~n15810 ;
  assign n16120 = n33154 & n16119 ;
  assign n33155 = ~n16119 ;
  assign n16121 = n15810 & n33155 ;
  assign n16122 = n16120 | n16121 ;
  assign n13462 = n4135 & n13456 ;
  assign n10868 = n4148 & n10865 ;
  assign n10906 = n4185 & n10892 ;
  assign n16123 = n10868 | n10906 ;
  assign n16124 = n4165 & n10841 ;
  assign n16125 = n16123 | n16124 ;
  assign n16126 = n13462 | n16125 ;
  assign n33156 = ~n16126 ;
  assign n16127 = x23 & n33156 ;
  assign n16128 = n30030 & n16126 ;
  assign n16129 = n16127 | n16128 ;
  assign n16130 = n16122 | n16129 ;
  assign n16131 = n16122 & n16129 ;
  assign n33157 = ~n16131 ;
  assign n16132 = n16130 & n33157 ;
  assign n13532 = n4135 & n32502 ;
  assign n10904 = n4148 & n10892 ;
  assign n10922 = n4185 & n32503 ;
  assign n16133 = n10904 | n10922 ;
  assign n16134 = n4165 & n10865 ;
  assign n16135 = n16133 | n16134 ;
  assign n16136 = n13532 | n16135 ;
  assign n16137 = x23 | n16136 ;
  assign n16138 = x23 & n16136 ;
  assign n33158 = ~n16138 ;
  assign n16139 = n16137 & n33158 ;
  assign n33159 = ~n15792 ;
  assign n15799 = n33159 & n15798 ;
  assign n33160 = ~n15798 ;
  assign n16140 = n15792 & n33160 ;
  assign n16141 = n15799 | n16140 ;
  assign n16143 = n16139 | n16141 ;
  assign n16142 = n16139 & n16141 ;
  assign n33161 = ~n16142 ;
  assign n16144 = n33161 & n16143 ;
  assign n16145 = n4132 & n32507 ;
  assign n14863 = n4135 & n14859 ;
  assign n16146 = n4165 & n31995 ;
  assign n16147 = n4148 & n32507 ;
  assign n16148 = n16146 | n16147 ;
  assign n16149 = n14863 | n16148 ;
  assign n16150 = n16145 | n16149 ;
  assign n16151 = x23 & n16150 ;
  assign n10959 = n4165 & n10940 ;
  assign n16152 = n4148 & n31995 ;
  assign n16153 = n4185 & n32507 ;
  assign n16154 = n16152 | n16153 ;
  assign n16155 = n10959 | n16154 ;
  assign n16156 = n4135 & n13637 ;
  assign n16157 = n16155 | n16156 ;
  assign n16159 = n16151 | n16157 ;
  assign n33162 = ~n16159 ;
  assign n16160 = x23 & n33162 ;
  assign n16162 = n15784 | n16160 ;
  assign n13694 = n4135 & n13690 ;
  assign n10958 = n4148 & n10940 ;
  assign n10981 = n4185 & n31995 ;
  assign n16163 = n10958 | n10981 ;
  assign n16164 = n4165 & n32503 ;
  assign n16165 = n16163 | n16164 ;
  assign n16166 = n13694 | n16165 ;
  assign n33163 = ~n16166 ;
  assign n16167 = x23 & n33163 ;
  assign n16168 = n30030 & n16166 ;
  assign n16169 = n16167 | n16168 ;
  assign n16170 = n16162 & n16169 ;
  assign n33164 = ~n15789 ;
  assign n15790 = n15785 & n33164 ;
  assign n33165 = ~n15785 ;
  assign n16171 = n33165 & n15789 ;
  assign n16172 = n15790 | n16171 ;
  assign n16174 = n16170 | n16172 ;
  assign n13762 = n4135 & n13756 ;
  assign n10921 = n4148 & n32503 ;
  assign n10949 = n4185 & n10940 ;
  assign n16175 = n10921 | n10949 ;
  assign n16176 = n4165 & n10892 ;
  assign n16177 = n16175 | n16176 ;
  assign n16178 = n13762 | n16177 ;
  assign n33166 = ~n16178 ;
  assign n16179 = x23 & n33166 ;
  assign n16180 = n30030 & n16178 ;
  assign n16181 = n16179 | n16180 ;
  assign n16173 = n16170 & n16172 ;
  assign n33167 = ~n16173 ;
  assign n16182 = n33167 & n16174 ;
  assign n33168 = ~n16181 ;
  assign n16183 = n33168 & n16182 ;
  assign n33169 = ~n16183 ;
  assign n16184 = n16174 & n33169 ;
  assign n33170 = ~n16184 ;
  assign n16186 = n16144 & n33170 ;
  assign n33171 = ~n16186 ;
  assign n16187 = n16143 & n33171 ;
  assign n33172 = ~n16187 ;
  assign n16189 = n16132 & n33172 ;
  assign n33173 = ~n16189 ;
  assign n16190 = n16130 & n33173 ;
  assign n33174 = ~n16190 ;
  assign n16192 = n16117 & n33174 ;
  assign n33175 = ~n16192 ;
  assign n16193 = n16115 & n33175 ;
  assign n33176 = ~n16193 ;
  assign n16195 = n16104 & n33176 ;
  assign n33177 = ~n16195 ;
  assign n16196 = n16103 & n33177 ;
  assign n33178 = ~n16196 ;
  assign n16198 = n16092 & n33178 ;
  assign n33179 = ~n16198 ;
  assign n16199 = n16091 & n33179 ;
  assign n16201 = n16080 | n16199 ;
  assign n33180 = ~n16079 ;
  assign n16202 = n33180 & n16201 ;
  assign n16204 = n16068 | n16202 ;
  assign n33181 = ~n16067 ;
  assign n16205 = n33181 & n16204 ;
  assign n33182 = ~n16205 ;
  assign n16207 = n16056 & n33182 ;
  assign n33183 = ~n16207 ;
  assign n16208 = n16054 & n33183 ;
  assign n16210 = n16044 | n16208 ;
  assign n33184 = ~n16042 ;
  assign n16211 = n33184 & n16210 ;
  assign n16213 = n16031 | n16211 ;
  assign n33185 = ~n16030 ;
  assign n16214 = n33185 & n16213 ;
  assign n33186 = ~n16214 ;
  assign n16216 = n16019 & n33186 ;
  assign n33187 = ~n16216 ;
  assign n16217 = n16017 & n33187 ;
  assign n33188 = ~n16217 ;
  assign n16219 = n16006 & n33188 ;
  assign n33189 = ~n16219 ;
  assign n16220 = n16004 & n33189 ;
  assign n33190 = ~n16220 ;
  assign n16222 = n15993 & n33190 ;
  assign n33191 = ~n16222 ;
  assign n16223 = n15992 & n33191 ;
  assign n33192 = ~n16223 ;
  assign n16225 = n15981 & n33192 ;
  assign n33193 = ~n16225 ;
  assign n16226 = n15979 & n33193 ;
  assign n33194 = ~n16226 ;
  assign n16228 = n15968 & n33194 ;
  assign n33195 = ~n16228 ;
  assign n16229 = n15966 & n33195 ;
  assign n16231 = n15955 | n16229 ;
  assign n33196 = ~n15953 ;
  assign n16232 = n33196 & n16231 ;
  assign n33197 = ~n15933 ;
  assign n15941 = n33197 & n15940 ;
  assign n33198 = ~n15940 ;
  assign n16233 = n15933 & n33198 ;
  assign n16234 = n15941 | n16233 ;
  assign n33199 = ~n16232 ;
  assign n16236 = n33199 & n16234 ;
  assign n33200 = ~n16236 ;
  assign n16237 = n15942 & n33200 ;
  assign n33201 = ~n15922 ;
  assign n15930 = n33201 & n15929 ;
  assign n16238 = n15930 | n15931 ;
  assign n16239 = n16237 | n16238 ;
  assign n33202 = ~n15931 ;
  assign n16240 = n33202 & n16239 ;
  assign n16242 = n15920 | n16240 ;
  assign n33203 = ~n15918 ;
  assign n16243 = n33203 & n16242 ;
  assign n33204 = ~n15905 ;
  assign n15906 = n15903 & n33204 ;
  assign n33205 = ~n15903 ;
  assign n16244 = n33205 & n15905 ;
  assign n16245 = n15906 | n16244 ;
  assign n33206 = ~n16243 ;
  assign n16246 = n33206 & n16245 ;
  assign n33207 = ~n16246 ;
  assign n16248 = n15907 & n33207 ;
  assign n16250 = n72 & n16248 ;
  assign n16251 = n15876 | n15877 ;
  assign n16252 = n33075 & n16251 ;
  assign n16249 = n30040 & n16248 ;
  assign n33208 = ~n16248 ;
  assign n16253 = n72 & n33208 ;
  assign n16254 = n16249 | n16253 ;
  assign n33209 = ~n16252 ;
  assign n16256 = n33209 & n16254 ;
  assign n16257 = n16250 | n16256 ;
  assign n33210 = ~n16257 ;
  assign n16258 = n15896 & n33210 ;
  assign n33211 = ~n15896 ;
  assign n16259 = n33211 & n16257 ;
  assign n16260 = n16258 | n16259 ;
  assign n16255 = n16252 & n16254 ;
  assign n16261 = n16252 | n16254 ;
  assign n33212 = ~n16255 ;
  assign n16262 = n33212 & n16261 ;
  assign n33213 = ~n15920 ;
  assign n16241 = n33213 & n16240 ;
  assign n33214 = ~n16240 ;
  assign n16263 = n15920 & n33214 ;
  assign n16264 = n16241 | n16263 ;
  assign n15187 = n6272 & n32875 ;
  assign n15067 = n6190 & n32856 ;
  assign n15098 = n6244 & n15081 ;
  assign n16265 = n15067 | n15098 ;
  assign n16266 = n6217 & n32876 ;
  assign n16267 = n16265 | n16266 ;
  assign n16268 = n15187 | n16267 ;
  assign n16269 = x11 | n16268 ;
  assign n16270 = x11 & n16268 ;
  assign n33215 = ~n16270 ;
  assign n16271 = n16269 & n33215 ;
  assign n33216 = ~n16271 ;
  assign n16273 = n16264 & n33216 ;
  assign n16272 = n16264 & n16271 ;
  assign n16274 = n16264 | n16271 ;
  assign n33217 = ~n16272 ;
  assign n16275 = n33217 & n16274 ;
  assign n16276 = n16237 & n16238 ;
  assign n33218 = ~n16276 ;
  assign n16277 = n16239 & n33218 ;
  assign n15115 = n6272 & n15111 ;
  assign n14498 = n6244 & n32707 ;
  assign n15096 = n6190 & n15081 ;
  assign n16278 = n14498 | n15096 ;
  assign n16279 = n6217 & n32856 ;
  assign n16280 = n16278 | n16279 ;
  assign n16281 = n15115 | n16280 ;
  assign n16282 = x11 | n16281 ;
  assign n16283 = x11 & n16281 ;
  assign n33219 = ~n16283 ;
  assign n16284 = n16282 & n33219 ;
  assign n33220 = ~n16284 ;
  assign n16286 = n16277 & n33220 ;
  assign n33221 = ~n16277 ;
  assign n16285 = n33221 & n16284 ;
  assign n16287 = n16285 | n16286 ;
  assign n16235 = n16232 & n16234 ;
  assign n16288 = n16232 | n16234 ;
  assign n33222 = ~n16235 ;
  assign n16289 = n33222 & n16288 ;
  assign n14970 = n5937 & n14965 ;
  assign n14104 = n5970 & n14101 ;
  assign n14131 = n5994 & n14124 ;
  assign n16290 = n14104 | n14131 ;
  assign n16291 = n6018 & n14536 ;
  assign n16292 = n16290 | n16291 ;
  assign n16293 = n14970 | n16292 ;
  assign n16294 = x14 | n16293 ;
  assign n16295 = x14 & n16293 ;
  assign n33223 = ~n16295 ;
  assign n16296 = n16294 & n33223 ;
  assign n16298 = n16289 | n16296 ;
  assign n16297 = n16289 & n16296 ;
  assign n33224 = ~n16297 ;
  assign n16299 = n33224 & n16298 ;
  assign n33225 = ~n15955 ;
  assign n16230 = n33225 & n16229 ;
  assign n33226 = ~n16229 ;
  assign n16300 = n15955 & n33226 ;
  assign n16301 = n16230 | n16300 ;
  assign n13119 = n37300 & n32455 ;
  assign n13058 = n5144 & n32456 ;
  assign n13079 = n5166 & n13077 ;
  assign n16302 = n13058 | n13079 ;
  assign n16303 = n5191 & n13027 ;
  assign n16304 = n16302 | n16303 ;
  assign n16305 = n13119 | n16304 ;
  assign n16306 = x17 | n16305 ;
  assign n16307 = x17 & n16305 ;
  assign n33227 = ~n16307 ;
  assign n16308 = n16306 & n33227 ;
  assign n33228 = ~n16308 ;
  assign n16310 = n16301 & n33228 ;
  assign n16227 = n15968 & n16226 ;
  assign n16311 = n15968 | n16226 ;
  assign n33229 = ~n16227 ;
  assign n16312 = n33229 & n16311 ;
  assign n12686 = n4686 & n12681 ;
  assign n12151 = n4726 & n32253 ;
  assign n12600 = n4706 & n12595 ;
  assign n16313 = n12151 | n12600 ;
  assign n16314 = n4748 & n12570 ;
  assign n16315 = n16313 | n16314 ;
  assign n16316 = n12686 | n16315 ;
  assign n16317 = x20 | n16316 ;
  assign n16318 = x20 & n16316 ;
  assign n33230 = ~n16318 ;
  assign n16319 = n16317 & n33230 ;
  assign n16321 = n16312 | n16319 ;
  assign n33231 = ~n16312 ;
  assign n16320 = n33231 & n16319 ;
  assign n33232 = ~n16319 ;
  assign n16322 = n16312 & n33232 ;
  assign n16323 = n16320 | n16322 ;
  assign n16224 = n15981 & n16223 ;
  assign n16324 = n15981 | n16223 ;
  assign n33233 = ~n16224 ;
  assign n16325 = n33233 & n16324 ;
  assign n13823 = n4686 & n32550 ;
  assign n12140 = n4706 & n32253 ;
  assign n12163 = n4726 & n12161 ;
  assign n16326 = n12140 | n12163 ;
  assign n16327 = n4748 & n12595 ;
  assign n16328 = n16326 | n16327 ;
  assign n16329 = n13823 | n16328 ;
  assign n16330 = x20 | n16329 ;
  assign n16331 = x20 & n16329 ;
  assign n33234 = ~n16331 ;
  assign n16332 = n16330 & n33234 ;
  assign n16334 = n16325 | n16332 ;
  assign n33235 = ~n16325 ;
  assign n16333 = n33235 & n16332 ;
  assign n33236 = ~n16332 ;
  assign n16335 = n16325 & n33236 ;
  assign n16336 = n16333 | n16335 ;
  assign n16221 = n15993 & n16220 ;
  assign n16337 = n15993 | n16220 ;
  assign n33237 = ~n16221 ;
  assign n16338 = n33237 & n16337 ;
  assign n12197 = n4686 & n32255 ;
  assign n11849 = n4726 & n32176 ;
  assign n12164 = n4706 & n12161 ;
  assign n16339 = n11849 | n12164 ;
  assign n16340 = n4748 & n32253 ;
  assign n16341 = n16339 | n16340 ;
  assign n16342 = n12197 | n16341 ;
  assign n16343 = x20 | n16342 ;
  assign n16344 = x20 & n16342 ;
  assign n33238 = ~n16344 ;
  assign n16345 = n16343 & n33238 ;
  assign n16347 = n16338 | n16345 ;
  assign n33239 = ~n16338 ;
  assign n16346 = n33239 & n16345 ;
  assign n33240 = ~n16345 ;
  assign n16348 = n16338 & n33240 ;
  assign n16349 = n16346 | n16348 ;
  assign n16218 = n16006 & n16217 ;
  assign n16350 = n16006 | n16217 ;
  assign n33241 = ~n16218 ;
  assign n16351 = n33241 & n16350 ;
  assign n12658 = n4686 & n32362 ;
  assign n11431 = n4726 & n11430 ;
  assign n11841 = n4706 & n32176 ;
  assign n16352 = n11431 | n11841 ;
  assign n16353 = n4748 & n12161 ;
  assign n16354 = n16352 | n16353 ;
  assign n16355 = n12658 | n16354 ;
  assign n16356 = x20 | n16355 ;
  assign n16357 = x20 & n16355 ;
  assign n33242 = ~n16357 ;
  assign n16358 = n16356 & n33242 ;
  assign n16360 = n16351 & n16358 ;
  assign n16215 = n16019 & n16214 ;
  assign n16361 = n16019 | n16214 ;
  assign n33243 = ~n16215 ;
  assign n16362 = n33243 & n16361 ;
  assign n11876 = n4686 & n32178 ;
  assign n11434 = n4706 & n11430 ;
  assign n11491 = n4726 & n11476 ;
  assign n16363 = n11434 | n11491 ;
  assign n16364 = n4748 & n32176 ;
  assign n16365 = n16363 | n16364 ;
  assign n16366 = n11876 | n16365 ;
  assign n16367 = x20 | n16366 ;
  assign n16368 = x20 & n16366 ;
  assign n33244 = ~n16368 ;
  assign n16369 = n16367 & n33244 ;
  assign n16371 = n16362 | n16369 ;
  assign n33245 = ~n16362 ;
  assign n16370 = n33245 & n16369 ;
  assign n33246 = ~n16369 ;
  assign n16372 = n16362 & n33246 ;
  assign n16373 = n16370 | n16372 ;
  assign n33247 = ~n16031 ;
  assign n16212 = n33247 & n16211 ;
  assign n33248 = ~n16211 ;
  assign n16374 = n16031 & n33248 ;
  assign n16375 = n16212 | n16374 ;
  assign n11471 = n4686 & n11463 ;
  assign n10657 = n4726 & n10656 ;
  assign n11477 = n4706 & n11476 ;
  assign n16376 = n10657 | n11477 ;
  assign n16377 = n4748 & n11430 ;
  assign n16378 = n16376 | n16377 ;
  assign n16379 = n11471 | n16378 ;
  assign n16380 = x20 | n16379 ;
  assign n16381 = x20 & n16379 ;
  assign n33249 = ~n16381 ;
  assign n16382 = n16380 & n33249 ;
  assign n33250 = ~n16382 ;
  assign n16384 = n16375 & n33250 ;
  assign n33251 = ~n16375 ;
  assign n16383 = n33251 & n16382 ;
  assign n16385 = n16383 | n16384 ;
  assign n33252 = ~n16044 ;
  assign n16209 = n33252 & n16208 ;
  assign n33253 = ~n16208 ;
  assign n16386 = n16044 & n33253 ;
  assign n16387 = n16209 | n16386 ;
  assign n11513 = n4686 & n11511 ;
  assign n10671 = n4706 & n10656 ;
  assign n11044 = n4726 & n10679 ;
  assign n16388 = n10671 | n11044 ;
  assign n16389 = n4748 & n11452 ;
  assign n16390 = n16388 | n16389 ;
  assign n16391 = n11513 | n16390 ;
  assign n16392 = x20 | n16391 ;
  assign n16393 = x20 & n16391 ;
  assign n33254 = ~n16393 ;
  assign n16394 = n16392 & n33254 ;
  assign n33255 = ~n16394 ;
  assign n16396 = n16387 & n33255 ;
  assign n16395 = n16387 & n16394 ;
  assign n16397 = n16387 | n16394 ;
  assign n33256 = ~n16395 ;
  assign n16398 = n33256 & n16397 ;
  assign n16206 = n16056 & n16205 ;
  assign n16399 = n16056 | n16205 ;
  assign n33257 = ~n16206 ;
  assign n16400 = n33257 & n16399 ;
  assign n11036 = n4686 & n11030 ;
  assign n10684 = n4726 & n10681 ;
  assign n11042 = n4706 & n10679 ;
  assign n16401 = n10684 | n11042 ;
  assign n16402 = n4748 & n10656 ;
  assign n16403 = n16401 | n16402 ;
  assign n16404 = n11036 | n16403 ;
  assign n16405 = x20 | n16404 ;
  assign n16406 = x20 & n16404 ;
  assign n33258 = ~n16406 ;
  assign n16407 = n16405 & n33258 ;
  assign n16409 = n16400 | n16407 ;
  assign n33259 = ~n16400 ;
  assign n16408 = n33259 & n16407 ;
  assign n33260 = ~n16407 ;
  assign n16410 = n16400 & n33260 ;
  assign n16411 = n16408 | n16410 ;
  assign n33261 = ~n16068 ;
  assign n16203 = n33261 & n16202 ;
  assign n33262 = ~n16202 ;
  assign n16412 = n16068 & n33262 ;
  assign n16413 = n16203 | n16412 ;
  assign n11541 = n4686 & n11536 ;
  assign n10693 = n4706 & n10681 ;
  assign n10708 = n4726 & n10703 ;
  assign n16414 = n10693 | n10708 ;
  assign n16415 = n4748 & n10679 ;
  assign n16416 = n16414 | n16415 ;
  assign n16417 = n11541 | n16416 ;
  assign n16418 = x20 | n16417 ;
  assign n16419 = x20 & n16417 ;
  assign n33263 = ~n16419 ;
  assign n16420 = n16418 & n33263 ;
  assign n33264 = ~n16420 ;
  assign n16422 = n16413 & n33264 ;
  assign n16421 = n16413 & n16420 ;
  assign n16423 = n16413 | n16420 ;
  assign n33265 = ~n16421 ;
  assign n16424 = n33265 & n16423 ;
  assign n33266 = ~n16080 ;
  assign n16200 = n33266 & n16199 ;
  assign n33267 = ~n16199 ;
  assign n16425 = n16080 & n33267 ;
  assign n16426 = n16200 | n16425 ;
  assign n13164 = n4686 & n13157 ;
  assign n10717 = n4706 & n10703 ;
  assign n10737 = n4726 & n10727 ;
  assign n16427 = n10717 | n10737 ;
  assign n16428 = n4748 & n10681 ;
  assign n16429 = n16427 | n16428 ;
  assign n16430 = n13164 | n16429 ;
  assign n16431 = x20 | n16430 ;
  assign n16432 = x20 & n16430 ;
  assign n33268 = ~n16432 ;
  assign n16433 = n16431 & n33268 ;
  assign n33269 = ~n16433 ;
  assign n16435 = n16426 & n33269 ;
  assign n16434 = n16426 & n16433 ;
  assign n16436 = n16426 | n16433 ;
  assign n33270 = ~n16434 ;
  assign n16437 = n33270 & n16436 ;
  assign n16197 = n16092 & n16196 ;
  assign n16438 = n16092 | n16196 ;
  assign n33271 = ~n16197 ;
  assign n16439 = n33271 & n16438 ;
  assign n13184 = n4686 & n13182 ;
  assign n10728 = n4706 & n10727 ;
  assign n10753 = n4726 & n31999 ;
  assign n16440 = n10728 | n10753 ;
  assign n16441 = n4748 & n13151 ;
  assign n16442 = n16440 | n16441 ;
  assign n16443 = n13184 | n16442 ;
  assign n16444 = x20 | n16443 ;
  assign n16445 = x20 & n16443 ;
  assign n33272 = ~n16445 ;
  assign n16446 = n16444 & n33272 ;
  assign n16448 = n16439 | n16446 ;
  assign n33273 = ~n16439 ;
  assign n16447 = n33273 & n16446 ;
  assign n33274 = ~n16446 ;
  assign n16449 = n16439 & n33274 ;
  assign n16450 = n16447 | n16449 ;
  assign n11691 = n4686 & n32125 ;
  assign n10766 = n4706 & n31999 ;
  assign n10784 = n4726 & n10773 ;
  assign n16451 = n10766 | n10784 ;
  assign n16452 = n4748 & n10727 ;
  assign n16453 = n16451 | n16452 ;
  assign n16454 = n11691 | n16453 ;
  assign n16455 = x20 | n16454 ;
  assign n16456 = x20 & n16454 ;
  assign n33275 = ~n16456 ;
  assign n16457 = n16455 & n33275 ;
  assign n16191 = n16117 & n16190 ;
  assign n16458 = n16117 | n16190 ;
  assign n33276 = ~n16191 ;
  assign n16459 = n33276 & n16458 ;
  assign n13235 = n4686 & n32477 ;
  assign n10783 = n4706 & n10773 ;
  assign n10801 = n4726 & n31998 ;
  assign n16460 = n10783 | n10801 ;
  assign n16461 = n4748 & n32478 ;
  assign n16462 = n16460 | n16461 ;
  assign n16463 = n13235 | n16462 ;
  assign n16464 = x20 | n16463 ;
  assign n16465 = x20 & n16463 ;
  assign n33277 = ~n16465 ;
  assign n16466 = n16464 & n33277 ;
  assign n16468 = n16459 | n16466 ;
  assign n33278 = ~n16459 ;
  assign n16467 = n33278 & n16466 ;
  assign n33279 = ~n16466 ;
  assign n16469 = n16459 & n33279 ;
  assign n16470 = n16467 | n16469 ;
  assign n16188 = n16132 & n16187 ;
  assign n16471 = n16132 | n16187 ;
  assign n33280 = ~n16188 ;
  assign n16472 = n33280 & n16471 ;
  assign n13286 = n4686 & n32482 ;
  assign n10799 = n4706 & n31998 ;
  assign n10820 = n4726 & n10818 ;
  assign n16473 = n10799 | n10820 ;
  assign n16474 = n4748 & n13292 ;
  assign n16475 = n16473 | n16474 ;
  assign n16476 = n13286 | n16475 ;
  assign n16477 = x20 | n16476 ;
  assign n16478 = x20 & n16476 ;
  assign n33281 = ~n16478 ;
  assign n16479 = n16477 & n33281 ;
  assign n16481 = n16472 | n16479 ;
  assign n16480 = n16472 & n16479 ;
  assign n33282 = ~n16480 ;
  assign n16482 = n33282 & n16481 ;
  assign n16185 = n16144 & n16184 ;
  assign n16483 = n16144 | n16184 ;
  assign n33283 = ~n16185 ;
  assign n16484 = n33283 & n16483 ;
  assign n13323 = n4686 & n32488 ;
  assign n10819 = n4706 & n10818 ;
  assign n10844 = n4726 & n10841 ;
  assign n16485 = n10819 | n10844 ;
  assign n16486 = n4748 & n31998 ;
  assign n16487 = n16485 | n16486 ;
  assign n16488 = n13323 | n16487 ;
  assign n16489 = x20 | n16488 ;
  assign n16490 = x20 & n16488 ;
  assign n33284 = ~n16490 ;
  assign n16491 = n16489 & n33284 ;
  assign n16493 = n16484 | n16491 ;
  assign n33285 = ~n16484 ;
  assign n16492 = n33285 & n16491 ;
  assign n33286 = ~n16491 ;
  assign n16494 = n16484 & n33286 ;
  assign n16495 = n16492 | n16494 ;
  assign n13390 = n4686 & n13382 ;
  assign n10856 = n4706 & n10841 ;
  assign n10866 = n4726 & n10865 ;
  assign n16496 = n10856 | n10866 ;
  assign n16497 = n4748 & n10818 ;
  assign n16498 = n16496 | n16497 ;
  assign n16499 = n13390 | n16498 ;
  assign n33287 = ~n16499 ;
  assign n16500 = x20 & n33287 ;
  assign n16501 = n30374 & n16499 ;
  assign n16502 = n16500 | n16501 ;
  assign n33288 = ~n16182 ;
  assign n16503 = n16181 & n33288 ;
  assign n16504 = n16183 | n16503 ;
  assign n16506 = n16502 & n16504 ;
  assign n33289 = ~n15784 ;
  assign n16161 = n33289 & n16160 ;
  assign n33290 = ~n16160 ;
  assign n16507 = n15784 & n33290 ;
  assign n16508 = n16161 | n16507 ;
  assign n33291 = ~n16169 ;
  assign n16509 = n33291 & n16508 ;
  assign n33292 = ~n16508 ;
  assign n16510 = n16169 & n33292 ;
  assign n16511 = n16509 | n16510 ;
  assign n13463 = n4686 & n13456 ;
  assign n10877 = n4706 & n10865 ;
  assign n10902 = n4726 & n10892 ;
  assign n16512 = n10877 | n10902 ;
  assign n16513 = n4748 & n10841 ;
  assign n16514 = n16512 | n16513 ;
  assign n16515 = n13463 | n16514 ;
  assign n16516 = x20 | n16515 ;
  assign n16517 = x20 & n16515 ;
  assign n33293 = ~n16517 ;
  assign n16518 = n16516 & n33293 ;
  assign n16519 = n16511 & n16518 ;
  assign n16520 = n16511 | n16518 ;
  assign n33294 = ~n16519 ;
  assign n16521 = n33294 & n16520 ;
  assign n16158 = n16151 & n16157 ;
  assign n33295 = ~n16158 ;
  assign n16522 = n33295 & n16159 ;
  assign n13533 = n4686 & n32502 ;
  assign n10895 = n4706 & n10892 ;
  assign n10919 = n4726 & n32503 ;
  assign n16523 = n10895 | n10919 ;
  assign n16524 = n4748 & n10865 ;
  assign n16525 = n16523 | n16524 ;
  assign n16526 = n13533 | n16525 ;
  assign n16527 = x20 | n16526 ;
  assign n16528 = x20 & n16526 ;
  assign n33296 = ~n16528 ;
  assign n16529 = n16527 & n33296 ;
  assign n16531 = n16522 | n16529 ;
  assign n16530 = n16522 & n16529 ;
  assign n33297 = ~n16530 ;
  assign n16532 = n33297 & n16531 ;
  assign n16533 = n4683 & n32507 ;
  assign n14865 = n4686 & n14859 ;
  assign n16534 = n4748 & n31995 ;
  assign n16535 = n4706 & n32507 ;
  assign n16536 = n16534 | n16535 ;
  assign n16537 = n14865 | n16536 ;
  assign n16538 = n16533 | n16537 ;
  assign n16539 = x20 & n16538 ;
  assign n10956 = n4748 & n10940 ;
  assign n16540 = n4706 & n31995 ;
  assign n16541 = n4726 & n32507 ;
  assign n16542 = n16540 | n16541 ;
  assign n16543 = n10956 | n16542 ;
  assign n16544 = n4686 & n13637 ;
  assign n16545 = n16543 | n16544 ;
  assign n16547 = n16539 | n16545 ;
  assign n33298 = ~n16547 ;
  assign n16548 = x20 & n33298 ;
  assign n16550 = n16145 | n16548 ;
  assign n13698 = n4686 & n13690 ;
  assign n10953 = n4706 & n10940 ;
  assign n10982 = n4726 & n31995 ;
  assign n16551 = n10953 | n10982 ;
  assign n16552 = n4748 & n32503 ;
  assign n16553 = n16551 | n16552 ;
  assign n16554 = n13698 | n16553 ;
  assign n33299 = ~n16554 ;
  assign n16555 = x20 & n33299 ;
  assign n16556 = n30374 & n16554 ;
  assign n16557 = n16555 | n16556 ;
  assign n16558 = n16550 & n16557 ;
  assign n16559 = x23 & n16145 ;
  assign n33300 = ~n16149 ;
  assign n16560 = n33300 & n16559 ;
  assign n33301 = ~n16559 ;
  assign n16561 = n16149 & n33301 ;
  assign n16562 = n16560 | n16561 ;
  assign n16564 = n16558 | n16562 ;
  assign n13764 = n4686 & n13756 ;
  assign n10918 = n4706 & n32503 ;
  assign n10957 = n4726 & n10940 ;
  assign n16565 = n10918 | n10957 ;
  assign n16566 = n4748 & n10892 ;
  assign n16567 = n16565 | n16566 ;
  assign n16568 = n13764 | n16567 ;
  assign n16569 = x20 | n16568 ;
  assign n16570 = x20 & n16568 ;
  assign n33302 = ~n16570 ;
  assign n16571 = n16569 & n33302 ;
  assign n16563 = n16558 & n16562 ;
  assign n33303 = ~n16563 ;
  assign n16572 = n33303 & n16564 ;
  assign n33304 = ~n16571 ;
  assign n16573 = n33304 & n16572 ;
  assign n33305 = ~n16573 ;
  assign n16575 = n16564 & n33305 ;
  assign n33306 = ~n16575 ;
  assign n16577 = n16532 & n33306 ;
  assign n33307 = ~n16577 ;
  assign n16578 = n16531 & n33307 ;
  assign n16579 = n16521 & n16578 ;
  assign n16580 = n16519 | n16579 ;
  assign n16505 = n16502 | n16504 ;
  assign n33308 = ~n16506 ;
  assign n16581 = n16505 & n33308 ;
  assign n16582 = n16580 & n16581 ;
  assign n16583 = n16506 | n16582 ;
  assign n33309 = ~n16583 ;
  assign n16584 = n16495 & n33309 ;
  assign n33310 = ~n16584 ;
  assign n16585 = n16493 & n33310 ;
  assign n33311 = ~n16585 ;
  assign n16587 = n16482 & n33311 ;
  assign n33312 = ~n16587 ;
  assign n16588 = n16481 & n33312 ;
  assign n33313 = ~n16588 ;
  assign n16590 = n16470 & n33313 ;
  assign n33314 = ~n16590 ;
  assign n16591 = n16468 & n33314 ;
  assign n16593 = n16457 | n16591 ;
  assign n16194 = n16104 & n16193 ;
  assign n16594 = n16104 | n16193 ;
  assign n33315 = ~n16194 ;
  assign n16595 = n33315 & n16594 ;
  assign n16592 = n16457 & n16591 ;
  assign n33316 = ~n16592 ;
  assign n16596 = n33316 & n16593 ;
  assign n33317 = ~n16595 ;
  assign n16597 = n33317 & n16596 ;
  assign n33318 = ~n16597 ;
  assign n16598 = n16593 & n33318 ;
  assign n33319 = ~n16598 ;
  assign n16600 = n16450 & n33319 ;
  assign n33320 = ~n16600 ;
  assign n16601 = n16448 & n33320 ;
  assign n16603 = n16437 | n16601 ;
  assign n33321 = ~n16435 ;
  assign n16604 = n33321 & n16603 ;
  assign n16606 = n16424 | n16604 ;
  assign n33322 = ~n16422 ;
  assign n16607 = n33322 & n16606 ;
  assign n33323 = ~n16607 ;
  assign n16609 = n16411 & n33323 ;
  assign n33324 = ~n16609 ;
  assign n16610 = n16409 & n33324 ;
  assign n16612 = n16398 | n16610 ;
  assign n33325 = ~n16396 ;
  assign n16613 = n33325 & n16612 ;
  assign n16615 = n16385 | n16613 ;
  assign n33326 = ~n16384 ;
  assign n16616 = n33326 & n16615 ;
  assign n33327 = ~n16616 ;
  assign n16618 = n16373 & n33327 ;
  assign n33328 = ~n16618 ;
  assign n16619 = n16371 & n33328 ;
  assign n33329 = ~n16351 ;
  assign n16359 = n33329 & n16358 ;
  assign n33330 = ~n16358 ;
  assign n16620 = n16351 & n33330 ;
  assign n16621 = n16359 | n16620 ;
  assign n16622 = n16619 & n16621 ;
  assign n16623 = n16360 | n16622 ;
  assign n33331 = ~n16623 ;
  assign n16624 = n16349 & n33331 ;
  assign n33332 = ~n16624 ;
  assign n16625 = n16347 & n33332 ;
  assign n33333 = ~n16625 ;
  assign n16627 = n16336 & n33333 ;
  assign n33334 = ~n16627 ;
  assign n16628 = n16334 & n33334 ;
  assign n33335 = ~n16628 ;
  assign n16630 = n16323 & n33335 ;
  assign n33336 = ~n16630 ;
  assign n16631 = n16321 & n33336 ;
  assign n33337 = ~n16301 ;
  assign n16309 = n33337 & n16308 ;
  assign n16632 = n16309 | n16310 ;
  assign n16634 = n16631 | n16632 ;
  assign n33338 = ~n16310 ;
  assign n16635 = n33338 & n16634 ;
  assign n33339 = ~n16635 ;
  assign n16637 = n16299 & n33339 ;
  assign n33340 = ~n16637 ;
  assign n16638 = n16298 & n33340 ;
  assign n16640 = n16287 | n16638 ;
  assign n33341 = ~n16286 ;
  assign n16641 = n33341 & n16640 ;
  assign n16643 = n16275 | n16641 ;
  assign n33342 = ~n16273 ;
  assign n16644 = n33342 & n16643 ;
  assign n15235 = x8 & n32883 ;
  assign n16645 = n70 | n15235 ;
  assign n16646 = x7 & n15221 ;
  assign n16647 = n16645 | n16646 ;
  assign n16648 = n30018 & n16647 ;
  assign n16650 = n16644 | n16648 ;
  assign n16247 = n16243 & n16245 ;
  assign n16651 = n16243 | n16245 ;
  assign n33343 = ~n16247 ;
  assign n16652 = n33343 & n16651 ;
  assign n16649 = n16644 & n16648 ;
  assign n33344 = ~n16649 ;
  assign n16653 = n33344 & n16650 ;
  assign n33345 = ~n16652 ;
  assign n16654 = n33345 & n16653 ;
  assign n33346 = ~n16654 ;
  assign n16655 = n16650 & n33346 ;
  assign n33347 = ~n16655 ;
  assign n16657 = n16262 & n33347 ;
  assign n33348 = ~n16262 ;
  assign n16656 = n33348 & n16655 ;
  assign n16658 = n16656 | n16657 ;
  assign n33349 = ~n16653 ;
  assign n16659 = n16652 & n33349 ;
  assign n16660 = n16654 | n16659 ;
  assign n33350 = ~n16275 ;
  assign n16642 = n33350 & n16641 ;
  assign n33351 = ~n16641 ;
  assign n16661 = n16275 & n33351 ;
  assign n16662 = n16642 | n16661 ;
  assign n15519 = n67 & n15516 ;
  assign n15222 = n69 & n15221 ;
  assign n16663 = n7017 | n15222 ;
  assign n16664 = n7041 & n32890 ;
  assign n16665 = n16663 | n16664 ;
  assign n16666 = n15519 | n16665 ;
  assign n16667 = x8 | n16666 ;
  assign n16668 = x8 & n16666 ;
  assign n33352 = ~n16668 ;
  assign n16669 = n16667 & n33352 ;
  assign n33353 = ~n16669 ;
  assign n16671 = n16662 & n33353 ;
  assign n16670 = n16662 & n16669 ;
  assign n16672 = n16662 | n16669 ;
  assign n33354 = ~n16670 ;
  assign n16673 = n33354 & n16672 ;
  assign n33355 = ~n16287 ;
  assign n16639 = n33355 & n16638 ;
  assign n33356 = ~n16638 ;
  assign n16674 = n16287 & n33356 ;
  assign n16675 = n16639 | n16674 ;
  assign n15530 = n7068 & n15526 ;
  assign n15170 = n7041 & n32876 ;
  assign n15226 = n7017 & n15221 ;
  assign n16676 = n15170 | n15226 ;
  assign n16677 = n69 & n32890 ;
  assign n16678 = n16676 | n16677 ;
  assign n16679 = n15530 | n16678 ;
  assign n16680 = x8 | n16679 ;
  assign n16681 = x8 & n16679 ;
  assign n33357 = ~n16681 ;
  assign n16682 = n16680 & n33357 ;
  assign n33358 = ~n16682 ;
  assign n16684 = n16675 & n33358 ;
  assign n16683 = n16675 & n16682 ;
  assign n16685 = n16675 | n16682 ;
  assign n33359 = ~n16683 ;
  assign n16686 = n33359 & n16685 ;
  assign n16636 = n16299 & n16635 ;
  assign n16687 = n16299 | n16635 ;
  assign n33360 = ~n16636 ;
  assign n16688 = n33360 & n16687 ;
  assign n15290 = n6272 & n15288 ;
  assign n14494 = n6190 & n32707 ;
  assign n14520 = n6244 & n32706 ;
  assign n16689 = n14494 | n14520 ;
  assign n16690 = n6217 & n15081 ;
  assign n16691 = n16689 | n16690 ;
  assign n16692 = n15290 | n16691 ;
  assign n16693 = x11 | n16692 ;
  assign n16694 = x11 & n16692 ;
  assign n33361 = ~n16694 ;
  assign n16695 = n16693 & n33361 ;
  assign n16697 = n16688 & n16695 ;
  assign n33362 = ~n16688 ;
  assign n16696 = n33362 & n16695 ;
  assign n33363 = ~n16695 ;
  assign n16698 = n16688 & n33363 ;
  assign n16699 = n16696 | n16698 ;
  assign n33364 = ~n16632 ;
  assign n16633 = n16631 & n33364 ;
  assign n33365 = ~n16631 ;
  assign n16700 = n33365 & n16632 ;
  assign n16701 = n16633 | n16700 ;
  assign n14188 = n5937 & n14183 ;
  assign n14129 = n5970 & n14124 ;
  assign n14152 = n5994 & n14147 ;
  assign n16702 = n14129 | n14152 ;
  assign n16703 = n6018 & n14196 ;
  assign n16704 = n16702 | n16703 ;
  assign n16705 = n14188 | n16704 ;
  assign n16706 = x14 | n16705 ;
  assign n16707 = x14 & n16705 ;
  assign n33366 = ~n16707 ;
  assign n16708 = n16706 & n33366 ;
  assign n33367 = ~n16708 ;
  assign n16710 = n16701 & n33367 ;
  assign n16629 = n16323 & n16628 ;
  assign n16711 = n16323 | n16628 ;
  assign n33368 = ~n16629 ;
  assign n16712 = n33368 & n16711 ;
  assign n13852 = n37300 & n32557 ;
  assign n12549 = n5166 & n32354 ;
  assign n13084 = n5144 & n13077 ;
  assign n16713 = n12549 | n13084 ;
  assign n16714 = n5191 & n32456 ;
  assign n16715 = n16713 | n16714 ;
  assign n16716 = n13852 | n16715 ;
  assign n16717 = x17 | n16716 ;
  assign n16718 = x17 & n16716 ;
  assign n33369 = ~n16718 ;
  assign n16719 = n16717 & n33369 ;
  assign n16721 = n16712 | n16719 ;
  assign n33370 = ~n16712 ;
  assign n16720 = n33370 & n16719 ;
  assign n33371 = ~n16719 ;
  assign n16722 = n16712 & n33371 ;
  assign n16723 = n16720 | n16722 ;
  assign n16626 = n16336 & n16625 ;
  assign n16724 = n16336 | n16625 ;
  assign n33372 = ~n16626 ;
  assign n16725 = n33372 & n16724 ;
  assign n14260 = n37300 & n32641 ;
  assign n12552 = n5144 & n32354 ;
  assign n12571 = n5166 & n12570 ;
  assign n16726 = n12552 | n12571 ;
  assign n16727 = n5191 & n13077 ;
  assign n16728 = n16726 | n16727 ;
  assign n16729 = n14260 | n16728 ;
  assign n16730 = x17 | n16729 ;
  assign n16731 = x17 & n16729 ;
  assign n33373 = ~n16731 ;
  assign n16732 = n16730 & n33373 ;
  assign n16734 = n16725 | n16732 ;
  assign n33374 = ~n16725 ;
  assign n16733 = n33374 & n16732 ;
  assign n33375 = ~n16732 ;
  assign n16735 = n16725 & n33375 ;
  assign n16736 = n16733 | n16735 ;
  assign n33376 = ~n16349 ;
  assign n16737 = n33376 & n16623 ;
  assign n16738 = n16624 | n16737 ;
  assign n12635 = n37300 & n32356 ;
  assign n12585 = n5144 & n12570 ;
  assign n12599 = n5166 & n12595 ;
  assign n16739 = n12585 | n12599 ;
  assign n16740 = n5191 & n32354 ;
  assign n16741 = n16739 | n16740 ;
  assign n16742 = n12635 | n16741 ;
  assign n16743 = x17 | n16742 ;
  assign n16744 = x17 & n16742 ;
  assign n33377 = ~n16744 ;
  assign n16745 = n16743 & n33377 ;
  assign n16747 = n16738 | n16745 ;
  assign n33378 = ~n16738 ;
  assign n16746 = n33378 & n16745 ;
  assign n33379 = ~n16745 ;
  assign n16748 = n16738 & n33379 ;
  assign n16749 = n16746 | n16748 ;
  assign n16750 = n16619 | n16621 ;
  assign n33380 = ~n16622 ;
  assign n16751 = n33380 & n16750 ;
  assign n12687 = n37300 & n12681 ;
  assign n12139 = n5166 & n32253 ;
  assign n12605 = n5144 & n12595 ;
  assign n16752 = n12139 | n12605 ;
  assign n16753 = n5191 & n12570 ;
  assign n16754 = n16752 | n16753 ;
  assign n16755 = n12687 | n16754 ;
  assign n16756 = x17 | n16755 ;
  assign n16757 = x17 & n16755 ;
  assign n33381 = ~n16757 ;
  assign n16758 = n16756 & n33381 ;
  assign n16759 = n16751 & n16758 ;
  assign n16617 = n16373 & n16616 ;
  assign n16760 = n16373 | n16616 ;
  assign n33382 = ~n16617 ;
  assign n16761 = n33382 & n16760 ;
  assign n13828 = n37300 & n32550 ;
  assign n12137 = n5144 & n32253 ;
  assign n12168 = n5166 & n12161 ;
  assign n16762 = n12137 | n12168 ;
  assign n16763 = n5191 & n12595 ;
  assign n16764 = n16762 | n16763 ;
  assign n16765 = n13828 | n16764 ;
  assign n16766 = x17 | n16765 ;
  assign n16767 = x17 & n16765 ;
  assign n33383 = ~n16767 ;
  assign n16768 = n16766 & n33383 ;
  assign n16770 = n16761 | n16768 ;
  assign n33384 = ~n16761 ;
  assign n16769 = n33384 & n16768 ;
  assign n33385 = ~n16768 ;
  assign n16771 = n16761 & n33385 ;
  assign n16772 = n16769 | n16771 ;
  assign n33386 = ~n16385 ;
  assign n16614 = n33386 & n16613 ;
  assign n33387 = ~n16613 ;
  assign n16773 = n16385 & n33387 ;
  assign n16774 = n16614 | n16773 ;
  assign n12198 = n37300 & n32255 ;
  assign n11850 = n5166 & n32176 ;
  assign n12162 = n5144 & n12161 ;
  assign n16775 = n11850 | n12162 ;
  assign n16776 = n5191 & n32253 ;
  assign n16777 = n16775 | n16776 ;
  assign n16778 = n12198 | n16777 ;
  assign n16779 = x17 | n16778 ;
  assign n16780 = x17 & n16778 ;
  assign n33388 = ~n16780 ;
  assign n16781 = n16779 & n33388 ;
  assign n33389 = ~n16781 ;
  assign n16783 = n16774 & n33389 ;
  assign n33390 = ~n16398 ;
  assign n16611 = n33390 & n16610 ;
  assign n33391 = ~n16610 ;
  assign n16784 = n16398 & n33391 ;
  assign n16785 = n16611 | n16784 ;
  assign n12661 = n37300 & n32362 ;
  assign n11440 = n5166 & n11430 ;
  assign n11855 = n5144 & n32176 ;
  assign n16786 = n11440 | n11855 ;
  assign n16787 = n5191 & n12161 ;
  assign n16788 = n16786 | n16787 ;
  assign n16789 = n12661 | n16788 ;
  assign n16790 = x17 | n16789 ;
  assign n16791 = x17 & n16789 ;
  assign n33392 = ~n16791 ;
  assign n16792 = n16790 & n33392 ;
  assign n33393 = ~n16792 ;
  assign n16794 = n16785 & n33393 ;
  assign n16793 = n16785 & n16792 ;
  assign n16795 = n16785 | n16792 ;
  assign n33394 = ~n16793 ;
  assign n16796 = n33394 & n16795 ;
  assign n16608 = n16411 & n16607 ;
  assign n16797 = n16411 | n16607 ;
  assign n33395 = ~n16608 ;
  assign n16798 = n33395 & n16797 ;
  assign n11877 = n37300 & n32178 ;
  assign n11435 = n5144 & n11430 ;
  assign n11478 = n5166 & n11476 ;
  assign n16799 = n11435 | n11478 ;
  assign n16800 = n5191 & n32176 ;
  assign n16801 = n16799 | n16800 ;
  assign n16802 = n11877 | n16801 ;
  assign n16803 = x17 | n16802 ;
  assign n16804 = x17 & n16802 ;
  assign n33396 = ~n16804 ;
  assign n16805 = n16803 & n33396 ;
  assign n16807 = n16798 & n16805 ;
  assign n33397 = ~n16798 ;
  assign n16806 = n33397 & n16805 ;
  assign n33398 = ~n16805 ;
  assign n16808 = n16798 & n33398 ;
  assign n16809 = n16806 | n16808 ;
  assign n11472 = n37300 & n11463 ;
  assign n10672 = n5166 & n10656 ;
  assign n11490 = n5144 & n11476 ;
  assign n16810 = n10672 | n11490 ;
  assign n16811 = n5191 & n11430 ;
  assign n16812 = n16810 | n16811 ;
  assign n16813 = n11472 | n16812 ;
  assign n16814 = x17 | n16813 ;
  assign n16815 = x17 & n16813 ;
  assign n33399 = ~n16815 ;
  assign n16816 = n16814 & n33399 ;
  assign n33400 = ~n16424 ;
  assign n16605 = n33400 & n16604 ;
  assign n33401 = ~n16604 ;
  assign n16817 = n16424 & n33401 ;
  assign n16818 = n16605 | n16817 ;
  assign n33402 = ~n16816 ;
  assign n16819 = n33402 & n16818 ;
  assign n33403 = ~n16818 ;
  assign n16820 = n16816 & n33403 ;
  assign n16821 = n16819 | n16820 ;
  assign n33404 = ~n16437 ;
  assign n16602 = n33404 & n16601 ;
  assign n33405 = ~n16601 ;
  assign n16822 = n16437 & n33405 ;
  assign n16823 = n16602 | n16822 ;
  assign n11520 = n37300 & n11511 ;
  assign n10670 = n5144 & n10656 ;
  assign n11041 = n5166 & n10679 ;
  assign n16824 = n10670 | n11041 ;
  assign n16825 = n5191 & n11452 ;
  assign n16826 = n16824 | n16825 ;
  assign n16827 = n11520 | n16826 ;
  assign n16828 = x17 | n16827 ;
  assign n16829 = x17 & n16827 ;
  assign n33406 = ~n16829 ;
  assign n16830 = n16828 & n33406 ;
  assign n33407 = ~n16830 ;
  assign n16832 = n16823 & n33407 ;
  assign n16831 = n16823 & n16830 ;
  assign n16833 = n16823 | n16830 ;
  assign n33408 = ~n16831 ;
  assign n16834 = n33408 & n16833 ;
  assign n16599 = n16450 & n16598 ;
  assign n16835 = n16450 | n16598 ;
  assign n33409 = ~n16599 ;
  assign n16836 = n33409 & n16835 ;
  assign n11038 = n37300 & n11030 ;
  assign n10695 = n5166 & n10681 ;
  assign n11056 = n5144 & n10679 ;
  assign n16837 = n10695 | n11056 ;
  assign n16838 = n5191 & n10656 ;
  assign n16839 = n16837 | n16838 ;
  assign n16840 = n11038 | n16839 ;
  assign n16841 = x17 | n16840 ;
  assign n16842 = x17 & n16840 ;
  assign n33410 = ~n16842 ;
  assign n16843 = n16841 & n33410 ;
  assign n16845 = n16836 | n16843 ;
  assign n33411 = ~n16836 ;
  assign n16844 = n33411 & n16843 ;
  assign n33412 = ~n16843 ;
  assign n16846 = n16836 & n33412 ;
  assign n16847 = n16844 | n16846 ;
  assign n33413 = ~n16596 ;
  assign n16848 = n16595 & n33413 ;
  assign n16849 = n16597 | n16848 ;
  assign n11542 = n37300 & n11536 ;
  assign n10696 = n5144 & n10681 ;
  assign n10704 = n5166 & n10703 ;
  assign n16850 = n10696 | n10704 ;
  assign n16851 = n5191 & n10679 ;
  assign n16852 = n16850 | n16851 ;
  assign n16853 = n11542 | n16852 ;
  assign n16854 = x17 | n16853 ;
  assign n16855 = x17 & n16853 ;
  assign n33414 = ~n16855 ;
  assign n16856 = n16854 & n33414 ;
  assign n16858 = n16849 | n16856 ;
  assign n33415 = ~n16849 ;
  assign n16857 = n33415 & n16856 ;
  assign n33416 = ~n16856 ;
  assign n16859 = n16849 & n33416 ;
  assign n16860 = n16857 | n16859 ;
  assign n16589 = n16470 & n16588 ;
  assign n16861 = n16470 | n16588 ;
  assign n33417 = ~n16589 ;
  assign n16862 = n33417 & n16861 ;
  assign n13163 = n37300 & n13157 ;
  assign n10723 = n5144 & n10703 ;
  assign n10739 = n5166 & n10727 ;
  assign n16863 = n10723 | n10739 ;
  assign n16864 = n5191 & n10681 ;
  assign n16865 = n16863 | n16864 ;
  assign n16866 = n13163 | n16865 ;
  assign n16867 = x17 | n16866 ;
  assign n16868 = x17 & n16866 ;
  assign n33418 = ~n16868 ;
  assign n16869 = n16867 & n33418 ;
  assign n16871 = n16862 | n16869 ;
  assign n33419 = ~n16862 ;
  assign n16870 = n33419 & n16869 ;
  assign n33420 = ~n16869 ;
  assign n16872 = n16862 & n33420 ;
  assign n16873 = n16870 | n16872 ;
  assign n16586 = n16482 & n16585 ;
  assign n16874 = n16482 | n16585 ;
  assign n33421 = ~n16586 ;
  assign n16875 = n33421 & n16874 ;
  assign n13186 = n37300 & n13182 ;
  assign n10741 = n5144 & n10727 ;
  assign n10751 = n5166 & n31999 ;
  assign n16876 = n10741 | n10751 ;
  assign n16877 = n5191 & n13151 ;
  assign n16878 = n16876 | n16877 ;
  assign n16879 = n13186 | n16878 ;
  assign n16880 = x17 | n16879 ;
  assign n16881 = x17 & n16879 ;
  assign n33422 = ~n16881 ;
  assign n16882 = n16880 & n33422 ;
  assign n16884 = n16875 | n16882 ;
  assign n16883 = n16875 & n16882 ;
  assign n33423 = ~n16883 ;
  assign n16885 = n33423 & n16884 ;
  assign n33424 = ~n16495 ;
  assign n16886 = n33424 & n16583 ;
  assign n16887 = n16584 | n16886 ;
  assign n11692 = n37300 & n32125 ;
  assign n10752 = n5144 & n31999 ;
  assign n10787 = n5166 & n10773 ;
  assign n16888 = n10752 | n10787 ;
  assign n16889 = n5191 & n10727 ;
  assign n16890 = n16888 | n16889 ;
  assign n16891 = n11692 | n16890 ;
  assign n16892 = x17 | n16891 ;
  assign n16893 = x17 & n16891 ;
  assign n33425 = ~n16893 ;
  assign n16894 = n16892 & n33425 ;
  assign n16896 = n16887 | n16894 ;
  assign n16895 = n16887 & n16894 ;
  assign n33426 = ~n16895 ;
  assign n16897 = n33426 & n16896 ;
  assign n13236 = n37300 & n32477 ;
  assign n10788 = n5144 & n10773 ;
  assign n10796 = n5166 & n31998 ;
  assign n16898 = n10788 | n10796 ;
  assign n16899 = n5191 & n32478 ;
  assign n16900 = n16898 | n16899 ;
  assign n16901 = n13236 | n16900 ;
  assign n16902 = x17 | n16901 ;
  assign n16903 = x17 & n16901 ;
  assign n33427 = ~n16903 ;
  assign n16904 = n16902 & n33427 ;
  assign n16905 = n16580 | n16581 ;
  assign n33428 = ~n16582 ;
  assign n16906 = n33428 & n16905 ;
  assign n16908 = n16904 | n16906 ;
  assign n16907 = n16904 & n16906 ;
  assign n33429 = ~n16907 ;
  assign n16909 = n33429 & n16908 ;
  assign n16910 = n16521 | n16578 ;
  assign n33430 = ~n16579 ;
  assign n16911 = n33430 & n16910 ;
  assign n13287 = n37300 & n32482 ;
  assign n10809 = n5144 & n31998 ;
  assign n10831 = n5166 & n10818 ;
  assign n16912 = n10809 | n10831 ;
  assign n16913 = n5191 & n13292 ;
  assign n16914 = n16912 | n16913 ;
  assign n16915 = n13287 | n16914 ;
  assign n16916 = x17 | n16915 ;
  assign n16917 = x17 & n16915 ;
  assign n33431 = ~n16917 ;
  assign n16918 = n16916 & n33431 ;
  assign n16920 = n16911 | n16918 ;
  assign n13324 = n37300 & n32488 ;
  assign n10832 = n5144 & n10818 ;
  assign n10842 = n5166 & n10841 ;
  assign n16921 = n10832 | n10842 ;
  assign n16922 = n5191 & n31998 ;
  assign n16923 = n16921 | n16922 ;
  assign n16924 = n13324 | n16923 ;
  assign n16925 = x17 | n16924 ;
  assign n16926 = x17 & n16924 ;
  assign n33432 = ~n16926 ;
  assign n16927 = n16925 & n33432 ;
  assign n13391 = n37300 & n13382 ;
  assign n10858 = n5144 & n10841 ;
  assign n10878 = n5166 & n10865 ;
  assign n16928 = n10858 | n10878 ;
  assign n16929 = n5191 & n10818 ;
  assign n16930 = n16928 | n16929 ;
  assign n16931 = n13391 | n16930 ;
  assign n33433 = ~n16931 ;
  assign n16932 = x17 & n33433 ;
  assign n16933 = n30580 & n16931 ;
  assign n16934 = n16932 | n16933 ;
  assign n16574 = n16571 & n16572 ;
  assign n16935 = n16571 | n16572 ;
  assign n33434 = ~n16574 ;
  assign n16936 = n33434 & n16935 ;
  assign n16937 = n16934 | n16936 ;
  assign n33435 = ~n16145 ;
  assign n16549 = n33435 & n16548 ;
  assign n33436 = ~n16548 ;
  assign n16938 = n16145 & n33436 ;
  assign n16939 = n16549 | n16938 ;
  assign n33437 = ~n16557 ;
  assign n16940 = n33437 & n16939 ;
  assign n33438 = ~n16939 ;
  assign n16941 = n16557 & n33438 ;
  assign n16942 = n16940 | n16941 ;
  assign n13459 = n37300 & n13456 ;
  assign n10880 = n5144 & n10865 ;
  assign n10893 = n5166 & n10892 ;
  assign n16943 = n10880 | n10893 ;
  assign n16944 = n5191 & n10841 ;
  assign n16945 = n16943 | n16944 ;
  assign n16946 = n13459 | n16945 ;
  assign n16947 = x17 | n16946 ;
  assign n16948 = x17 & n16946 ;
  assign n33439 = ~n16948 ;
  assign n16949 = n16947 & n33439 ;
  assign n16950 = n16942 & n16949 ;
  assign n16951 = n16942 | n16949 ;
  assign n33440 = ~n16950 ;
  assign n16952 = n33440 & n16951 ;
  assign n16546 = n16539 & n16545 ;
  assign n33441 = ~n16546 ;
  assign n16953 = n33441 & n16547 ;
  assign n13534 = n37300 & n32502 ;
  assign n10909 = n5144 & n10892 ;
  assign n10933 = n5166 & n32503 ;
  assign n16954 = n10909 | n10933 ;
  assign n16955 = n5191 & n10865 ;
  assign n16956 = n16954 | n16955 ;
  assign n16957 = n13534 | n16956 ;
  assign n16958 = x17 | n16957 ;
  assign n16959 = x17 & n16957 ;
  assign n33442 = ~n16959 ;
  assign n16960 = n16958 & n33442 ;
  assign n16961 = n16953 & n16960 ;
  assign n16962 = x20 & n16533 ;
  assign n33443 = ~n16537 ;
  assign n16963 = n33443 & n16962 ;
  assign n33444 = ~n16962 ;
  assign n16964 = n16537 & n33444 ;
  assign n16965 = n16963 | n16964 ;
  assign n13758 = n37300 & n13756 ;
  assign n10927 = n5144 & n32503 ;
  assign n10951 = n5166 & n10940 ;
  assign n16966 = n10927 | n10951 ;
  assign n16967 = n5191 & n10892 ;
  assign n16968 = n16966 | n16967 ;
  assign n16969 = n13758 | n16968 ;
  assign n16970 = x17 | n16969 ;
  assign n16971 = x17 & n16969 ;
  assign n33445 = ~n16971 ;
  assign n16972 = n16970 & n33445 ;
  assign n16974 = n16965 | n16972 ;
  assign n16975 = n37297 & n32507 ;
  assign n14861 = n37300 & n14859 ;
  assign n16976 = n5191 & n31995 ;
  assign n16977 = n5144 & n32507 ;
  assign n16978 = n16976 | n16977 ;
  assign n16979 = n14861 | n16978 ;
  assign n16980 = n16975 | n16979 ;
  assign n16981 = x17 & n16980 ;
  assign n10948 = n5191 & n10940 ;
  assign n16982 = n5144 & n31995 ;
  assign n16983 = n5166 & n32507 ;
  assign n16984 = n16982 | n16983 ;
  assign n16985 = n10948 | n16984 ;
  assign n16986 = n37300 & n13637 ;
  assign n16987 = n16985 | n16986 ;
  assign n16989 = n16981 | n16987 ;
  assign n33446 = ~n16989 ;
  assign n16990 = x17 & n33446 ;
  assign n16992 = n16533 | n16990 ;
  assign n13696 = n37300 & n13690 ;
  assign n10947 = n5144 & n10940 ;
  assign n10980 = n5166 & n31995 ;
  assign n16993 = n10947 | n10980 ;
  assign n16994 = n5191 & n32503 ;
  assign n16995 = n16993 | n16994 ;
  assign n16996 = n13696 | n16995 ;
  assign n33447 = ~n16996 ;
  assign n16997 = x17 & n33447 ;
  assign n16998 = n30580 & n16996 ;
  assign n16999 = n16997 | n16998 ;
  assign n17000 = n16992 & n16999 ;
  assign n16973 = n16965 & n16972 ;
  assign n33448 = ~n16973 ;
  assign n17001 = n33448 & n16974 ;
  assign n33449 = ~n17000 ;
  assign n17002 = n33449 & n17001 ;
  assign n33450 = ~n17002 ;
  assign n17003 = n16974 & n33450 ;
  assign n17004 = n16953 | n16960 ;
  assign n33451 = ~n16961 ;
  assign n17005 = n33451 & n17004 ;
  assign n17006 = n17003 & n17005 ;
  assign n17007 = n16961 | n17006 ;
  assign n17009 = n16952 & n17007 ;
  assign n17010 = n16950 | n17009 ;
  assign n17011 = n16934 & n16936 ;
  assign n33452 = ~n17011 ;
  assign n17012 = n16937 & n33452 ;
  assign n33453 = ~n17010 ;
  assign n17014 = n33453 & n17012 ;
  assign n33454 = ~n17014 ;
  assign n17015 = n16937 & n33454 ;
  assign n17016 = n16927 & n17015 ;
  assign n16576 = n16532 & n16575 ;
  assign n17017 = n16532 | n16575 ;
  assign n33455 = ~n16576 ;
  assign n17018 = n33455 & n17017 ;
  assign n17019 = n16927 | n17015 ;
  assign n33456 = ~n17016 ;
  assign n17020 = n33456 & n17019 ;
  assign n17022 = n17018 & n17020 ;
  assign n17023 = n17016 | n17022 ;
  assign n16919 = n16911 & n16918 ;
  assign n33457 = ~n16919 ;
  assign n17024 = n33457 & n16920 ;
  assign n33458 = ~n17023 ;
  assign n17025 = n33458 & n17024 ;
  assign n33459 = ~n17025 ;
  assign n17026 = n16920 & n33459 ;
  assign n33460 = ~n17026 ;
  assign n17028 = n16909 & n33460 ;
  assign n33461 = ~n17028 ;
  assign n17029 = n16908 & n33461 ;
  assign n33462 = ~n17029 ;
  assign n17031 = n16897 & n33462 ;
  assign n33463 = ~n17031 ;
  assign n17032 = n16896 & n33463 ;
  assign n33464 = ~n17032 ;
  assign n17034 = n16885 & n33464 ;
  assign n33465 = ~n17034 ;
  assign n17035 = n16884 & n33465 ;
  assign n33466 = ~n17035 ;
  assign n17037 = n16873 & n33466 ;
  assign n33467 = ~n17037 ;
  assign n17038 = n16871 & n33467 ;
  assign n33468 = ~n17038 ;
  assign n17040 = n16860 & n33468 ;
  assign n33469 = ~n17040 ;
  assign n17041 = n16858 & n33469 ;
  assign n33470 = ~n17041 ;
  assign n17043 = n16847 & n33470 ;
  assign n33471 = ~n17043 ;
  assign n17044 = n16845 & n33471 ;
  assign n17046 = n16834 | n17044 ;
  assign n33472 = ~n16832 ;
  assign n17047 = n33472 & n17046 ;
  assign n17049 = n16821 | n17047 ;
  assign n33473 = ~n16819 ;
  assign n17050 = n33473 & n17049 ;
  assign n17051 = n16809 & n17050 ;
  assign n17052 = n16807 | n17051 ;
  assign n17053 = n16796 | n17052 ;
  assign n33474 = ~n16794 ;
  assign n17054 = n33474 & n17053 ;
  assign n33475 = ~n16774 ;
  assign n16782 = n33475 & n16781 ;
  assign n17055 = n16782 | n16783 ;
  assign n17057 = n17054 | n17055 ;
  assign n33476 = ~n16783 ;
  assign n17058 = n33476 & n17057 ;
  assign n33477 = ~n17058 ;
  assign n17060 = n16772 & n33477 ;
  assign n33478 = ~n17060 ;
  assign n17061 = n16770 & n33478 ;
  assign n17062 = n16751 | n16758 ;
  assign n33479 = ~n16759 ;
  assign n17063 = n33479 & n17062 ;
  assign n17064 = n17061 & n17063 ;
  assign n17065 = n16759 | n17064 ;
  assign n33480 = ~n17065 ;
  assign n17066 = n16749 & n33480 ;
  assign n33481 = ~n17066 ;
  assign n17067 = n16747 & n33481 ;
  assign n33482 = ~n17067 ;
  assign n17069 = n16736 & n33482 ;
  assign n33483 = ~n17069 ;
  assign n17070 = n16734 & n33483 ;
  assign n33484 = ~n17070 ;
  assign n17072 = n16723 & n33484 ;
  assign n33485 = ~n17072 ;
  assign n17073 = n16721 & n33485 ;
  assign n33486 = ~n16701 ;
  assign n16709 = n33486 & n16708 ;
  assign n17074 = n16709 | n16710 ;
  assign n17076 = n17073 | n17074 ;
  assign n33487 = ~n16710 ;
  assign n17077 = n33487 & n17076 ;
  assign n17078 = n16699 & n17077 ;
  assign n17079 = n16697 | n17078 ;
  assign n17080 = n16686 | n17079 ;
  assign n33488 = ~n16684 ;
  assign n17081 = n33488 & n17080 ;
  assign n17083 = n16673 | n17081 ;
  assign n33489 = ~n16671 ;
  assign n17084 = n33489 & n17083 ;
  assign n17086 = n16660 | n17084 ;
  assign n33490 = ~n16660 ;
  assign n17085 = n33490 & n17084 ;
  assign n33491 = ~n17084 ;
  assign n17087 = n16660 & n33491 ;
  assign n17088 = n17085 | n17087 ;
  assign n33492 = ~n16673 ;
  assign n17082 = n33492 & n17081 ;
  assign n33493 = ~n17081 ;
  assign n17089 = n16673 & n33493 ;
  assign n17090 = n17082 | n17089 ;
  assign n17091 = n16686 & n17079 ;
  assign n33494 = ~n17091 ;
  assign n17092 = n17080 & n33494 ;
  assign n33495 = ~n743 ;
  assign n17093 = n33495 & n17092 ;
  assign n33496 = ~n17092 ;
  assign n17094 = n743 & n33496 ;
  assign n17095 = n17093 | n17094 ;
  assign n17096 = n16699 | n17077 ;
  assign n33497 = ~n17078 ;
  assign n17097 = n33497 & n17096 ;
  assign n15269 = n7068 & n32889 ;
  assign n15065 = n7041 & n32856 ;
  assign n15165 = n69 & n32876 ;
  assign n17098 = n15065 | n15165 ;
  assign n17099 = n7017 & n32890 ;
  assign n17100 = n17098 | n17099 ;
  assign n17101 = n15269 | n17100 ;
  assign n17102 = x8 | n17101 ;
  assign n17103 = x8 & n17101 ;
  assign n33498 = ~n17103 ;
  assign n17104 = n17102 & n33498 ;
  assign n17106 = n17097 | n17104 ;
  assign n33499 = ~n17074 ;
  assign n17075 = n17073 & n33499 ;
  assign n33500 = ~n17073 ;
  assign n17107 = n33500 & n17074 ;
  assign n17108 = n17075 | n17107 ;
  assign n14574 = n6272 & n14570 ;
  assign n14522 = n6190 & n32706 ;
  assign n14549 = n6244 & n14536 ;
  assign n17109 = n14522 | n14549 ;
  assign n17110 = n6217 & n32707 ;
  assign n17111 = n17109 | n17110 ;
  assign n17112 = n14574 | n17111 ;
  assign n17113 = x11 | n17112 ;
  assign n17114 = x11 & n17112 ;
  assign n33501 = ~n17114 ;
  assign n17115 = n17113 & n33501 ;
  assign n33502 = ~n17115 ;
  assign n17117 = n17108 & n33502 ;
  assign n17116 = n17108 & n17115 ;
  assign n17118 = n17108 | n17115 ;
  assign n33503 = ~n17116 ;
  assign n17119 = n33503 & n17118 ;
  assign n17071 = n16723 & n17070 ;
  assign n17120 = n16723 | n17070 ;
  assign n33504 = ~n17071 ;
  assign n17121 = n33504 & n17120 ;
  assign n14285 = n5937 & n14283 ;
  assign n13028 = n5994 & n13027 ;
  assign n14149 = n5970 & n14147 ;
  assign n17122 = n13028 | n14149 ;
  assign n17123 = n6018 & n14295 ;
  assign n17124 = n17122 | n17123 ;
  assign n17125 = n14285 | n17124 ;
  assign n17126 = x14 | n17125 ;
  assign n17127 = x14 & n17125 ;
  assign n33505 = ~n17127 ;
  assign n17128 = n17126 & n33505 ;
  assign n17130 = n17121 | n17128 ;
  assign n17068 = n16736 & n17067 ;
  assign n17131 = n16736 | n17067 ;
  assign n33506 = ~n17068 ;
  assign n17132 = n33506 & n17131 ;
  assign n14661 = n5937 & n14655 ;
  assign n13038 = n5970 & n13027 ;
  assign n13065 = n5994 & n32456 ;
  assign n17133 = n13038 | n13065 ;
  assign n17134 = n6018 & n14147 ;
  assign n17135 = n17133 | n17134 ;
  assign n17136 = n14661 | n17135 ;
  assign n17137 = x14 | n17136 ;
  assign n17138 = x14 & n17136 ;
  assign n33507 = ~n17138 ;
  assign n17139 = n17137 & n33507 ;
  assign n17141 = n17132 | n17139 ;
  assign n33508 = ~n16749 ;
  assign n17142 = n33508 & n17065 ;
  assign n17143 = n17066 | n17142 ;
  assign n13115 = n5937 & n32455 ;
  assign n13055 = n5970 & n32456 ;
  assign n13081 = n5994 & n13077 ;
  assign n17144 = n13055 | n13081 ;
  assign n17145 = n6018 & n13027 ;
  assign n17146 = n17144 | n17145 ;
  assign n17147 = n13115 | n17146 ;
  assign n17148 = x14 | n17147 ;
  assign n17149 = x14 & n17147 ;
  assign n33509 = ~n17149 ;
  assign n17150 = n17148 & n33509 ;
  assign n17152 = n17143 | n17150 ;
  assign n33510 = ~n17143 ;
  assign n17151 = n33510 & n17150 ;
  assign n33511 = ~n17150 ;
  assign n17153 = n17143 & n33511 ;
  assign n17154 = n17151 | n17153 ;
  assign n17155 = n17061 | n17063 ;
  assign n33512 = ~n17064 ;
  assign n17156 = n33512 & n17155 ;
  assign n13854 = n5937 & n32557 ;
  assign n12545 = n5994 & n32354 ;
  assign n13078 = n5970 & n13077 ;
  assign n17157 = n12545 | n13078 ;
  assign n17158 = n6018 & n32456 ;
  assign n17159 = n17157 | n17158 ;
  assign n17160 = n13854 | n17159 ;
  assign n17161 = x14 | n17160 ;
  assign n17162 = x14 & n17160 ;
  assign n33513 = ~n17162 ;
  assign n17163 = n17161 & n33513 ;
  assign n17165 = n17156 | n17163 ;
  assign n17164 = n17156 & n17163 ;
  assign n33514 = ~n17164 ;
  assign n17166 = n33514 & n17165 ;
  assign n17059 = n16772 & n17058 ;
  assign n17167 = n16772 | n17058 ;
  assign n33515 = ~n17059 ;
  assign n17168 = n33515 & n17167 ;
  assign n14262 = n5937 & n32641 ;
  assign n12558 = n5970 & n32354 ;
  assign n12574 = n5994 & n12570 ;
  assign n17169 = n12558 | n12574 ;
  assign n17170 = n6018 & n13077 ;
  assign n17171 = n17169 | n17170 ;
  assign n17172 = n14262 | n17171 ;
  assign n17173 = x14 | n17172 ;
  assign n17174 = x14 & n17172 ;
  assign n33516 = ~n17174 ;
  assign n17175 = n17173 & n33516 ;
  assign n17177 = n17168 | n17175 ;
  assign n33517 = ~n17168 ;
  assign n17176 = n33517 & n17175 ;
  assign n33518 = ~n17175 ;
  assign n17178 = n17168 & n33518 ;
  assign n17179 = n17176 | n17178 ;
  assign n33519 = ~n17055 ;
  assign n17056 = n17054 & n33519 ;
  assign n33520 = ~n17054 ;
  assign n17180 = n33520 & n17055 ;
  assign n17181 = n17056 | n17180 ;
  assign n12636 = n5937 & n32356 ;
  assign n12584 = n5970 & n12570 ;
  assign n12596 = n5994 & n12595 ;
  assign n17182 = n12584 | n12596 ;
  assign n17183 = n6018 & n32354 ;
  assign n17184 = n17182 | n17183 ;
  assign n17185 = n12636 | n17184 ;
  assign n17186 = x14 | n17185 ;
  assign n17187 = x14 & n17185 ;
  assign n33521 = ~n17187 ;
  assign n17188 = n17186 & n33521 ;
  assign n33522 = ~n17188 ;
  assign n17190 = n17181 & n33522 ;
  assign n17189 = n17181 & n17188 ;
  assign n17191 = n17181 | n17188 ;
  assign n33523 = ~n17189 ;
  assign n17192 = n33523 & n17191 ;
  assign n17193 = n16796 & n17052 ;
  assign n33524 = ~n17193 ;
  assign n17194 = n17053 & n33524 ;
  assign n12689 = n5937 & n12681 ;
  assign n12143 = n5994 & n32253 ;
  assign n12612 = n5970 & n12595 ;
  assign n17195 = n12143 | n12612 ;
  assign n17196 = n6018 & n12570 ;
  assign n17197 = n17195 | n17196 ;
  assign n17198 = n12689 | n17197 ;
  assign n17199 = x14 | n17198 ;
  assign n17200 = x14 & n17198 ;
  assign n33525 = ~n17200 ;
  assign n17201 = n17199 & n33525 ;
  assign n33526 = ~n17201 ;
  assign n17203 = n17194 & n33526 ;
  assign n17202 = n17194 & n17201 ;
  assign n17204 = n17194 | n17201 ;
  assign n33527 = ~n17202 ;
  assign n17205 = n33527 & n17204 ;
  assign n17206 = n16809 | n17050 ;
  assign n33528 = ~n17051 ;
  assign n17207 = n33528 & n17206 ;
  assign n13829 = n5937 & n32550 ;
  assign n12153 = n5970 & n32253 ;
  assign n12176 = n5994 & n12161 ;
  assign n17208 = n12153 | n12176 ;
  assign n17209 = n6018 & n12595 ;
  assign n17210 = n17208 | n17209 ;
  assign n17211 = n13829 | n17210 ;
  assign n17212 = x14 | n17211 ;
  assign n17213 = x14 & n17211 ;
  assign n33529 = ~n17213 ;
  assign n17214 = n17212 & n33529 ;
  assign n17216 = n17207 | n17214 ;
  assign n17215 = n17207 & n17214 ;
  assign n33530 = ~n17215 ;
  assign n17217 = n33530 & n17216 ;
  assign n12201 = n5937 & n32255 ;
  assign n11856 = n5994 & n32176 ;
  assign n12177 = n5970 & n12161 ;
  assign n17218 = n11856 | n12177 ;
  assign n17219 = n6018 & n32253 ;
  assign n17220 = n17218 | n17219 ;
  assign n17221 = n12201 | n17220 ;
  assign n17222 = x14 | n17221 ;
  assign n17223 = x14 & n17221 ;
  assign n33531 = ~n17223 ;
  assign n17224 = n17222 & n33531 ;
  assign n33532 = ~n16834 ;
  assign n17045 = n33532 & n17044 ;
  assign n33533 = ~n17044 ;
  assign n17225 = n16834 & n33533 ;
  assign n17226 = n17045 | n17225 ;
  assign n12660 = n5937 & n32362 ;
  assign n11446 = n5994 & n11430 ;
  assign n11851 = n5970 & n32176 ;
  assign n17227 = n11446 | n11851 ;
  assign n17228 = n6018 & n12161 ;
  assign n17229 = n17227 | n17228 ;
  assign n17230 = n12660 | n17229 ;
  assign n17231 = x14 | n17230 ;
  assign n17232 = x14 & n17230 ;
  assign n33534 = ~n17232 ;
  assign n17233 = n17231 & n33534 ;
  assign n33535 = ~n17233 ;
  assign n17235 = n17226 & n33535 ;
  assign n17234 = n17226 & n17233 ;
  assign n17236 = n17226 | n17233 ;
  assign n33536 = ~n17234 ;
  assign n17237 = n33536 & n17236 ;
  assign n17042 = n16847 & n17041 ;
  assign n17238 = n16847 | n17041 ;
  assign n33537 = ~n17042 ;
  assign n17239 = n33537 & n17238 ;
  assign n11871 = n5937 & n32178 ;
  assign n11448 = n5970 & n11430 ;
  assign n11492 = n5994 & n11476 ;
  assign n17240 = n11448 | n11492 ;
  assign n17241 = n6018 & n32176 ;
  assign n17242 = n17240 | n17241 ;
  assign n17243 = n11871 | n17242 ;
  assign n17244 = x14 | n17243 ;
  assign n17245 = x14 & n17243 ;
  assign n33538 = ~n17245 ;
  assign n17246 = n17244 & n33538 ;
  assign n17248 = n17239 | n17246 ;
  assign n33539 = ~n17239 ;
  assign n17247 = n33539 & n17246 ;
  assign n33540 = ~n17246 ;
  assign n17249 = n17239 & n33540 ;
  assign n17250 = n17247 | n17249 ;
  assign n17039 = n16860 & n17038 ;
  assign n17251 = n16860 | n17038 ;
  assign n33541 = ~n17039 ;
  assign n17252 = n33541 & n17251 ;
  assign n11473 = n5937 & n11463 ;
  assign n10664 = n5994 & n10656 ;
  assign n11493 = n5970 & n11476 ;
  assign n17253 = n10664 | n11493 ;
  assign n17254 = n6018 & n11430 ;
  assign n17255 = n17253 | n17254 ;
  assign n17256 = n11473 | n17255 ;
  assign n17257 = x14 | n17256 ;
  assign n17258 = x14 & n17256 ;
  assign n33542 = ~n17258 ;
  assign n17259 = n17257 & n33542 ;
  assign n17261 = n17252 | n17259 ;
  assign n33543 = ~n17252 ;
  assign n17260 = n33543 & n17259 ;
  assign n33544 = ~n17259 ;
  assign n17262 = n17252 & n33544 ;
  assign n17263 = n17260 | n17262 ;
  assign n17036 = n16873 & n17035 ;
  assign n17264 = n16873 | n17035 ;
  assign n33545 = ~n17036 ;
  assign n17265 = n33545 & n17264 ;
  assign n11517 = n5937 & n11511 ;
  assign n10674 = n5970 & n10656 ;
  assign n11057 = n5994 & n10679 ;
  assign n17266 = n10674 | n11057 ;
  assign n17267 = n6018 & n11452 ;
  assign n17268 = n17266 | n17267 ;
  assign n17269 = n11517 | n17268 ;
  assign n17270 = x14 | n17269 ;
  assign n17271 = x14 & n17269 ;
  assign n33546 = ~n17271 ;
  assign n17272 = n17270 & n33546 ;
  assign n17274 = n17265 | n17272 ;
  assign n33547 = ~n17265 ;
  assign n17273 = n33547 & n17272 ;
  assign n33548 = ~n17272 ;
  assign n17275 = n17265 & n33548 ;
  assign n17276 = n17273 | n17275 ;
  assign n17033 = n16885 & n17032 ;
  assign n17277 = n16885 | n17032 ;
  assign n33549 = ~n17033 ;
  assign n17278 = n33549 & n17277 ;
  assign n11037 = n5937 & n11030 ;
  assign n10698 = n5994 & n10681 ;
  assign n11058 = n5970 & n10679 ;
  assign n17279 = n10698 | n11058 ;
  assign n17280 = n6018 & n10656 ;
  assign n17281 = n17279 | n17280 ;
  assign n17282 = n11037 | n17281 ;
  assign n17283 = x14 | n17282 ;
  assign n17284 = x14 & n17282 ;
  assign n33550 = ~n17284 ;
  assign n17285 = n17283 & n33550 ;
  assign n17287 = n17278 & n17285 ;
  assign n17030 = n16897 & n17029 ;
  assign n17288 = n16897 | n17029 ;
  assign n33551 = ~n17030 ;
  assign n17289 = n33551 & n17288 ;
  assign n11543 = n5937 & n11536 ;
  assign n10686 = n5970 & n10681 ;
  assign n10724 = n5994 & n10703 ;
  assign n17290 = n10686 | n10724 ;
  assign n17291 = n6018 & n10679 ;
  assign n17292 = n17290 | n17291 ;
  assign n17293 = n11543 | n17292 ;
  assign n17294 = x14 | n17293 ;
  assign n17295 = x14 & n17293 ;
  assign n33552 = ~n17295 ;
  assign n17296 = n17294 & n33552 ;
  assign n17298 = n17289 | n17296 ;
  assign n33553 = ~n17289 ;
  assign n17297 = n33553 & n17296 ;
  assign n33554 = ~n17296 ;
  assign n17299 = n17289 & n33554 ;
  assign n17300 = n17297 | n17299 ;
  assign n17027 = n16909 & n17026 ;
  assign n17301 = n16909 | n17026 ;
  assign n33555 = ~n17027 ;
  assign n17302 = n33555 & n17301 ;
  assign n13166 = n5937 & n13157 ;
  assign n10713 = n5970 & n10703 ;
  assign n10743 = n5994 & n10727 ;
  assign n17303 = n10713 | n10743 ;
  assign n17304 = n6018 & n10681 ;
  assign n17305 = n17303 | n17304 ;
  assign n17306 = n13166 | n17305 ;
  assign n17307 = x14 | n17306 ;
  assign n17308 = x14 & n17306 ;
  assign n33556 = ~n17308 ;
  assign n17309 = n17307 & n33556 ;
  assign n17311 = n17302 | n17309 ;
  assign n33557 = ~n17302 ;
  assign n17310 = n33557 & n17309 ;
  assign n33558 = ~n17309 ;
  assign n17312 = n17302 & n33558 ;
  assign n17313 = n17310 | n17312 ;
  assign n33559 = ~n17024 ;
  assign n17314 = n17023 & n33559 ;
  assign n17315 = n17025 | n17314 ;
  assign n13187 = n5937 & n13182 ;
  assign n10744 = n5970 & n10727 ;
  assign n10769 = n5994 & n31999 ;
  assign n17316 = n10744 | n10769 ;
  assign n17317 = n6018 & n13151 ;
  assign n17318 = n17316 | n17317 ;
  assign n17319 = n13187 | n17318 ;
  assign n33560 = ~n17319 ;
  assign n17320 = x14 & n33560 ;
  assign n17321 = n30547 & n17319 ;
  assign n17322 = n17320 | n17321 ;
  assign n17323 = n17315 | n17322 ;
  assign n17324 = n17315 & n17322 ;
  assign n33561 = ~n17324 ;
  assign n17325 = n17323 & n33561 ;
  assign n33562 = ~n17018 ;
  assign n17021 = n33562 & n17020 ;
  assign n33563 = ~n17020 ;
  assign n17326 = n17018 & n33563 ;
  assign n17327 = n17021 | n17326 ;
  assign n11694 = n5937 & n32125 ;
  assign n10759 = n5970 & n31999 ;
  assign n10789 = n5994 & n10773 ;
  assign n17328 = n10759 | n10789 ;
  assign n17329 = n6018 & n10727 ;
  assign n17330 = n17328 | n17329 ;
  assign n17331 = n11694 | n17330 ;
  assign n17332 = x14 | n17331 ;
  assign n17333 = x14 & n17331 ;
  assign n33564 = ~n17333 ;
  assign n17334 = n17332 & n33564 ;
  assign n17336 = n17327 | n17334 ;
  assign n17335 = n17327 & n17334 ;
  assign n33565 = ~n17335 ;
  assign n17337 = n33565 & n17336 ;
  assign n17013 = n17010 & n17012 ;
  assign n17338 = n17010 | n17012 ;
  assign n33566 = ~n17013 ;
  assign n17339 = n33566 & n17338 ;
  assign n13237 = n5937 & n32477 ;
  assign n10790 = n5970 & n10773 ;
  assign n10810 = n5994 & n31998 ;
  assign n17340 = n10790 | n10810 ;
  assign n17341 = n6018 & n32478 ;
  assign n17342 = n17340 | n17341 ;
  assign n17343 = n13237 | n17342 ;
  assign n17344 = x14 | n17343 ;
  assign n17345 = x14 & n17343 ;
  assign n33567 = ~n17345 ;
  assign n17346 = n17344 & n33567 ;
  assign n17348 = n17339 | n17346 ;
  assign n33568 = ~n17007 ;
  assign n17008 = n16952 & n33568 ;
  assign n33569 = ~n16952 ;
  assign n17349 = n33569 & n17007 ;
  assign n17350 = n17008 | n17349 ;
  assign n13288 = n5937 & n32482 ;
  assign n10797 = n5970 & n31998 ;
  assign n10823 = n5994 & n10818 ;
  assign n17351 = n10797 | n10823 ;
  assign n17352 = n6018 & n13292 ;
  assign n17353 = n17351 | n17352 ;
  assign n17354 = n13288 | n17353 ;
  assign n17355 = x14 | n17354 ;
  assign n17356 = x14 & n17354 ;
  assign n33570 = ~n17356 ;
  assign n17357 = n17355 & n33570 ;
  assign n17359 = n17350 | n17357 ;
  assign n17358 = n17350 & n17357 ;
  assign n33571 = ~n17358 ;
  assign n17360 = n33571 & n17359 ;
  assign n13319 = n5937 & n32488 ;
  assign n10834 = n5970 & n10818 ;
  assign n10859 = n5994 & n10841 ;
  assign n17361 = n10834 | n10859 ;
  assign n17362 = n6018 & n31998 ;
  assign n17363 = n17361 | n17362 ;
  assign n17364 = n13319 | n17363 ;
  assign n17365 = x14 | n17364 ;
  assign n17366 = x14 & n17364 ;
  assign n33572 = ~n17366 ;
  assign n17367 = n17365 & n33572 ;
  assign n17368 = n17003 | n17005 ;
  assign n33573 = ~n17006 ;
  assign n17369 = n33573 & n17368 ;
  assign n17371 = n17367 | n17369 ;
  assign n17370 = n17367 & n17369 ;
  assign n33574 = ~n17370 ;
  assign n17372 = n33574 & n17371 ;
  assign n13389 = n5937 & n13382 ;
  assign n10860 = n5970 & n10841 ;
  assign n10881 = n5994 & n10865 ;
  assign n17373 = n10860 | n10881 ;
  assign n17374 = n6018 & n10818 ;
  assign n17375 = n17373 | n17374 ;
  assign n17376 = n13389 | n17375 ;
  assign n33575 = ~n17376 ;
  assign n17377 = x14 & n33575 ;
  assign n17378 = n30547 & n17376 ;
  assign n17379 = n17377 | n17378 ;
  assign n33576 = ~n17001 ;
  assign n17380 = n17000 & n33576 ;
  assign n17381 = n17002 | n17380 ;
  assign n17383 = n17379 & n17381 ;
  assign n17382 = n17379 | n17381 ;
  assign n33577 = ~n17383 ;
  assign n17384 = n17382 & n33577 ;
  assign n33578 = ~n16533 ;
  assign n16991 = n33578 & n16990 ;
  assign n33579 = ~n16990 ;
  assign n17385 = n16533 & n33579 ;
  assign n17386 = n16991 | n17385 ;
  assign n33580 = ~n16999 ;
  assign n17387 = n33580 & n17386 ;
  assign n33581 = ~n17386 ;
  assign n17388 = n16999 & n33581 ;
  assign n17389 = n17387 | n17388 ;
  assign n13464 = n5937 & n13456 ;
  assign n10876 = n5970 & n10865 ;
  assign n10910 = n5994 & n10892 ;
  assign n17390 = n10876 | n10910 ;
  assign n17391 = n6018 & n10841 ;
  assign n17392 = n17390 | n17391 ;
  assign n17393 = n13464 | n17392 ;
  assign n17394 = x14 | n17393 ;
  assign n17395 = x14 & n17393 ;
  assign n33582 = ~n17395 ;
  assign n17396 = n17394 & n33582 ;
  assign n17397 = n17389 & n17396 ;
  assign n17398 = n17389 | n17396 ;
  assign n33583 = ~n17397 ;
  assign n17399 = n33583 & n17398 ;
  assign n16988 = n16981 & n16987 ;
  assign n33584 = ~n16988 ;
  assign n17400 = n33584 & n16989 ;
  assign n13530 = n5937 & n32502 ;
  assign n10899 = n5970 & n10892 ;
  assign n10934 = n5994 & n32503 ;
  assign n17401 = n10899 | n10934 ;
  assign n17402 = n6018 & n10865 ;
  assign n17403 = n17401 | n17402 ;
  assign n17404 = n13530 | n17403 ;
  assign n33585 = ~n17404 ;
  assign n17405 = x14 & n33585 ;
  assign n17406 = n30547 & n17404 ;
  assign n17407 = n17405 | n17406 ;
  assign n17409 = n17400 & n17407 ;
  assign n33586 = ~n17407 ;
  assign n17408 = n17400 & n33586 ;
  assign n33587 = ~n17400 ;
  assign n17410 = n33587 & n17407 ;
  assign n17411 = n17408 | n17410 ;
  assign n17412 = x17 & n16975 ;
  assign n33588 = ~n16979 ;
  assign n17413 = n33588 & n17412 ;
  assign n33589 = ~n17412 ;
  assign n17414 = n16979 & n33589 ;
  assign n17415 = n17413 | n17414 ;
  assign n13761 = n5937 & n13756 ;
  assign n10935 = n5970 & n32503 ;
  assign n10950 = n5994 & n10940 ;
  assign n17416 = n10935 | n10950 ;
  assign n17417 = n6018 & n10892 ;
  assign n17418 = n17416 | n17417 ;
  assign n17419 = n13761 | n17418 ;
  assign n17420 = x14 | n17419 ;
  assign n17421 = x14 & n17419 ;
  assign n33590 = ~n17421 ;
  assign n17422 = n17420 & n33590 ;
  assign n17424 = n17415 | n17422 ;
  assign n17425 = n5934 & n32507 ;
  assign n14867 = n5937 & n14859 ;
  assign n17426 = n6018 & n31995 ;
  assign n17427 = n5970 & n32507 ;
  assign n17428 = n17426 | n17427 ;
  assign n17429 = n14867 | n17428 ;
  assign n17430 = n17425 | n17429 ;
  assign n17431 = x14 & n17430 ;
  assign n10945 = n6018 & n10940 ;
  assign n17432 = n5970 & n31995 ;
  assign n17433 = n5994 & n32507 ;
  assign n17434 = n17432 | n17433 ;
  assign n17435 = n10945 | n17434 ;
  assign n17436 = n5937 & n13637 ;
  assign n17437 = n17435 | n17436 ;
  assign n17439 = n17431 | n17437 ;
  assign n33591 = ~n17439 ;
  assign n17440 = x14 & n33591 ;
  assign n17442 = n16975 | n17440 ;
  assign n13699 = n5937 & n13690 ;
  assign n10954 = n5970 & n10940 ;
  assign n10976 = n5994 & n31995 ;
  assign n17443 = n10954 | n10976 ;
  assign n17444 = n6018 & n32503 ;
  assign n17445 = n17443 | n17444 ;
  assign n17446 = n13699 | n17445 ;
  assign n33592 = ~n17446 ;
  assign n17447 = x14 & n33592 ;
  assign n17448 = n30547 & n17446 ;
  assign n17449 = n17447 | n17448 ;
  assign n17450 = n17442 & n17449 ;
  assign n17423 = n17415 & n17422 ;
  assign n33593 = ~n17423 ;
  assign n17451 = n33593 & n17424 ;
  assign n33594 = ~n17450 ;
  assign n17452 = n33594 & n17451 ;
  assign n33595 = ~n17452 ;
  assign n17453 = n17424 & n33595 ;
  assign n17455 = n17411 & n17453 ;
  assign n17456 = n17409 | n17455 ;
  assign n17458 = n17399 & n17456 ;
  assign n17459 = n17397 | n17458 ;
  assign n17461 = n17384 & n17459 ;
  assign n17462 = n17383 | n17461 ;
  assign n33596 = ~n17462 ;
  assign n17463 = n17372 & n33596 ;
  assign n33597 = ~n17463 ;
  assign n17465 = n17371 & n33597 ;
  assign n33598 = ~n17465 ;
  assign n17467 = n17360 & n33598 ;
  assign n33599 = ~n17467 ;
  assign n17468 = n17359 & n33599 ;
  assign n17347 = n17339 & n17346 ;
  assign n33600 = ~n17347 ;
  assign n17469 = n33600 & n17348 ;
  assign n33601 = ~n17468 ;
  assign n17471 = n33601 & n17469 ;
  assign n33602 = ~n17471 ;
  assign n17472 = n17348 & n33602 ;
  assign n33603 = ~n17472 ;
  assign n17474 = n17337 & n33603 ;
  assign n33604 = ~n17474 ;
  assign n17475 = n17336 & n33604 ;
  assign n33605 = ~n17475 ;
  assign n17477 = n17325 & n33605 ;
  assign n33606 = ~n17477 ;
  assign n17478 = n17323 & n33606 ;
  assign n33607 = ~n17478 ;
  assign n17480 = n17313 & n33607 ;
  assign n33608 = ~n17480 ;
  assign n17481 = n17311 & n33608 ;
  assign n33609 = ~n17481 ;
  assign n17483 = n17300 & n33609 ;
  assign n33610 = ~n17483 ;
  assign n17484 = n17298 & n33610 ;
  assign n33611 = ~n17278 ;
  assign n17286 = n33611 & n17285 ;
  assign n33612 = ~n17285 ;
  assign n17485 = n17278 & n33612 ;
  assign n17486 = n17286 | n17485 ;
  assign n17487 = n17484 & n17486 ;
  assign n17488 = n17287 | n17487 ;
  assign n33613 = ~n17488 ;
  assign n17489 = n17276 & n33613 ;
  assign n33614 = ~n17489 ;
  assign n17490 = n17274 & n33614 ;
  assign n33615 = ~n17490 ;
  assign n17492 = n17263 & n33615 ;
  assign n33616 = ~n17492 ;
  assign n17493 = n17261 & n33616 ;
  assign n33617 = ~n17493 ;
  assign n17495 = n17250 & n33617 ;
  assign n33618 = ~n17495 ;
  assign n17496 = n17248 & n33618 ;
  assign n17498 = n17237 | n17496 ;
  assign n33619 = ~n17235 ;
  assign n17499 = n33619 & n17498 ;
  assign n17501 = n17224 | n17499 ;
  assign n33620 = ~n16821 ;
  assign n17048 = n33620 & n17047 ;
  assign n33621 = ~n17047 ;
  assign n17502 = n16821 & n33621 ;
  assign n17503 = n17048 | n17502 ;
  assign n17500 = n17224 & n17499 ;
  assign n33622 = ~n17500 ;
  assign n17504 = n33622 & n17501 ;
  assign n17505 = n17503 & n17504 ;
  assign n33623 = ~n17505 ;
  assign n17506 = n17501 & n33623 ;
  assign n33624 = ~n17506 ;
  assign n17508 = n17217 & n33624 ;
  assign n33625 = ~n17508 ;
  assign n17509 = n17216 & n33625 ;
  assign n17511 = n17205 | n17509 ;
  assign n33626 = ~n17203 ;
  assign n17512 = n33626 & n17511 ;
  assign n17514 = n17192 | n17512 ;
  assign n33627 = ~n17190 ;
  assign n17515 = n33627 & n17514 ;
  assign n33628 = ~n17515 ;
  assign n17517 = n17179 & n33628 ;
  assign n33629 = ~n17517 ;
  assign n17518 = n17177 & n33629 ;
  assign n33630 = ~n17518 ;
  assign n17520 = n17166 & n33630 ;
  assign n33631 = ~n17520 ;
  assign n17521 = n17165 & n33631 ;
  assign n33632 = ~n17521 ;
  assign n17523 = n17154 & n33632 ;
  assign n33633 = ~n17523 ;
  assign n17524 = n17152 & n33633 ;
  assign n33634 = ~n17132 ;
  assign n17140 = n33634 & n17139 ;
  assign n33635 = ~n17139 ;
  assign n17525 = n17132 & n33635 ;
  assign n17526 = n17140 | n17525 ;
  assign n33636 = ~n17524 ;
  assign n17527 = n33636 & n17526 ;
  assign n33637 = ~n17527 ;
  assign n17528 = n17141 & n33637 ;
  assign n17129 = n17121 & n17128 ;
  assign n33638 = ~n17129 ;
  assign n17529 = n33638 & n17130 ;
  assign n33639 = ~n17528 ;
  assign n17530 = n33639 & n17529 ;
  assign n33640 = ~n17530 ;
  assign n17531 = n17130 & n33640 ;
  assign n17533 = n17119 | n17531 ;
  assign n33641 = ~n17117 ;
  assign n17534 = n33641 & n17533 ;
  assign n17105 = n17097 & n17104 ;
  assign n33642 = ~n17105 ;
  assign n17535 = n33642 & n17106 ;
  assign n33643 = ~n17534 ;
  assign n17537 = n33643 & n17535 ;
  assign n33644 = ~n17537 ;
  assign n17538 = n17106 & n33644 ;
  assign n17540 = n17095 | n17538 ;
  assign n33645 = ~n17093 ;
  assign n17541 = n33645 & n17540 ;
  assign n33646 = ~n17541 ;
  assign n17543 = n17090 & n33646 ;
  assign n17542 = n17090 & n17541 ;
  assign n17544 = n17090 | n17541 ;
  assign n33647 = ~n17542 ;
  assign n17545 = n33647 & n17544 ;
  assign n33648 = ~n17095 ;
  assign n17539 = n33648 & n17538 ;
  assign n33649 = ~n17538 ;
  assign n17546 = n17095 & n33649 ;
  assign n17547 = n17539 | n17546 ;
  assign n17536 = n17534 & n17535 ;
  assign n17548 = n17534 | n17535 ;
  assign n33650 = ~n17536 ;
  assign n17549 = n33650 & n17548 ;
  assign n15232 = n8156 & n15221 ;
  assign n17550 = n741 | n15232 ;
  assign n33651 = ~n17550 ;
  assign n17551 = x5 & n33651 ;
  assign n17552 = n30053 & n17550 ;
  assign n17553 = n17551 | n17552 ;
  assign n17555 = n17549 & n17553 ;
  assign n15188 = n7068 & n32875 ;
  assign n15063 = n69 & n32856 ;
  assign n15094 = n7041 & n15081 ;
  assign n17556 = n15063 | n15094 ;
  assign n17557 = n7017 & n32876 ;
  assign n17558 = n17556 | n17557 ;
  assign n17559 = n15188 | n17558 ;
  assign n17560 = x8 | n17559 ;
  assign n17561 = x8 & n17559 ;
  assign n33652 = ~n17561 ;
  assign n17562 = n17560 & n33652 ;
  assign n33653 = ~n17119 ;
  assign n17532 = n33653 & n17531 ;
  assign n33654 = ~n17531 ;
  assign n17563 = n17119 & n33654 ;
  assign n17564 = n17532 | n17563 ;
  assign n33655 = ~n17562 ;
  assign n17566 = n33655 & n17564 ;
  assign n17565 = n17562 & n17564 ;
  assign n17567 = n17562 | n17564 ;
  assign n33656 = ~n17565 ;
  assign n17568 = n33656 & n17567 ;
  assign n14688 = n6272 & n32735 ;
  assign n14103 = n6244 & n14101 ;
  assign n14542 = n6190 & n14536 ;
  assign n17569 = n14103 | n14542 ;
  assign n17570 = n6217 & n32706 ;
  assign n17571 = n17569 | n17570 ;
  assign n17572 = n14688 | n17571 ;
  assign n17573 = x11 | n17572 ;
  assign n17574 = x11 & n17572 ;
  assign n33657 = ~n17574 ;
  assign n17575 = n17573 & n33657 ;
  assign n33658 = ~n17529 ;
  assign n17576 = n17528 & n33658 ;
  assign n17577 = n17530 | n17576 ;
  assign n17578 = n17575 | n17577 ;
  assign n17579 = n17575 & n17577 ;
  assign n33659 = ~n17579 ;
  assign n17580 = n17578 & n33659 ;
  assign n33660 = ~n17526 ;
  assign n17581 = n17524 & n33660 ;
  assign n17582 = n17527 | n17581 ;
  assign n14969 = n6272 & n14965 ;
  assign n14102 = n6190 & n14101 ;
  assign n14125 = n6244 & n14124 ;
  assign n17583 = n14102 | n14125 ;
  assign n17584 = n6217 & n14536 ;
  assign n17585 = n17583 | n17584 ;
  assign n17586 = n14969 | n17585 ;
  assign n17587 = x11 | n17586 ;
  assign n17588 = x11 & n17586 ;
  assign n33661 = ~n17588 ;
  assign n17589 = n17587 & n33661 ;
  assign n17591 = n17582 | n17589 ;
  assign n33662 = ~n17582 ;
  assign n17590 = n33662 & n17589 ;
  assign n33663 = ~n17589 ;
  assign n17592 = n17582 & n33663 ;
  assign n17593 = n17590 | n17592 ;
  assign n33664 = ~n17154 ;
  assign n17522 = n33664 & n17521 ;
  assign n17594 = n17522 | n17523 ;
  assign n14186 = n6272 & n14183 ;
  assign n14137 = n6190 & n14124 ;
  assign n14150 = n6244 & n14147 ;
  assign n17595 = n14137 | n14150 ;
  assign n17596 = n6217 & n14196 ;
  assign n17597 = n17595 | n17596 ;
  assign n17598 = n14186 | n17597 ;
  assign n17599 = x11 | n17598 ;
  assign n17600 = x11 & n17598 ;
  assign n33665 = ~n17600 ;
  assign n17601 = n17599 & n33665 ;
  assign n17603 = n17594 | n17601 ;
  assign n33666 = ~n17594 ;
  assign n17602 = n33666 & n17601 ;
  assign n33667 = ~n17601 ;
  assign n17604 = n17594 & n33667 ;
  assign n17605 = n17602 | n17604 ;
  assign n17519 = n17166 & n17518 ;
  assign n17606 = n17166 | n17518 ;
  assign n33668 = ~n17519 ;
  assign n17607 = n33668 & n17606 ;
  assign n14290 = n6272 & n14283 ;
  assign n13029 = n6244 & n13027 ;
  assign n14148 = n6190 & n14147 ;
  assign n17608 = n13029 | n14148 ;
  assign n17609 = n6217 & n14295 ;
  assign n17610 = n17608 | n17609 ;
  assign n17611 = n14290 | n17610 ;
  assign n17612 = x11 | n17611 ;
  assign n17613 = x11 & n17611 ;
  assign n33669 = ~n17613 ;
  assign n17614 = n17612 & n33669 ;
  assign n17616 = n17607 | n17614 ;
  assign n17615 = n17607 & n17614 ;
  assign n33670 = ~n17615 ;
  assign n17617 = n33670 & n17616 ;
  assign n17516 = n17179 & n17515 ;
  assign n17618 = n17179 | n17515 ;
  assign n33671 = ~n17516 ;
  assign n17619 = n33671 & n17618 ;
  assign n14659 = n6272 & n14655 ;
  assign n13044 = n6190 & n13027 ;
  assign n13063 = n6244 & n32456 ;
  assign n17620 = n13044 | n13063 ;
  assign n17621 = n6217 & n14147 ;
  assign n17622 = n17620 | n17621 ;
  assign n17623 = n14659 | n17622 ;
  assign n17624 = x11 | n17623 ;
  assign n17625 = x11 & n17623 ;
  assign n33672 = ~n17625 ;
  assign n17626 = n17624 & n33672 ;
  assign n17628 = n17619 | n17626 ;
  assign n33673 = ~n17619 ;
  assign n17627 = n33673 & n17626 ;
  assign n33674 = ~n17626 ;
  assign n17629 = n17619 & n33674 ;
  assign n17630 = n17627 | n17629 ;
  assign n33675 = ~n17192 ;
  assign n17513 = n33675 & n17512 ;
  assign n33676 = ~n17512 ;
  assign n17631 = n17192 & n33676 ;
  assign n17632 = n17513 | n17631 ;
  assign n13120 = n6272 & n32455 ;
  assign n13053 = n6190 & n32456 ;
  assign n13089 = n6244 & n13077 ;
  assign n17633 = n13053 | n13089 ;
  assign n17634 = n6217 & n13027 ;
  assign n17635 = n17633 | n17634 ;
  assign n17636 = n13120 | n17635 ;
  assign n17637 = x11 | n17636 ;
  assign n17638 = x11 & n17636 ;
  assign n33677 = ~n17638 ;
  assign n17639 = n17637 & n33677 ;
  assign n33678 = ~n17639 ;
  assign n17641 = n17632 & n33678 ;
  assign n17640 = n17632 & n17639 ;
  assign n17642 = n17632 | n17639 ;
  assign n33679 = ~n17640 ;
  assign n17643 = n33679 & n17642 ;
  assign n33680 = ~n17205 ;
  assign n17510 = n33680 & n17509 ;
  assign n33681 = ~n17509 ;
  assign n17644 = n17205 & n33681 ;
  assign n17645 = n17510 | n17644 ;
  assign n13855 = n6272 & n32557 ;
  assign n12547 = n6244 & n32354 ;
  assign n13090 = n6190 & n13077 ;
  assign n17646 = n12547 | n13090 ;
  assign n17647 = n6217 & n32456 ;
  assign n17648 = n17646 | n17647 ;
  assign n17649 = n13855 | n17648 ;
  assign n17650 = x11 | n17649 ;
  assign n17651 = x11 & n17649 ;
  assign n33682 = ~n17651 ;
  assign n17652 = n17650 & n33682 ;
  assign n33683 = ~n17652 ;
  assign n17654 = n17645 & n33683 ;
  assign n17653 = n17645 & n17652 ;
  assign n17655 = n17645 | n17652 ;
  assign n33684 = ~n17653 ;
  assign n17656 = n33684 & n17655 ;
  assign n17507 = n17217 & n17506 ;
  assign n17657 = n17217 | n17506 ;
  assign n33685 = ~n17507 ;
  assign n17658 = n33685 & n17657 ;
  assign n14258 = n6272 & n32641 ;
  assign n12559 = n6190 & n32354 ;
  assign n12589 = n6244 & n12570 ;
  assign n17659 = n12559 | n12589 ;
  assign n17660 = n6217 & n13077 ;
  assign n17661 = n17659 | n17660 ;
  assign n17662 = n14258 | n17661 ;
  assign n17663 = x11 | n17662 ;
  assign n17664 = x11 & n17662 ;
  assign n33686 = ~n17664 ;
  assign n17665 = n17663 & n33686 ;
  assign n17667 = n17658 | n17665 ;
  assign n17666 = n17658 & n17665 ;
  assign n33687 = ~n17666 ;
  assign n17668 = n33687 & n17667 ;
  assign n17669 = n17503 | n17504 ;
  assign n17670 = n33623 & n17669 ;
  assign n12637 = n6272 & n32356 ;
  assign n12583 = n6190 & n12570 ;
  assign n12597 = n6244 & n12595 ;
  assign n17671 = n12583 | n12597 ;
  assign n17672 = n6217 & n32354 ;
  assign n17673 = n17671 | n17672 ;
  assign n17674 = n12637 | n17673 ;
  assign n17675 = x11 | n17674 ;
  assign n17676 = x11 & n17674 ;
  assign n33688 = ~n17676 ;
  assign n17677 = n17675 & n33688 ;
  assign n33689 = ~n17677 ;
  assign n17679 = n17670 & n33689 ;
  assign n17678 = n17670 & n17677 ;
  assign n17680 = n17670 | n17677 ;
  assign n33690 = ~n17678 ;
  assign n17681 = n33690 & n17680 ;
  assign n33691 = ~n17237 ;
  assign n17497 = n33691 & n17496 ;
  assign n33692 = ~n17496 ;
  assign n17682 = n17237 & n33692 ;
  assign n17683 = n17497 | n17682 ;
  assign n12683 = n6272 & n12681 ;
  assign n12150 = n6244 & n32253 ;
  assign n12611 = n6190 & n12595 ;
  assign n17684 = n12150 | n12611 ;
  assign n17685 = n6217 & n12570 ;
  assign n17686 = n17684 | n17685 ;
  assign n17687 = n12683 | n17686 ;
  assign n17688 = x11 | n17687 ;
  assign n17689 = x11 & n17687 ;
  assign n33693 = ~n17689 ;
  assign n17690 = n17688 & n33693 ;
  assign n33694 = ~n17690 ;
  assign n17692 = n17683 & n33694 ;
  assign n17691 = n17683 & n17690 ;
  assign n17693 = n17683 | n17690 ;
  assign n33695 = ~n17691 ;
  assign n17694 = n33695 & n17693 ;
  assign n17494 = n17250 & n17493 ;
  assign n17695 = n17250 | n17493 ;
  assign n33696 = ~n17494 ;
  assign n17696 = n33696 & n17695 ;
  assign n13826 = n6272 & n32550 ;
  assign n12154 = n6190 & n32253 ;
  assign n12175 = n6244 & n12161 ;
  assign n17697 = n12154 | n12175 ;
  assign n17698 = n6217 & n12595 ;
  assign n17699 = n17697 | n17698 ;
  assign n17700 = n13826 | n17699 ;
  assign n17701 = x11 | n17700 ;
  assign n17702 = x11 & n17700 ;
  assign n33697 = ~n17702 ;
  assign n17703 = n17701 & n33697 ;
  assign n17705 = n17696 | n17703 ;
  assign n33698 = ~n17696 ;
  assign n17704 = n33698 & n17703 ;
  assign n33699 = ~n17703 ;
  assign n17706 = n17696 & n33699 ;
  assign n17707 = n17704 | n17706 ;
  assign n17491 = n17263 & n17490 ;
  assign n17708 = n17263 | n17490 ;
  assign n33700 = ~n17491 ;
  assign n17709 = n33700 & n17708 ;
  assign n12199 = n6272 & n32255 ;
  assign n11846 = n6244 & n32176 ;
  assign n12173 = n6190 & n12161 ;
  assign n17710 = n11846 | n12173 ;
  assign n17711 = n6217 & n32253 ;
  assign n17712 = n17710 | n17711 ;
  assign n17713 = n12199 | n17712 ;
  assign n17714 = x11 | n17713 ;
  assign n17715 = x11 & n17713 ;
  assign n33701 = ~n17715 ;
  assign n17716 = n17714 & n33701 ;
  assign n17718 = n17709 | n17716 ;
  assign n33702 = ~n17709 ;
  assign n17717 = n33702 & n17716 ;
  assign n33703 = ~n17716 ;
  assign n17719 = n17709 & n33703 ;
  assign n17720 = n17717 | n17719 ;
  assign n33704 = ~n17276 ;
  assign n17721 = n33704 & n17488 ;
  assign n17722 = n17489 | n17721 ;
  assign n12662 = n6272 & n32362 ;
  assign n11445 = n6244 & n11430 ;
  assign n11857 = n6190 & n32176 ;
  assign n17723 = n11445 | n11857 ;
  assign n17724 = n6217 & n12161 ;
  assign n17725 = n17723 | n17724 ;
  assign n17726 = n12662 | n17725 ;
  assign n17727 = x11 | n17726 ;
  assign n17728 = x11 & n17726 ;
  assign n33705 = ~n17728 ;
  assign n17729 = n17727 & n33705 ;
  assign n17731 = n17722 | n17729 ;
  assign n17730 = n17722 & n17729 ;
  assign n33706 = ~n17730 ;
  assign n17732 = n33706 & n17731 ;
  assign n17733 = n17484 | n17486 ;
  assign n33707 = ~n17487 ;
  assign n17734 = n33707 & n17733 ;
  assign n11878 = n6272 & n32178 ;
  assign n11433 = n6190 & n11430 ;
  assign n11494 = n6244 & n11476 ;
  assign n17735 = n11433 | n11494 ;
  assign n17736 = n6217 & n32176 ;
  assign n17737 = n17735 | n17736 ;
  assign n17738 = n11878 | n17737 ;
  assign n17739 = x11 | n17738 ;
  assign n17740 = x11 & n17738 ;
  assign n33708 = ~n17740 ;
  assign n17741 = n17739 & n33708 ;
  assign n17743 = n17734 | n17741 ;
  assign n17482 = n17300 & n17481 ;
  assign n17744 = n17300 | n17481 ;
  assign n33709 = ~n17482 ;
  assign n17745 = n33709 & n17744 ;
  assign n11474 = n6272 & n11463 ;
  assign n10666 = n6244 & n10656 ;
  assign n11484 = n6190 & n11476 ;
  assign n17746 = n10666 | n11484 ;
  assign n17747 = n6217 & n11430 ;
  assign n17748 = n17746 | n17747 ;
  assign n17749 = n11474 | n17748 ;
  assign n17750 = x11 | n17749 ;
  assign n17751 = x11 & n17749 ;
  assign n33710 = ~n17751 ;
  assign n17752 = n17750 & n33710 ;
  assign n17754 = n17745 | n17752 ;
  assign n33711 = ~n17745 ;
  assign n17753 = n33711 & n17752 ;
  assign n33712 = ~n17752 ;
  assign n17755 = n17745 & n33712 ;
  assign n17756 = n17753 | n17755 ;
  assign n17479 = n17313 & n17478 ;
  assign n17757 = n17313 | n17478 ;
  assign n33713 = ~n17479 ;
  assign n17758 = n33713 & n17757 ;
  assign n11521 = n6272 & n11511 ;
  assign n10675 = n6190 & n10656 ;
  assign n11059 = n6244 & n10679 ;
  assign n17759 = n10675 | n11059 ;
  assign n17760 = n6217 & n11452 ;
  assign n17761 = n17759 | n17760 ;
  assign n17762 = n11521 | n17761 ;
  assign n17763 = x11 | n17762 ;
  assign n17764 = x11 & n17762 ;
  assign n33714 = ~n17764 ;
  assign n17765 = n17763 & n33714 ;
  assign n17767 = n17758 | n17765 ;
  assign n33715 = ~n17758 ;
  assign n17766 = n33715 & n17765 ;
  assign n33716 = ~n17765 ;
  assign n17768 = n17758 & n33716 ;
  assign n17769 = n17766 | n17768 ;
  assign n17476 = n17325 & n17475 ;
  assign n17770 = n17325 | n17475 ;
  assign n33717 = ~n17476 ;
  assign n17771 = n33717 & n17770 ;
  assign n11039 = n6272 & n11030 ;
  assign n10699 = n6244 & n10681 ;
  assign n11046 = n6190 & n10679 ;
  assign n17772 = n10699 | n11046 ;
  assign n17773 = n6217 & n10656 ;
  assign n17774 = n17772 | n17773 ;
  assign n17775 = n11039 | n17774 ;
  assign n17776 = x11 | n17775 ;
  assign n17777 = x11 & n17775 ;
  assign n33718 = ~n17777 ;
  assign n17778 = n17776 & n33718 ;
  assign n17780 = n17771 | n17778 ;
  assign n33719 = ~n17771 ;
  assign n17779 = n33719 & n17778 ;
  assign n33720 = ~n17778 ;
  assign n17781 = n17771 & n33720 ;
  assign n17782 = n17779 | n17781 ;
  assign n17473 = n17337 & n17472 ;
  assign n17783 = n17337 | n17472 ;
  assign n33721 = ~n17473 ;
  assign n17784 = n33721 & n17783 ;
  assign n11545 = n6272 & n11536 ;
  assign n10692 = n6190 & n10681 ;
  assign n10725 = n6244 & n10703 ;
  assign n17785 = n10692 | n10725 ;
  assign n17786 = n6217 & n10679 ;
  assign n17787 = n17785 | n17786 ;
  assign n17788 = n11545 | n17787 ;
  assign n17789 = x11 | n17788 ;
  assign n17790 = x11 & n17788 ;
  assign n33722 = ~n17790 ;
  assign n17791 = n17789 & n33722 ;
  assign n17793 = n17784 | n17791 ;
  assign n33723 = ~n17784 ;
  assign n17792 = n33723 & n17791 ;
  assign n33724 = ~n17791 ;
  assign n17794 = n17784 & n33724 ;
  assign n17795 = n17792 | n17794 ;
  assign n17470 = n17468 & n17469 ;
  assign n17796 = n17468 | n17469 ;
  assign n33725 = ~n17470 ;
  assign n17797 = n33725 & n17796 ;
  assign n13167 = n6272 & n13157 ;
  assign n10705 = n6190 & n10703 ;
  assign n10745 = n6244 & n10727 ;
  assign n17798 = n10705 | n10745 ;
  assign n17799 = n6217 & n10681 ;
  assign n17800 = n17798 | n17799 ;
  assign n17801 = n13167 | n17800 ;
  assign n17802 = x11 | n17801 ;
  assign n17803 = x11 & n17801 ;
  assign n33726 = ~n17803 ;
  assign n17804 = n17802 & n33726 ;
  assign n17806 = n17797 | n17804 ;
  assign n33727 = ~n17797 ;
  assign n17805 = n33727 & n17804 ;
  assign n33728 = ~n17804 ;
  assign n17807 = n17797 & n33728 ;
  assign n17808 = n17805 | n17807 ;
  assign n17466 = n17360 & n17465 ;
  assign n17809 = n17360 | n17465 ;
  assign n33729 = ~n17466 ;
  assign n17810 = n33729 & n17809 ;
  assign n13191 = n6272 & n13182 ;
  assign n10732 = n6190 & n10727 ;
  assign n10767 = n6244 & n31999 ;
  assign n17811 = n10732 | n10767 ;
  assign n17812 = n6217 & n13151 ;
  assign n17813 = n17811 | n17812 ;
  assign n17814 = n13191 | n17813 ;
  assign n17815 = x11 | n17814 ;
  assign n17816 = x11 & n17814 ;
  assign n33730 = ~n17816 ;
  assign n17817 = n17815 & n33730 ;
  assign n17819 = n17810 | n17817 ;
  assign n33731 = ~n17810 ;
  assign n17818 = n33731 & n17817 ;
  assign n33732 = ~n17817 ;
  assign n17820 = n17810 & n33732 ;
  assign n17821 = n17818 | n17820 ;
  assign n17464 = n17372 | n17462 ;
  assign n17822 = n17372 & n17462 ;
  assign n33733 = ~n17822 ;
  assign n17823 = n17464 & n33733 ;
  assign n11693 = n6272 & n32125 ;
  assign n10768 = n6190 & n31999 ;
  assign n10791 = n6244 & n10773 ;
  assign n17824 = n10768 | n10791 ;
  assign n17825 = n6217 & n10727 ;
  assign n17826 = n17824 | n17825 ;
  assign n17827 = n11693 | n17826 ;
  assign n17828 = x11 | n17827 ;
  assign n17829 = x11 & n17827 ;
  assign n33734 = ~n17829 ;
  assign n17830 = n17828 & n33734 ;
  assign n17832 = n17823 | n17830 ;
  assign n33735 = ~n17823 ;
  assign n17831 = n33735 & n17830 ;
  assign n33736 = ~n17830 ;
  assign n17833 = n17823 & n33736 ;
  assign n17834 = n17831 | n17833 ;
  assign n33737 = ~n17459 ;
  assign n17460 = n17384 & n33737 ;
  assign n33738 = ~n17384 ;
  assign n17835 = n33738 & n17459 ;
  assign n17836 = n17460 | n17835 ;
  assign n13238 = n6272 & n32477 ;
  assign n10792 = n6190 & n10773 ;
  assign n10798 = n6244 & n31998 ;
  assign n17837 = n10792 | n10798 ;
  assign n17838 = n6217 & n32478 ;
  assign n17839 = n17837 | n17838 ;
  assign n17840 = n13238 | n17839 ;
  assign n17841 = x11 | n17840 ;
  assign n17842 = x11 & n17840 ;
  assign n33739 = ~n17842 ;
  assign n17843 = n17841 & n33739 ;
  assign n17845 = n17836 | n17843 ;
  assign n17844 = n17836 & n17843 ;
  assign n33740 = ~n17844 ;
  assign n17846 = n33740 & n17845 ;
  assign n33741 = ~n17456 ;
  assign n17457 = n17399 & n33741 ;
  assign n33742 = ~n17399 ;
  assign n17847 = n33742 & n17456 ;
  assign n17848 = n17457 | n17847 ;
  assign n13289 = n6272 & n32482 ;
  assign n10812 = n6190 & n31998 ;
  assign n10837 = n6244 & n10818 ;
  assign n17849 = n10812 | n10837 ;
  assign n17850 = n6217 & n13292 ;
  assign n17851 = n17849 | n17850 ;
  assign n17852 = n13289 | n17851 ;
  assign n17853 = x11 | n17852 ;
  assign n17854 = x11 & n17852 ;
  assign n33743 = ~n17854 ;
  assign n17855 = n17853 & n33743 ;
  assign n17856 = n17848 & n17855 ;
  assign n17857 = n17848 | n17855 ;
  assign n33744 = ~n17856 ;
  assign n17858 = n33744 & n17857 ;
  assign n33745 = ~n17411 ;
  assign n17454 = n33745 & n17453 ;
  assign n33746 = ~n17453 ;
  assign n17859 = n17411 & n33746 ;
  assign n17860 = n17454 | n17859 ;
  assign n13325 = n6272 & n32488 ;
  assign n10835 = n6190 & n10818 ;
  assign n10845 = n6244 & n10841 ;
  assign n17861 = n10835 | n10845 ;
  assign n17862 = n6217 & n31998 ;
  assign n17863 = n17861 | n17862 ;
  assign n17864 = n13325 | n17863 ;
  assign n17865 = x11 | n17864 ;
  assign n17866 = x11 & n17864 ;
  assign n33747 = ~n17866 ;
  assign n17867 = n17865 & n33747 ;
  assign n17869 = n17860 | n17867 ;
  assign n13392 = n6272 & n13382 ;
  assign n10847 = n6190 & n10841 ;
  assign n10882 = n6244 & n10865 ;
  assign n17870 = n10847 | n10882 ;
  assign n17871 = n6217 & n10818 ;
  assign n17872 = n17870 | n17871 ;
  assign n17873 = n13392 | n17872 ;
  assign n17874 = x11 | n17873 ;
  assign n17875 = x11 & n17873 ;
  assign n33748 = ~n17875 ;
  assign n17876 = n17874 & n33748 ;
  assign n33749 = ~n17451 ;
  assign n17877 = n17450 & n33749 ;
  assign n17878 = n17452 | n17877 ;
  assign n17880 = n17876 | n17878 ;
  assign n17879 = n17876 & n17878 ;
  assign n33750 = ~n17879 ;
  assign n17881 = n33750 & n17880 ;
  assign n13466 = n6272 & n13456 ;
  assign n10884 = n6190 & n10865 ;
  assign n10894 = n6244 & n10892 ;
  assign n17882 = n10884 | n10894 ;
  assign n17883 = n6217 & n10841 ;
  assign n17884 = n17882 | n17883 ;
  assign n17885 = n13466 | n17884 ;
  assign n17886 = x11 | n17885 ;
  assign n17887 = x11 & n17885 ;
  assign n33751 = ~n17887 ;
  assign n17888 = n17886 & n33751 ;
  assign n33752 = ~n16975 ;
  assign n17441 = n33752 & n17440 ;
  assign n33753 = ~n17440 ;
  assign n17889 = n16975 & n33753 ;
  assign n17890 = n17441 | n17889 ;
  assign n33754 = ~n17449 ;
  assign n17891 = n33754 & n17890 ;
  assign n33755 = ~n17890 ;
  assign n17892 = n17449 & n33755 ;
  assign n17893 = n17891 | n17892 ;
  assign n17895 = n17888 | n17893 ;
  assign n17894 = n17888 & n17893 ;
  assign n33756 = ~n17894 ;
  assign n17896 = n33756 & n17895 ;
  assign n17438 = n17431 & n17437 ;
  assign n33757 = ~n17438 ;
  assign n17897 = n33757 & n17439 ;
  assign n13535 = n6272 & n32502 ;
  assign n10911 = n6190 & n10892 ;
  assign n10920 = n6244 & n32503 ;
  assign n17898 = n10911 | n10920 ;
  assign n17899 = n6217 & n10865 ;
  assign n17900 = n17898 | n17899 ;
  assign n17901 = n13535 | n17900 ;
  assign n17902 = x11 | n17901 ;
  assign n17903 = x11 & n17901 ;
  assign n33758 = ~n17903 ;
  assign n17904 = n17902 & n33758 ;
  assign n17905 = n17897 & n17904 ;
  assign n17906 = x14 & n17425 ;
  assign n33759 = ~n17429 ;
  assign n17907 = n33759 & n17906 ;
  assign n33760 = ~n17906 ;
  assign n17908 = n17429 & n33760 ;
  assign n17909 = n17907 | n17908 ;
  assign n13765 = n6272 & n13756 ;
  assign n10936 = n6190 & n32503 ;
  assign n10943 = n6244 & n10940 ;
  assign n17910 = n10936 | n10943 ;
  assign n17911 = n6217 & n10892 ;
  assign n17912 = n17910 | n17911 ;
  assign n17913 = n13765 | n17912 ;
  assign n17914 = x11 | n17913 ;
  assign n17915 = x11 & n17913 ;
  assign n33761 = ~n17915 ;
  assign n17916 = n17914 & n33761 ;
  assign n17918 = n17909 | n17916 ;
  assign n17919 = n6188 & n32507 ;
  assign n14864 = n6272 & n14859 ;
  assign n17920 = n6217 & n31995 ;
  assign n17921 = n6190 & n32507 ;
  assign n17922 = n17920 | n17921 ;
  assign n17923 = n14864 | n17922 ;
  assign n17924 = n17919 | n17923 ;
  assign n17925 = x11 & n17924 ;
  assign n10942 = n6217 & n10940 ;
  assign n17926 = n6190 & n31995 ;
  assign n17927 = n6244 & n32507 ;
  assign n17928 = n17926 | n17927 ;
  assign n17929 = n10942 | n17928 ;
  assign n17930 = n6272 & n13637 ;
  assign n17931 = n17929 | n17930 ;
  assign n17933 = n17925 | n17931 ;
  assign n33762 = ~n17933 ;
  assign n17934 = x11 & n33762 ;
  assign n17936 = n17425 | n17934 ;
  assign n13700 = n6272 & n13690 ;
  assign n10963 = n6190 & n10940 ;
  assign n10983 = n6244 & n31995 ;
  assign n17937 = n10963 | n10983 ;
  assign n17938 = n6217 & n32503 ;
  assign n17939 = n17937 | n17938 ;
  assign n17940 = n13700 | n17939 ;
  assign n33763 = ~n17940 ;
  assign n17941 = x11 & n33763 ;
  assign n17942 = n30180 & n17940 ;
  assign n17943 = n17941 | n17942 ;
  assign n17944 = n17936 & n17943 ;
  assign n17917 = n17909 & n17916 ;
  assign n33764 = ~n17917 ;
  assign n17945 = n33764 & n17918 ;
  assign n33765 = ~n17944 ;
  assign n17946 = n33765 & n17945 ;
  assign n33766 = ~n17946 ;
  assign n17947 = n17918 & n33766 ;
  assign n17948 = n17897 | n17904 ;
  assign n33767 = ~n17905 ;
  assign n17949 = n33767 & n17948 ;
  assign n17950 = n17947 & n17949 ;
  assign n17951 = n17905 | n17950 ;
  assign n33768 = ~n17951 ;
  assign n17953 = n17896 & n33768 ;
  assign n33769 = ~n17953 ;
  assign n17954 = n17895 & n33769 ;
  assign n33770 = ~n17954 ;
  assign n17956 = n17881 & n33770 ;
  assign n33771 = ~n17956 ;
  assign n17957 = n17880 & n33771 ;
  assign n17868 = n17860 & n17867 ;
  assign n33772 = ~n17868 ;
  assign n17958 = n33772 & n17869 ;
  assign n33773 = ~n17957 ;
  assign n17960 = n33773 & n17958 ;
  assign n33774 = ~n17960 ;
  assign n17961 = n17869 & n33774 ;
  assign n17963 = n17858 & n17961 ;
  assign n17964 = n17856 | n17963 ;
  assign n33775 = ~n17964 ;
  assign n17965 = n17846 & n33775 ;
  assign n33776 = ~n17965 ;
  assign n17966 = n17845 & n33776 ;
  assign n33777 = ~n17966 ;
  assign n17968 = n17834 & n33777 ;
  assign n33778 = ~n17968 ;
  assign n17969 = n17832 & n33778 ;
  assign n33779 = ~n17969 ;
  assign n17971 = n17821 & n33779 ;
  assign n33780 = ~n17971 ;
  assign n17972 = n17819 & n33780 ;
  assign n33781 = ~n17972 ;
  assign n17974 = n17808 & n33781 ;
  assign n33782 = ~n17974 ;
  assign n17975 = n17806 & n33782 ;
  assign n33783 = ~n17975 ;
  assign n17977 = n17795 & n33783 ;
  assign n33784 = ~n17977 ;
  assign n17978 = n17793 & n33784 ;
  assign n33785 = ~n17978 ;
  assign n17980 = n17782 & n33785 ;
  assign n33786 = ~n17980 ;
  assign n17981 = n17780 & n33786 ;
  assign n33787 = ~n17981 ;
  assign n17983 = n17769 & n33787 ;
  assign n33788 = ~n17983 ;
  assign n17984 = n17767 & n33788 ;
  assign n33789 = ~n17984 ;
  assign n17986 = n17756 & n33789 ;
  assign n33790 = ~n17986 ;
  assign n17987 = n17754 & n33790 ;
  assign n17742 = n17734 & n17741 ;
  assign n33791 = ~n17742 ;
  assign n17988 = n33791 & n17743 ;
  assign n33792 = ~n17987 ;
  assign n17989 = n33792 & n17988 ;
  assign n33793 = ~n17989 ;
  assign n17990 = n17743 & n33793 ;
  assign n33794 = ~n17990 ;
  assign n17992 = n17732 & n33794 ;
  assign n33795 = ~n17992 ;
  assign n17993 = n17731 & n33795 ;
  assign n33796 = ~n17993 ;
  assign n17995 = n17720 & n33796 ;
  assign n33797 = ~n17995 ;
  assign n17996 = n17718 & n33797 ;
  assign n33798 = ~n17996 ;
  assign n17998 = n17707 & n33798 ;
  assign n33799 = ~n17998 ;
  assign n17999 = n17705 & n33799 ;
  assign n18001 = n17694 | n17999 ;
  assign n33800 = ~n17692 ;
  assign n18002 = n33800 & n18001 ;
  assign n18004 = n17681 | n18002 ;
  assign n33801 = ~n17679 ;
  assign n18005 = n33801 & n18004 ;
  assign n33802 = ~n18005 ;
  assign n18007 = n17668 & n33802 ;
  assign n33803 = ~n18007 ;
  assign n18008 = n17667 & n33803 ;
  assign n18010 = n17656 | n18008 ;
  assign n33804 = ~n17654 ;
  assign n18011 = n33804 & n18010 ;
  assign n18013 = n17643 | n18011 ;
  assign n33805 = ~n17641 ;
  assign n18014 = n33805 & n18013 ;
  assign n33806 = ~n18014 ;
  assign n18016 = n17630 & n33806 ;
  assign n33807 = ~n18016 ;
  assign n18017 = n17628 & n33807 ;
  assign n33808 = ~n18017 ;
  assign n18019 = n17617 & n33808 ;
  assign n33809 = ~n18019 ;
  assign n18020 = n17616 & n33809 ;
  assign n33810 = ~n18020 ;
  assign n18022 = n17605 & n33810 ;
  assign n33811 = ~n18022 ;
  assign n18023 = n17603 & n33811 ;
  assign n33812 = ~n18023 ;
  assign n18024 = n17593 & n33812 ;
  assign n33813 = ~n18024 ;
  assign n18025 = n17591 & n33813 ;
  assign n33814 = ~n18025 ;
  assign n18027 = n17580 & n33814 ;
  assign n33815 = ~n18027 ;
  assign n18028 = n17578 & n33815 ;
  assign n18030 = n17568 | n18028 ;
  assign n33816 = ~n17566 ;
  assign n18031 = n33816 & n18030 ;
  assign n17554 = n17549 | n17553 ;
  assign n33817 = ~n17555 ;
  assign n18032 = n17554 & n33817 ;
  assign n18034 = n18031 & n18032 ;
  assign n18035 = n17555 | n18034 ;
  assign n33818 = ~n18035 ;
  assign n18036 = n17547 & n33818 ;
  assign n33819 = ~n17547 ;
  assign n18037 = n33819 & n18035 ;
  assign n18038 = n18036 | n18037 ;
  assign n33820 = ~n18031 ;
  assign n18033 = n33820 & n18032 ;
  assign n33821 = ~n18032 ;
  assign n18039 = n18031 & n33821 ;
  assign n18040 = n18033 | n18039 ;
  assign n15522 = n738 & n15516 ;
  assign n15253 = n8195 & n32890 ;
  assign n18041 = n9052 | n15253 ;
  assign n18042 = n740 & n15221 ;
  assign n18043 = n18041 | n18042 ;
  assign n18044 = n15522 | n18043 ;
  assign n33822 = ~n18044 ;
  assign n18045 = x5 & n33822 ;
  assign n18046 = n30053 & n18044 ;
  assign n18047 = n18045 | n18046 ;
  assign n33823 = ~n17568 ;
  assign n18029 = n33823 & n18028 ;
  assign n33824 = ~n18028 ;
  assign n18048 = n17568 & n33824 ;
  assign n18049 = n18029 | n18048 ;
  assign n33825 = ~n18047 ;
  assign n18050 = n33825 & n18049 ;
  assign n33826 = ~n18049 ;
  assign n18051 = n18047 & n33826 ;
  assign n18052 = n18050 | n18051 ;
  assign n15116 = n7068 & n15111 ;
  assign n14492 = n7041 & n32707 ;
  assign n15092 = n69 & n15081 ;
  assign n18053 = n14492 | n15092 ;
  assign n18054 = n7017 & n32856 ;
  assign n18055 = n18053 | n18054 ;
  assign n18056 = n15116 | n18055 ;
  assign n18057 = x8 | n18056 ;
  assign n18058 = x8 & n18056 ;
  assign n33827 = ~n18058 ;
  assign n18059 = n18057 & n33827 ;
  assign n18026 = n17580 & n18025 ;
  assign n18060 = n17580 | n18025 ;
  assign n33828 = ~n18026 ;
  assign n18061 = n33828 & n18060 ;
  assign n18062 = n18059 | n18061 ;
  assign n18063 = n18059 & n18061 ;
  assign n33829 = ~n18063 ;
  assign n18064 = n18062 & n33829 ;
  assign n33830 = ~n17593 ;
  assign n18065 = n33830 & n18023 ;
  assign n18066 = n18024 | n18065 ;
  assign n15292 = n7068 & n15288 ;
  assign n14491 = n69 & n32707 ;
  assign n14519 = n7041 & n32706 ;
  assign n18067 = n14491 | n14519 ;
  assign n18068 = n7017 & n15081 ;
  assign n18069 = n18067 | n18068 ;
  assign n18070 = n15292 | n18069 ;
  assign n18071 = x8 | n18070 ;
  assign n18072 = x8 & n18070 ;
  assign n33831 = ~n18072 ;
  assign n18073 = n18071 & n33831 ;
  assign n18075 = n18066 | n18073 ;
  assign n33832 = ~n18066 ;
  assign n18074 = n33832 & n18073 ;
  assign n33833 = ~n18073 ;
  assign n18076 = n18066 & n33833 ;
  assign n18077 = n18074 | n18076 ;
  assign n18021 = n17605 & n18020 ;
  assign n18078 = n17605 | n18020 ;
  assign n33834 = ~n18021 ;
  assign n18079 = n33834 & n18078 ;
  assign n14572 = n7068 & n14570 ;
  assign n14525 = n69 & n32706 ;
  assign n14541 = n7041 & n14536 ;
  assign n18080 = n14525 | n14541 ;
  assign n18081 = n7017 & n32707 ;
  assign n18082 = n18080 | n18081 ;
  assign n18083 = n14572 | n18082 ;
  assign n18084 = x8 | n18083 ;
  assign n18085 = x8 & n18083 ;
  assign n33835 = ~n18085 ;
  assign n18086 = n18084 & n33835 ;
  assign n18088 = n18079 | n18086 ;
  assign n33836 = ~n18079 ;
  assign n18087 = n33836 & n18086 ;
  assign n33837 = ~n18086 ;
  assign n18089 = n18079 & n33837 ;
  assign n18090 = n18087 | n18089 ;
  assign n18018 = n17617 & n18017 ;
  assign n18091 = n17617 | n18017 ;
  assign n33838 = ~n18018 ;
  assign n18092 = n33838 & n18091 ;
  assign n14686 = n7068 & n32735 ;
  assign n14114 = n7041 & n14101 ;
  assign n14539 = n69 & n14536 ;
  assign n18093 = n14114 | n14539 ;
  assign n18094 = n7017 & n32706 ;
  assign n18095 = n18093 | n18094 ;
  assign n18096 = n14686 | n18095 ;
  assign n18097 = x8 | n18096 ;
  assign n18098 = x8 & n18096 ;
  assign n33839 = ~n18098 ;
  assign n18099 = n18097 & n33839 ;
  assign n18101 = n18092 | n18099 ;
  assign n18100 = n18092 & n18099 ;
  assign n33840 = ~n18100 ;
  assign n18102 = n33840 & n18101 ;
  assign n18015 = n17630 & n18014 ;
  assign n18103 = n17630 | n18014 ;
  assign n33841 = ~n18015 ;
  assign n18104 = n33841 & n18103 ;
  assign n14971 = n7068 & n14965 ;
  assign n14106 = n69 & n14101 ;
  assign n14132 = n7041 & n14124 ;
  assign n18105 = n14106 | n14132 ;
  assign n18106 = n7017 & n14536 ;
  assign n18107 = n18105 | n18106 ;
  assign n18108 = n14971 | n18107 ;
  assign n18109 = x8 | n18108 ;
  assign n18110 = x8 & n18108 ;
  assign n33842 = ~n18110 ;
  assign n18111 = n18109 & n33842 ;
  assign n18113 = n18104 | n18111 ;
  assign n33843 = ~n18104 ;
  assign n18112 = n33843 & n18111 ;
  assign n33844 = ~n18111 ;
  assign n18114 = n18104 & n33844 ;
  assign n18115 = n18112 | n18114 ;
  assign n33845 = ~n17643 ;
  assign n18012 = n33845 & n18011 ;
  assign n33846 = ~n18011 ;
  assign n18116 = n17643 & n33846 ;
  assign n18117 = n18012 | n18116 ;
  assign n14189 = n7068 & n14183 ;
  assign n14128 = n69 & n14124 ;
  assign n14159 = n7041 & n14147 ;
  assign n18118 = n14128 | n14159 ;
  assign n18119 = n7017 & n14196 ;
  assign n18120 = n18118 | n18119 ;
  assign n18121 = n14189 | n18120 ;
  assign n18122 = x8 | n18121 ;
  assign n18123 = x8 & n18121 ;
  assign n33847 = ~n18123 ;
  assign n18124 = n18122 & n33847 ;
  assign n33848 = ~n18124 ;
  assign n18126 = n18117 & n33848 ;
  assign n33849 = ~n18117 ;
  assign n18125 = n33849 & n18124 ;
  assign n18127 = n18125 | n18126 ;
  assign n33850 = ~n17656 ;
  assign n18009 = n33850 & n18008 ;
  assign n33851 = ~n18008 ;
  assign n18128 = n17656 & n33851 ;
  assign n18129 = n18009 | n18128 ;
  assign n14291 = n7068 & n14283 ;
  assign n13037 = n7041 & n13027 ;
  assign n14161 = n69 & n14147 ;
  assign n18130 = n13037 | n14161 ;
  assign n18131 = n7017 & n14295 ;
  assign n18132 = n18130 | n18131 ;
  assign n18133 = n14291 | n18132 ;
  assign n18134 = x8 | n18133 ;
  assign n18135 = x8 & n18133 ;
  assign n33852 = ~n18135 ;
  assign n18136 = n18134 & n33852 ;
  assign n33853 = ~n18136 ;
  assign n18138 = n18129 & n33853 ;
  assign n33854 = ~n18129 ;
  assign n18137 = n33854 & n18136 ;
  assign n18139 = n18137 | n18138 ;
  assign n18006 = n17668 & n18005 ;
  assign n18140 = n17668 | n18005 ;
  assign n33855 = ~n18006 ;
  assign n18141 = n33855 & n18140 ;
  assign n14657 = n7068 & n14655 ;
  assign n13030 = n69 & n13027 ;
  assign n13064 = n7041 & n32456 ;
  assign n18142 = n13030 | n13064 ;
  assign n18143 = n7017 & n14147 ;
  assign n18144 = n18142 | n18143 ;
  assign n18145 = n14657 | n18144 ;
  assign n18146 = x8 | n18145 ;
  assign n18147 = x8 & n18145 ;
  assign n33856 = ~n18147 ;
  assign n18148 = n18146 & n33856 ;
  assign n18150 = n18141 | n18148 ;
  assign n18149 = n18141 & n18148 ;
  assign n33857 = ~n18149 ;
  assign n18151 = n33857 & n18150 ;
  assign n33858 = ~n18002 ;
  assign n18003 = n17681 & n33858 ;
  assign n33859 = ~n17681 ;
  assign n18152 = n33859 & n18002 ;
  assign n18153 = n18003 | n18152 ;
  assign n13122 = n7068 & n32455 ;
  assign n13068 = n69 & n32456 ;
  assign n13091 = n7041 & n13077 ;
  assign n18154 = n13068 | n13091 ;
  assign n18155 = n7017 & n13027 ;
  assign n18156 = n18154 | n18155 ;
  assign n18157 = n13122 | n18156 ;
  assign n18158 = x8 | n18157 ;
  assign n18159 = x8 & n18157 ;
  assign n33860 = ~n18159 ;
  assign n18160 = n18158 & n33860 ;
  assign n33861 = ~n18160 ;
  assign n18162 = n18153 & n33861 ;
  assign n18161 = n18153 & n18160 ;
  assign n18163 = n18153 | n18160 ;
  assign n33862 = ~n18161 ;
  assign n18164 = n33862 & n18163 ;
  assign n33863 = ~n17694 ;
  assign n18000 = n33863 & n17999 ;
  assign n33864 = ~n17999 ;
  assign n18165 = n17694 & n33864 ;
  assign n18166 = n18000 | n18165 ;
  assign n13856 = n7068 & n32557 ;
  assign n12560 = n7041 & n32354 ;
  assign n13092 = n69 & n13077 ;
  assign n18167 = n12560 | n13092 ;
  assign n18168 = n7017 & n32456 ;
  assign n18169 = n18167 | n18168 ;
  assign n18170 = n13856 | n18169 ;
  assign n18171 = x8 | n18170 ;
  assign n18172 = x8 & n18170 ;
  assign n33865 = ~n18172 ;
  assign n18173 = n18171 & n33865 ;
  assign n33866 = ~n18173 ;
  assign n18175 = n18166 & n33866 ;
  assign n33867 = ~n18166 ;
  assign n18174 = n33867 & n18173 ;
  assign n18176 = n18174 | n18175 ;
  assign n17997 = n17707 & n17996 ;
  assign n18177 = n17707 | n17996 ;
  assign n33868 = ~n17997 ;
  assign n18178 = n33868 & n18177 ;
  assign n14263 = n7068 & n32641 ;
  assign n12562 = n69 & n32354 ;
  assign n12577 = n7041 & n12570 ;
  assign n18179 = n12562 | n12577 ;
  assign n18180 = n7017 & n13077 ;
  assign n18181 = n18179 | n18180 ;
  assign n18182 = n14263 | n18181 ;
  assign n18183 = x8 | n18182 ;
  assign n18184 = x8 & n18182 ;
  assign n33869 = ~n18184 ;
  assign n18185 = n18183 & n33869 ;
  assign n18187 = n18178 | n18185 ;
  assign n18186 = n18178 & n18185 ;
  assign n33870 = ~n18186 ;
  assign n18188 = n33870 & n18187 ;
  assign n12634 = n7068 & n32356 ;
  assign n12590 = n69 & n12570 ;
  assign n12606 = n7041 & n12595 ;
  assign n18189 = n12590 | n12606 ;
  assign n18190 = n7017 & n32354 ;
  assign n18191 = n18189 | n18190 ;
  assign n18192 = n12634 | n18191 ;
  assign n18193 = x8 | n18192 ;
  assign n18194 = x8 & n18192 ;
  assign n33871 = ~n18194 ;
  assign n18195 = n18193 & n33871 ;
  assign n17994 = n17720 & n17993 ;
  assign n18196 = n17720 | n17993 ;
  assign n33872 = ~n17994 ;
  assign n18197 = n33872 & n18196 ;
  assign n18198 = n18195 | n18197 ;
  assign n18199 = n18195 & n18197 ;
  assign n33873 = ~n18199 ;
  assign n18200 = n18198 & n33873 ;
  assign n17991 = n17732 & n17990 ;
  assign n18201 = n17732 | n17990 ;
  assign n33874 = ~n17991 ;
  assign n18202 = n33874 & n18201 ;
  assign n12690 = n7068 & n12681 ;
  assign n12155 = n7041 & n32253 ;
  assign n12613 = n69 & n12595 ;
  assign n18203 = n12155 | n12613 ;
  assign n18204 = n7017 & n12570 ;
  assign n18205 = n18203 | n18204 ;
  assign n18206 = n12690 | n18205 ;
  assign n18207 = x8 | n18206 ;
  assign n18208 = x8 & n18206 ;
  assign n33875 = ~n18208 ;
  assign n18209 = n18207 & n33875 ;
  assign n18211 = n18202 | n18209 ;
  assign n18210 = n18202 & n18209 ;
  assign n33876 = ~n18210 ;
  assign n18212 = n33876 & n18211 ;
  assign n33877 = ~n17988 ;
  assign n18213 = n17987 & n33877 ;
  assign n18214 = n17989 | n18213 ;
  assign n13830 = n7068 & n32550 ;
  assign n12152 = n69 & n32253 ;
  assign n12178 = n7041 & n12161 ;
  assign n18215 = n12152 | n12178 ;
  assign n18216 = n7017 & n12595 ;
  assign n18217 = n18215 | n18216 ;
  assign n18218 = n13830 | n18217 ;
  assign n18219 = x8 | n18218 ;
  assign n18220 = x8 & n18218 ;
  assign n33878 = ~n18220 ;
  assign n18221 = n18219 & n33878 ;
  assign n18223 = n18214 | n18221 ;
  assign n18222 = n18214 & n18221 ;
  assign n33879 = ~n18222 ;
  assign n18224 = n33879 & n18223 ;
  assign n17985 = n17756 & n17984 ;
  assign n18225 = n17756 | n17984 ;
  assign n33880 = ~n17985 ;
  assign n18226 = n33880 & n18225 ;
  assign n12200 = n7068 & n32255 ;
  assign n11847 = n7041 & n32176 ;
  assign n12180 = n69 & n12161 ;
  assign n18227 = n11847 | n12180 ;
  assign n18228 = n7017 & n32253 ;
  assign n18229 = n18227 | n18228 ;
  assign n18230 = n12200 | n18229 ;
  assign n18231 = x8 | n18230 ;
  assign n18232 = x8 & n18230 ;
  assign n33881 = ~n18232 ;
  assign n18233 = n18231 & n33881 ;
  assign n18234 = n18226 & n18233 ;
  assign n17982 = n17769 | n17981 ;
  assign n18235 = n17769 & n17981 ;
  assign n33882 = ~n18235 ;
  assign n18236 = n17982 & n33882 ;
  assign n12664 = n7068 & n32362 ;
  assign n11447 = n7041 & n11430 ;
  assign n11858 = n69 & n32176 ;
  assign n18237 = n11447 | n11858 ;
  assign n18238 = n7017 & n12161 ;
  assign n18239 = n18237 | n18238 ;
  assign n18240 = n12664 | n18239 ;
  assign n18241 = x8 | n18240 ;
  assign n18242 = x8 & n18240 ;
  assign n33883 = ~n18242 ;
  assign n18243 = n18241 & n33883 ;
  assign n18245 = n18236 | n18243 ;
  assign n18244 = n18236 & n18243 ;
  assign n33884 = ~n18244 ;
  assign n18246 = n33884 & n18245 ;
  assign n33885 = ~n17782 ;
  assign n17979 = n33885 & n17978 ;
  assign n18247 = n17979 | n17980 ;
  assign n11879 = n7068 & n32178 ;
  assign n11449 = n69 & n11430 ;
  assign n11485 = n7041 & n11476 ;
  assign n18248 = n11449 | n11485 ;
  assign n18249 = n7017 & n32176 ;
  assign n18250 = n18248 | n18249 ;
  assign n18251 = n11879 | n18250 ;
  assign n18252 = x8 | n18251 ;
  assign n18253 = x8 & n18251 ;
  assign n33886 = ~n18253 ;
  assign n18254 = n18252 & n33886 ;
  assign n18256 = n18247 | n18254 ;
  assign n33887 = ~n18247 ;
  assign n18255 = n33887 & n18254 ;
  assign n33888 = ~n18254 ;
  assign n18257 = n18247 & n33888 ;
  assign n18258 = n18255 | n18257 ;
  assign n17976 = n17795 & n17975 ;
  assign n18259 = n17795 | n17975 ;
  assign n33889 = ~n17976 ;
  assign n18260 = n33889 & n18259 ;
  assign n11465 = n7068 & n11463 ;
  assign n10676 = n7041 & n10656 ;
  assign n11495 = n69 & n11476 ;
  assign n18261 = n10676 | n11495 ;
  assign n18262 = n7017 & n11430 ;
  assign n18263 = n18261 | n18262 ;
  assign n18264 = n11465 | n18263 ;
  assign n18265 = x8 | n18264 ;
  assign n18266 = x8 & n18264 ;
  assign n33890 = ~n18266 ;
  assign n18267 = n18265 & n33890 ;
  assign n18269 = n18260 | n18267 ;
  assign n33891 = ~n18260 ;
  assign n18268 = n33891 & n18267 ;
  assign n33892 = ~n18267 ;
  assign n18270 = n18260 & n33892 ;
  assign n18271 = n18268 | n18270 ;
  assign n17973 = n17808 & n17972 ;
  assign n18272 = n17808 | n17972 ;
  assign n33893 = ~n17973 ;
  assign n18273 = n33893 & n18272 ;
  assign n11518 = n7068 & n11511 ;
  assign n10662 = n69 & n10656 ;
  assign n11054 = n7041 & n10679 ;
  assign n18274 = n10662 | n11054 ;
  assign n18275 = n7017 & n11452 ;
  assign n18276 = n18274 | n18275 ;
  assign n18277 = n11518 | n18276 ;
  assign n18278 = x8 | n18277 ;
  assign n18279 = x8 & n18277 ;
  assign n33894 = ~n18279 ;
  assign n18280 = n18278 & n33894 ;
  assign n18282 = n18273 | n18280 ;
  assign n33895 = ~n18273 ;
  assign n18281 = n33895 & n18280 ;
  assign n33896 = ~n18280 ;
  assign n18283 = n18273 & n33896 ;
  assign n18284 = n18281 | n18283 ;
  assign n17970 = n17821 & n17969 ;
  assign n18285 = n17821 | n17969 ;
  assign n33897 = ~n17970 ;
  assign n18286 = n33897 & n18285 ;
  assign n11035 = n7068 & n11030 ;
  assign n10697 = n7041 & n10681 ;
  assign n11061 = n69 & n10679 ;
  assign n18287 = n10697 | n11061 ;
  assign n18288 = n7017 & n10656 ;
  assign n18289 = n18287 | n18288 ;
  assign n18290 = n11035 | n18289 ;
  assign n18291 = x8 | n18290 ;
  assign n18292 = x8 & n18290 ;
  assign n33898 = ~n18292 ;
  assign n18293 = n18291 & n33898 ;
  assign n18294 = n18286 & n18293 ;
  assign n17967 = n17834 & n17966 ;
  assign n18295 = n17834 | n17966 ;
  assign n33899 = ~n17967 ;
  assign n18296 = n33899 & n18295 ;
  assign n11544 = n7068 & n11536 ;
  assign n10700 = n69 & n10681 ;
  assign n10714 = n7041 & n10703 ;
  assign n18297 = n10700 | n10714 ;
  assign n18298 = n7017 & n10679 ;
  assign n18299 = n18297 | n18298 ;
  assign n18300 = n11544 | n18299 ;
  assign n18301 = x8 | n18300 ;
  assign n18302 = x8 & n18300 ;
  assign n33900 = ~n18302 ;
  assign n18303 = n18301 & n33900 ;
  assign n18305 = n18296 | n18303 ;
  assign n33901 = ~n18296 ;
  assign n18304 = n33901 & n18303 ;
  assign n33902 = ~n18303 ;
  assign n18306 = n18296 & n33902 ;
  assign n18307 = n18304 | n18306 ;
  assign n33903 = ~n17846 ;
  assign n18308 = n33903 & n17964 ;
  assign n18309 = n17965 | n18308 ;
  assign n13165 = n7068 & n13157 ;
  assign n10706 = n69 & n10703 ;
  assign n10746 = n7041 & n10727 ;
  assign n18310 = n10706 | n10746 ;
  assign n18311 = n7017 & n10681 ;
  assign n18312 = n18310 | n18311 ;
  assign n18313 = n13165 | n18312 ;
  assign n18314 = x8 | n18313 ;
  assign n18315 = x8 & n18313 ;
  assign n33904 = ~n18315 ;
  assign n18316 = n18314 & n33904 ;
  assign n18318 = n18309 | n18316 ;
  assign n33905 = ~n18309 ;
  assign n18317 = n33905 & n18316 ;
  assign n33906 = ~n18316 ;
  assign n18319 = n18309 & n33906 ;
  assign n18320 = n18317 | n18319 ;
  assign n33907 = ~n17858 ;
  assign n17962 = n33907 & n17961 ;
  assign n33908 = ~n17961 ;
  assign n18321 = n17858 & n33908 ;
  assign n18322 = n17962 | n18321 ;
  assign n13189 = n7068 & n13182 ;
  assign n10736 = n69 & n10727 ;
  assign n10755 = n7041 & n31999 ;
  assign n18323 = n10736 | n10755 ;
  assign n18324 = n7017 & n13151 ;
  assign n18325 = n18323 | n18324 ;
  assign n18326 = n13189 | n18325 ;
  assign n18327 = x8 | n18326 ;
  assign n18328 = x8 & n18326 ;
  assign n33909 = ~n18328 ;
  assign n18329 = n18327 & n33909 ;
  assign n18331 = n18322 | n18329 ;
  assign n17959 = n17957 & n17958 ;
  assign n18332 = n17957 | n17958 ;
  assign n33910 = ~n17959 ;
  assign n18333 = n33910 & n18332 ;
  assign n11695 = n7068 & n32125 ;
  assign n10765 = n69 & n31999 ;
  assign n10781 = n7041 & n10773 ;
  assign n18334 = n10765 | n10781 ;
  assign n18335 = n7017 & n10727 ;
  assign n18336 = n18334 | n18335 ;
  assign n18337 = n11695 | n18336 ;
  assign n18338 = x8 | n18337 ;
  assign n18339 = x8 & n18337 ;
  assign n33911 = ~n18339 ;
  assign n18340 = n18338 & n33911 ;
  assign n18342 = n18333 | n18340 ;
  assign n33912 = ~n18333 ;
  assign n18341 = n33912 & n18340 ;
  assign n33913 = ~n18340 ;
  assign n18343 = n18333 & n33913 ;
  assign n18344 = n18341 | n18343 ;
  assign n13231 = n7068 & n32477 ;
  assign n10780 = n69 & n10773 ;
  assign n10813 = n7041 & n31998 ;
  assign n18345 = n10780 | n10813 ;
  assign n18346 = n7017 & n32478 ;
  assign n18347 = n18345 | n18346 ;
  assign n18348 = n13231 | n18347 ;
  assign n33914 = ~n18348 ;
  assign n18349 = x8 & n33914 ;
  assign n18350 = n30185 & n18348 ;
  assign n18351 = n18349 | n18350 ;
  assign n17955 = n17881 & n17954 ;
  assign n18352 = n17881 | n17954 ;
  assign n33915 = ~n17955 ;
  assign n18353 = n33915 & n18352 ;
  assign n18354 = n18351 | n18353 ;
  assign n18355 = n18351 & n18353 ;
  assign n33916 = ~n18355 ;
  assign n18356 = n18354 & n33916 ;
  assign n17952 = n17896 | n17951 ;
  assign n18357 = n17896 & n17951 ;
  assign n33917 = ~n18357 ;
  assign n18358 = n17952 & n33917 ;
  assign n13285 = n7068 & n32482 ;
  assign n10814 = n69 & n31998 ;
  assign n10836 = n7041 & n10818 ;
  assign n18359 = n10814 | n10836 ;
  assign n18360 = n7017 & n13292 ;
  assign n18361 = n18359 | n18360 ;
  assign n18362 = n13285 | n18361 ;
  assign n18363 = x8 | n18362 ;
  assign n18364 = x8 & n18362 ;
  assign n33918 = ~n18364 ;
  assign n18365 = n18363 & n33918 ;
  assign n18367 = n18358 | n18365 ;
  assign n18366 = n18358 & n18365 ;
  assign n33919 = ~n18366 ;
  assign n18368 = n33919 & n18367 ;
  assign n13326 = n7068 & n32488 ;
  assign n10833 = n69 & n10818 ;
  assign n10861 = n7041 & n10841 ;
  assign n18369 = n10833 | n10861 ;
  assign n18370 = n7017 & n31998 ;
  assign n18371 = n18369 | n18370 ;
  assign n18372 = n13326 | n18371 ;
  assign n18373 = x8 | n18372 ;
  assign n18374 = x8 & n18372 ;
  assign n33920 = ~n18374 ;
  assign n18375 = n18373 & n33920 ;
  assign n18376 = n17947 | n17949 ;
  assign n33921 = ~n17950 ;
  assign n18377 = n33921 & n18376 ;
  assign n18379 = n18375 | n18377 ;
  assign n18378 = n18375 & n18377 ;
  assign n33922 = ~n18378 ;
  assign n18380 = n33922 & n18379 ;
  assign n13386 = n7068 & n13382 ;
  assign n10853 = n69 & n10841 ;
  assign n10885 = n7041 & n10865 ;
  assign n18381 = n10853 | n10885 ;
  assign n18382 = n7017 & n10818 ;
  assign n18383 = n18381 | n18382 ;
  assign n18384 = n13386 | n18383 ;
  assign n18385 = x8 | n18384 ;
  assign n18386 = x8 & n18384 ;
  assign n33923 = ~n18386 ;
  assign n18387 = n18385 & n33923 ;
  assign n33924 = ~n17945 ;
  assign n18388 = n17944 & n33924 ;
  assign n18389 = n17946 | n18388 ;
  assign n18391 = n18387 | n18389 ;
  assign n33925 = ~n18389 ;
  assign n18390 = n18387 & n33925 ;
  assign n33926 = ~n18387 ;
  assign n18392 = n33926 & n18389 ;
  assign n18393 = n18390 | n18392 ;
  assign n33927 = ~n17425 ;
  assign n17935 = n33927 & n17934 ;
  assign n33928 = ~n17934 ;
  assign n18394 = n17425 & n33928 ;
  assign n18395 = n17935 | n18394 ;
  assign n33929 = ~n17943 ;
  assign n18396 = n33929 & n18395 ;
  assign n33930 = ~n18395 ;
  assign n18397 = n17943 & n33930 ;
  assign n18398 = n18396 | n18397 ;
  assign n13461 = n7068 & n13456 ;
  assign n10886 = n69 & n10865 ;
  assign n10912 = n7041 & n10892 ;
  assign n18399 = n10886 | n10912 ;
  assign n18400 = n7017 & n10841 ;
  assign n18401 = n18399 | n18400 ;
  assign n18402 = n13461 | n18401 ;
  assign n18403 = x8 | n18402 ;
  assign n18404 = x8 & n18402 ;
  assign n33931 = ~n18404 ;
  assign n18405 = n18403 & n33931 ;
  assign n18406 = n18398 & n18405 ;
  assign n18407 = n18398 | n18405 ;
  assign n33932 = ~n18406 ;
  assign n18408 = n33932 & n18407 ;
  assign n17932 = n17925 & n17931 ;
  assign n33933 = ~n17932 ;
  assign n18409 = n33933 & n17933 ;
  assign n13526 = n7068 & n32502 ;
  assign n10913 = n69 & n10892 ;
  assign n10925 = n7041 & n32503 ;
  assign n18410 = n10913 | n10925 ;
  assign n18411 = n7017 & n10865 ;
  assign n18412 = n18410 | n18411 ;
  assign n18413 = n13526 | n18412 ;
  assign n18414 = x8 | n18413 ;
  assign n18415 = x8 & n18413 ;
  assign n33934 = ~n18415 ;
  assign n18416 = n18414 & n33934 ;
  assign n18418 = n18409 | n18416 ;
  assign n18417 = n18409 & n18416 ;
  assign n33935 = ~n18417 ;
  assign n18419 = n33935 & n18418 ;
  assign n18420 = n67 & n32507 ;
  assign n18421 = x8 & n18420 ;
  assign n14866 = n7068 & n14859 ;
  assign n18422 = n7017 & n31995 ;
  assign n18423 = n69 & n32507 ;
  assign n18424 = n18422 | n18423 ;
  assign n18425 = n14866 | n18424 ;
  assign n18426 = n18421 | n18425 ;
  assign n10941 = n7017 & n10940 ;
  assign n18427 = n69 & n31995 ;
  assign n18428 = n7041 & n32507 ;
  assign n18429 = n18427 | n18428 ;
  assign n18430 = n10941 | n18429 ;
  assign n18431 = n7068 & n13637 ;
  assign n18432 = n18430 | n18431 ;
  assign n18433 = n18426 | n18432 ;
  assign n33936 = ~n18433 ;
  assign n18435 = x8 & n33936 ;
  assign n18436 = n17919 | n18435 ;
  assign n13697 = n7068 & n13690 ;
  assign n10968 = n69 & n10940 ;
  assign n10984 = n7041 & n31995 ;
  assign n18438 = n10968 | n10984 ;
  assign n18439 = n7017 & n32503 ;
  assign n18440 = n18438 | n18439 ;
  assign n18441 = n13697 | n18440 ;
  assign n33937 = ~n18441 ;
  assign n18442 = x8 & n33937 ;
  assign n18443 = n30185 & n18441 ;
  assign n18444 = n18442 | n18443 ;
  assign n18445 = n18436 & n18444 ;
  assign n18446 = x11 & n17919 ;
  assign n33938 = ~n17923 ;
  assign n18447 = n33938 & n18446 ;
  assign n33939 = ~n18446 ;
  assign n18448 = n17923 & n33939 ;
  assign n18449 = n18447 | n18448 ;
  assign n18451 = n18445 | n18449 ;
  assign n13763 = n7068 & n13756 ;
  assign n10923 = n69 & n32503 ;
  assign n10969 = n7041 & n10940 ;
  assign n18452 = n10923 | n10969 ;
  assign n18453 = n7017 & n10892 ;
  assign n18454 = n18452 | n18453 ;
  assign n18455 = n13763 | n18454 ;
  assign n33940 = ~n18455 ;
  assign n18456 = x8 & n33940 ;
  assign n18457 = n30185 & n18455 ;
  assign n18458 = n18456 | n18457 ;
  assign n18450 = n18445 & n18449 ;
  assign n33941 = ~n18450 ;
  assign n18459 = n33941 & n18451 ;
  assign n33942 = ~n18458 ;
  assign n18460 = n33942 & n18459 ;
  assign n33943 = ~n18460 ;
  assign n18461 = n18451 & n33943 ;
  assign n33944 = ~n18461 ;
  assign n18463 = n18419 & n33944 ;
  assign n33945 = ~n18463 ;
  assign n18464 = n18418 & n33945 ;
  assign n18466 = n18408 & n18464 ;
  assign n18467 = n18406 | n18466 ;
  assign n33946 = ~n18467 ;
  assign n18468 = n18393 & n33946 ;
  assign n33947 = ~n18468 ;
  assign n18469 = n18391 & n33947 ;
  assign n33948 = ~n18469 ;
  assign n18471 = n18380 & n33948 ;
  assign n33949 = ~n18471 ;
  assign n18472 = n18379 & n33949 ;
  assign n33950 = ~n18472 ;
  assign n18474 = n18368 & n33950 ;
  assign n33951 = ~n18474 ;
  assign n18475 = n18367 & n33951 ;
  assign n33952 = ~n18475 ;
  assign n18477 = n18356 & n33952 ;
  assign n33953 = ~n18477 ;
  assign n18478 = n18354 & n33953 ;
  assign n33954 = ~n18478 ;
  assign n18480 = n18344 & n33954 ;
  assign n33955 = ~n18480 ;
  assign n18481 = n18342 & n33955 ;
  assign n18330 = n18322 & n18329 ;
  assign n33956 = ~n18330 ;
  assign n18482 = n33956 & n18331 ;
  assign n33957 = ~n18481 ;
  assign n18484 = n33957 & n18482 ;
  assign n33958 = ~n18484 ;
  assign n18485 = n18331 & n33958 ;
  assign n33959 = ~n18485 ;
  assign n18487 = n18320 & n33959 ;
  assign n33960 = ~n18487 ;
  assign n18488 = n18318 & n33960 ;
  assign n33961 = ~n18488 ;
  assign n18489 = n18307 & n33961 ;
  assign n33962 = ~n18489 ;
  assign n18490 = n18305 & n33962 ;
  assign n18491 = n18286 | n18293 ;
  assign n33963 = ~n18294 ;
  assign n18492 = n33963 & n18491 ;
  assign n18493 = n18490 & n18492 ;
  assign n18494 = n18294 | n18493 ;
  assign n33964 = ~n18494 ;
  assign n18496 = n18284 & n33964 ;
  assign n33965 = ~n18496 ;
  assign n18497 = n18282 & n33965 ;
  assign n33966 = ~n18497 ;
  assign n18499 = n18271 & n33966 ;
  assign n33967 = ~n18499 ;
  assign n18500 = n18269 & n33967 ;
  assign n33968 = ~n18500 ;
  assign n18501 = n18258 & n33968 ;
  assign n33969 = ~n18501 ;
  assign n18502 = n18256 & n33969 ;
  assign n33970 = ~n18502 ;
  assign n18504 = n18246 & n33970 ;
  assign n33971 = ~n18504 ;
  assign n18505 = n18245 & n33971 ;
  assign n18506 = n18226 | n18233 ;
  assign n33972 = ~n18234 ;
  assign n18507 = n33972 & n18506 ;
  assign n18509 = n18505 & n18507 ;
  assign n18510 = n18234 | n18509 ;
  assign n33973 = ~n18510 ;
  assign n18511 = n18224 & n33973 ;
  assign n33974 = ~n18511 ;
  assign n18512 = n18223 & n33974 ;
  assign n33975 = ~n18512 ;
  assign n18514 = n18212 & n33975 ;
  assign n33976 = ~n18514 ;
  assign n18515 = n18211 & n33976 ;
  assign n33977 = ~n18515 ;
  assign n18517 = n18200 & n33977 ;
  assign n33978 = ~n18517 ;
  assign n18518 = n18198 & n33978 ;
  assign n33979 = ~n18518 ;
  assign n18520 = n18188 & n33979 ;
  assign n33980 = ~n18520 ;
  assign n18521 = n18187 & n33980 ;
  assign n18523 = n18176 | n18521 ;
  assign n33981 = ~n18175 ;
  assign n18524 = n33981 & n18523 ;
  assign n18525 = n18164 | n18524 ;
  assign n33982 = ~n18162 ;
  assign n18526 = n33982 & n18525 ;
  assign n33983 = ~n18526 ;
  assign n18528 = n18151 & n33983 ;
  assign n33984 = ~n18528 ;
  assign n18529 = n18150 & n33984 ;
  assign n18531 = n18139 | n18529 ;
  assign n33985 = ~n18138 ;
  assign n18532 = n33985 & n18531 ;
  assign n18534 = n18127 | n18532 ;
  assign n33986 = ~n18126 ;
  assign n18535 = n33986 & n18534 ;
  assign n33987 = ~n18535 ;
  assign n18537 = n18115 & n33987 ;
  assign n33988 = ~n18537 ;
  assign n18538 = n18113 & n33988 ;
  assign n33989 = ~n18538 ;
  assign n18540 = n18102 & n33989 ;
  assign n33990 = ~n18540 ;
  assign n18541 = n18101 & n33990 ;
  assign n33991 = ~n18541 ;
  assign n18543 = n18090 & n33991 ;
  assign n33992 = ~n18543 ;
  assign n18544 = n18088 & n33992 ;
  assign n33993 = ~n18544 ;
  assign n18545 = n18077 & n33993 ;
  assign n33994 = ~n18545 ;
  assign n18546 = n18075 & n33994 ;
  assign n33995 = ~n18546 ;
  assign n18548 = n18064 & n33995 ;
  assign n33996 = ~n18548 ;
  assign n18549 = n18062 & n33996 ;
  assign n18551 = n18052 | n18549 ;
  assign n33997 = ~n18050 ;
  assign n18552 = n33997 & n18551 ;
  assign n18554 = n18040 | n18552 ;
  assign n18553 = n18040 & n18552 ;
  assign n33998 = ~n18553 ;
  assign n18555 = n33998 & n18554 ;
  assign n33999 = ~n18052 ;
  assign n18550 = n33999 & n18549 ;
  assign n34000 = ~n18549 ;
  assign n18556 = n18052 & n34000 ;
  assign n18557 = n18550 | n18556 ;
  assign n15531 = n8157 & n15526 ;
  assign n15163 = n8195 & n32876 ;
  assign n15254 = n740 & n32890 ;
  assign n18558 = n15163 | n15254 ;
  assign n18559 = n9052 & n15221 ;
  assign n18560 = n18558 | n18559 ;
  assign n18561 = n15531 | n18560 ;
  assign n18562 = x5 | n18561 ;
  assign n18563 = x5 & n18561 ;
  assign n34001 = ~n18563 ;
  assign n18564 = n18562 & n34001 ;
  assign n18565 = n734 & n18564 ;
  assign n18547 = n18064 & n18546 ;
  assign n18566 = n18064 | n18546 ;
  assign n34002 = ~n18547 ;
  assign n18567 = n34002 & n18566 ;
  assign n18568 = n734 | n18564 ;
  assign n34003 = ~n18565 ;
  assign n18569 = n34003 & n18568 ;
  assign n18570 = n18567 & n18569 ;
  assign n18571 = n18565 | n18570 ;
  assign n34004 = ~n18557 ;
  assign n18573 = n34004 & n18571 ;
  assign n34005 = ~n18571 ;
  assign n18572 = n18557 & n34005 ;
  assign n18574 = n18572 | n18573 ;
  assign n18575 = n18567 | n18569 ;
  assign n34006 = ~n18570 ;
  assign n18576 = n34006 & n18575 ;
  assign n34007 = ~n18077 ;
  assign n18577 = n34007 & n18544 ;
  assign n18578 = n18545 | n18577 ;
  assign n15270 = n8157 & n32889 ;
  assign n15062 = n8195 & n32856 ;
  assign n15162 = n740 & n32876 ;
  assign n18579 = n15062 | n15162 ;
  assign n18580 = n9052 & n32890 ;
  assign n18581 = n18579 | n18580 ;
  assign n18582 = n15270 | n18581 ;
  assign n18583 = x5 | n18582 ;
  assign n18584 = x5 & n18582 ;
  assign n34008 = ~n18584 ;
  assign n18585 = n18583 & n34008 ;
  assign n18587 = n18578 | n18585 ;
  assign n34009 = ~n18578 ;
  assign n18586 = n34009 & n18585 ;
  assign n34010 = ~n18585 ;
  assign n18588 = n18578 & n34010 ;
  assign n18589 = n18586 | n18588 ;
  assign n18542 = n18090 & n18541 ;
  assign n18590 = n18090 | n18541 ;
  assign n34011 = ~n18542 ;
  assign n18591 = n34011 & n18590 ;
  assign n15186 = n8157 & n32875 ;
  assign n15068 = n740 & n32856 ;
  assign n15091 = n8195 & n15081 ;
  assign n18592 = n15068 | n15091 ;
  assign n18593 = n9052 & n32876 ;
  assign n18594 = n18592 | n18593 ;
  assign n18595 = n15186 | n18594 ;
  assign n18596 = x5 | n18595 ;
  assign n18597 = x5 & n18595 ;
  assign n34012 = ~n18597 ;
  assign n18598 = n18596 & n34012 ;
  assign n18600 = n18591 | n18598 ;
  assign n18599 = n18591 & n18598 ;
  assign n34013 = ~n18599 ;
  assign n18601 = n34013 & n18600 ;
  assign n18539 = n18102 & n18538 ;
  assign n18602 = n18102 | n18538 ;
  assign n34014 = ~n18539 ;
  assign n18603 = n34014 & n18602 ;
  assign n15118 = n8157 & n15111 ;
  assign n14502 = n8195 & n32707 ;
  assign n15090 = n740 & n15081 ;
  assign n18604 = n14502 | n15090 ;
  assign n18605 = n9052 & n32856 ;
  assign n18606 = n18604 | n18605 ;
  assign n18607 = n15118 | n18606 ;
  assign n18608 = x5 | n18607 ;
  assign n18609 = x5 & n18607 ;
  assign n34015 = ~n18609 ;
  assign n18610 = n18608 & n34015 ;
  assign n18612 = n18603 | n18610 ;
  assign n18611 = n18603 & n18610 ;
  assign n34016 = ~n18611 ;
  assign n18613 = n34016 & n18612 ;
  assign n18536 = n18115 & n18535 ;
  assign n18614 = n18115 | n18535 ;
  assign n34017 = ~n18536 ;
  assign n18615 = n34017 & n18614 ;
  assign n15293 = n8157 & n15288 ;
  assign n14495 = n740 & n32707 ;
  assign n14515 = n8195 & n32706 ;
  assign n18616 = n14495 | n14515 ;
  assign n18617 = n9052 & n15081 ;
  assign n18618 = n18616 | n18617 ;
  assign n18619 = n15293 | n18618 ;
  assign n18620 = x5 | n18619 ;
  assign n18621 = x5 & n18619 ;
  assign n34018 = ~n18621 ;
  assign n18622 = n18620 & n34018 ;
  assign n18624 = n18615 | n18622 ;
  assign n18623 = n18615 & n18622 ;
  assign n34019 = ~n18623 ;
  assign n18625 = n34019 & n18624 ;
  assign n34020 = ~n18127 ;
  assign n18533 = n34020 & n18532 ;
  assign n34021 = ~n18532 ;
  assign n18626 = n18127 & n34021 ;
  assign n18627 = n18533 | n18626 ;
  assign n14575 = n8157 & n14570 ;
  assign n14517 = n740 & n32706 ;
  assign n14546 = n8195 & n14536 ;
  assign n18628 = n14517 | n14546 ;
  assign n18629 = n9052 & n32707 ;
  assign n18630 = n18628 | n18629 ;
  assign n18631 = n14575 | n18630 ;
  assign n18632 = x5 | n18631 ;
  assign n18633 = x5 & n18631 ;
  assign n34022 = ~n18633 ;
  assign n18634 = n18632 & n34022 ;
  assign n34023 = ~n18634 ;
  assign n18636 = n18627 & n34023 ;
  assign n34024 = ~n18627 ;
  assign n18635 = n34024 & n18634 ;
  assign n18637 = n18635 | n18636 ;
  assign n34025 = ~n18139 ;
  assign n18530 = n34025 & n18529 ;
  assign n34026 = ~n18529 ;
  assign n18638 = n18139 & n34026 ;
  assign n18639 = n18530 | n18638 ;
  assign n14683 = n8157 & n32735 ;
  assign n14115 = n8195 & n14101 ;
  assign n14538 = n740 & n14536 ;
  assign n18640 = n14115 | n14538 ;
  assign n18641 = n9052 & n32706 ;
  assign n18642 = n18640 | n18641 ;
  assign n18643 = n14683 | n18642 ;
  assign n18644 = x5 | n18643 ;
  assign n18645 = x5 & n18643 ;
  assign n34027 = ~n18645 ;
  assign n18646 = n18644 & n34027 ;
  assign n34028 = ~n18646 ;
  assign n18648 = n18639 & n34028 ;
  assign n34029 = ~n18639 ;
  assign n18647 = n34029 & n18646 ;
  assign n18649 = n18647 | n18648 ;
  assign n18527 = n18151 & n18526 ;
  assign n18650 = n18151 | n18526 ;
  assign n34030 = ~n18527 ;
  assign n18651 = n34030 & n18650 ;
  assign n14972 = n8157 & n14965 ;
  assign n14108 = n740 & n14101 ;
  assign n14133 = n8195 & n14124 ;
  assign n18652 = n14108 | n14133 ;
  assign n18653 = n9052 & n14536 ;
  assign n18654 = n18652 | n18653 ;
  assign n18655 = n14972 | n18654 ;
  assign n18656 = x5 | n18655 ;
  assign n18657 = x5 & n18655 ;
  assign n34031 = ~n18657 ;
  assign n18658 = n18656 & n34031 ;
  assign n18660 = n18651 | n18658 ;
  assign n18659 = n18651 & n18658 ;
  assign n34032 = ~n18659 ;
  assign n18661 = n34032 & n18660 ;
  assign n18662 = n18164 & n18524 ;
  assign n34033 = ~n18662 ;
  assign n18663 = n18525 & n34033 ;
  assign n14187 = n8157 & n14183 ;
  assign n14134 = n740 & n14124 ;
  assign n14162 = n8195 & n14147 ;
  assign n18664 = n14134 | n14162 ;
  assign n18665 = n9052 & n14196 ;
  assign n18666 = n18664 | n18665 ;
  assign n18667 = n14187 | n18666 ;
  assign n18668 = x5 | n18667 ;
  assign n18669 = x5 & n18667 ;
  assign n34034 = ~n18669 ;
  assign n18670 = n18668 & n34034 ;
  assign n34035 = ~n18670 ;
  assign n18672 = n18663 & n34035 ;
  assign n18671 = n18663 & n18670 ;
  assign n18673 = n18663 | n18670 ;
  assign n34036 = ~n18671 ;
  assign n18674 = n34036 & n18673 ;
  assign n34037 = ~n18176 ;
  assign n18522 = n34037 & n18521 ;
  assign n34038 = ~n18521 ;
  assign n18675 = n18176 & n34038 ;
  assign n18676 = n18522 | n18675 ;
  assign n14292 = n8157 & n14283 ;
  assign n13046 = n8195 & n13027 ;
  assign n14163 = n740 & n14147 ;
  assign n18677 = n13046 | n14163 ;
  assign n18678 = n9052 & n14295 ;
  assign n18679 = n18677 | n18678 ;
  assign n18680 = n14292 | n18679 ;
  assign n18681 = x5 | n18680 ;
  assign n18682 = x5 & n18680 ;
  assign n34039 = ~n18682 ;
  assign n18683 = n18681 & n34039 ;
  assign n34040 = ~n18683 ;
  assign n18685 = n18676 & n34040 ;
  assign n18684 = n18676 & n18683 ;
  assign n18686 = n18676 | n18683 ;
  assign n34041 = ~n18684 ;
  assign n18687 = n34041 & n18686 ;
  assign n18519 = n18188 & n18518 ;
  assign n18688 = n18188 | n18518 ;
  assign n34042 = ~n18519 ;
  assign n18689 = n34042 & n18688 ;
  assign n14663 = n8157 & n14655 ;
  assign n13036 = n740 & n13027 ;
  assign n13061 = n8195 & n32456 ;
  assign n18690 = n13036 | n13061 ;
  assign n18691 = n9052 & n14147 ;
  assign n18692 = n18690 | n18691 ;
  assign n18693 = n14663 | n18692 ;
  assign n18694 = x5 | n18693 ;
  assign n18695 = x5 & n18693 ;
  assign n34043 = ~n18695 ;
  assign n18696 = n18694 & n34043 ;
  assign n18698 = n18689 | n18696 ;
  assign n18516 = n18200 & n18515 ;
  assign n18699 = n18200 | n18515 ;
  assign n34044 = ~n18516 ;
  assign n18700 = n34044 & n18699 ;
  assign n13123 = n8157 & n32455 ;
  assign n13069 = n740 & n32456 ;
  assign n13093 = n8195 & n13077 ;
  assign n18701 = n13069 | n13093 ;
  assign n18702 = n9052 & n13027 ;
  assign n18703 = n18701 | n18702 ;
  assign n18704 = n13123 | n18703 ;
  assign n18705 = x5 | n18704 ;
  assign n18706 = x5 & n18704 ;
  assign n34045 = ~n18706 ;
  assign n18707 = n18705 & n34045 ;
  assign n18709 = n18700 | n18707 ;
  assign n18708 = n18700 & n18707 ;
  assign n18513 = n18212 & n18512 ;
  assign n18710 = n18212 | n18512 ;
  assign n34046 = ~n18513 ;
  assign n18711 = n34046 & n18710 ;
  assign n14264 = n8157 & n32641 ;
  assign n12563 = n740 & n32354 ;
  assign n12587 = n8195 & n12570 ;
  assign n18712 = n12563 | n12587 ;
  assign n18713 = n9052 & n13077 ;
  assign n18714 = n18712 | n18713 ;
  assign n18715 = n14264 | n18714 ;
  assign n18716 = x5 | n18715 ;
  assign n18717 = x5 & n18715 ;
  assign n34047 = ~n18717 ;
  assign n18718 = n18716 & n34047 ;
  assign n34048 = ~n18505 ;
  assign n18508 = n34048 & n18507 ;
  assign n34049 = ~n18507 ;
  assign n18719 = n18505 & n34049 ;
  assign n18720 = n18508 | n18719 ;
  assign n12638 = n8157 & n32356 ;
  assign n12591 = n740 & n12570 ;
  assign n12614 = n8195 & n12595 ;
  assign n18721 = n12591 | n12614 ;
  assign n18722 = n9052 & n32354 ;
  assign n18723 = n18721 | n18722 ;
  assign n18724 = n12638 | n18723 ;
  assign n18725 = x5 | n18724 ;
  assign n18726 = x5 & n18724 ;
  assign n34050 = ~n18726 ;
  assign n18727 = n18725 & n34050 ;
  assign n18729 = n18720 | n18727 ;
  assign n34051 = ~n18720 ;
  assign n18728 = n34051 & n18727 ;
  assign n34052 = ~n18727 ;
  assign n18730 = n18720 & n34052 ;
  assign n18731 = n18728 | n18730 ;
  assign n34053 = ~n18246 ;
  assign n18503 = n34053 & n18502 ;
  assign n18732 = n18503 | n18504 ;
  assign n12688 = n8157 & n12681 ;
  assign n12148 = n8195 & n32253 ;
  assign n12607 = n740 & n12595 ;
  assign n18733 = n12148 | n12607 ;
  assign n18734 = n9052 & n12570 ;
  assign n18735 = n18733 | n18734 ;
  assign n18736 = n12688 | n18735 ;
  assign n18737 = x5 | n18736 ;
  assign n18738 = x5 & n18736 ;
  assign n34054 = ~n18738 ;
  assign n18739 = n18737 & n34054 ;
  assign n18741 = n18732 | n18739 ;
  assign n34055 = ~n18732 ;
  assign n18740 = n34055 & n18739 ;
  assign n34056 = ~n18739 ;
  assign n18742 = n18732 & n34056 ;
  assign n18743 = n18740 | n18742 ;
  assign n34057 = ~n18258 ;
  assign n18744 = n34057 & n18500 ;
  assign n18745 = n18501 | n18744 ;
  assign n13824 = n8157 & n32550 ;
  assign n12156 = n740 & n32253 ;
  assign n12170 = n8195 & n12161 ;
  assign n18746 = n12156 | n12170 ;
  assign n18747 = n9052 & n12595 ;
  assign n18748 = n18746 | n18747 ;
  assign n18749 = n13824 | n18748 ;
  assign n18750 = x5 | n18749 ;
  assign n18751 = x5 & n18749 ;
  assign n34058 = ~n18751 ;
  assign n18752 = n18750 & n34058 ;
  assign n18754 = n18745 | n18752 ;
  assign n34059 = ~n18271 ;
  assign n18498 = n34059 & n18497 ;
  assign n18755 = n18498 | n18499 ;
  assign n12663 = n8157 & n32362 ;
  assign n11450 = n8195 & n11430 ;
  assign n11859 = n740 & n32176 ;
  assign n18756 = n11450 | n11859 ;
  assign n18757 = n9052 & n12161 ;
  assign n18758 = n18756 | n18757 ;
  assign n18759 = n12663 | n18758 ;
  assign n34060 = ~n18759 ;
  assign n18760 = x5 & n34060 ;
  assign n18761 = n30053 & n18759 ;
  assign n18762 = n18760 | n18761 ;
  assign n18763 = n18490 | n18492 ;
  assign n34061 = ~n18493 ;
  assign n18764 = n34061 & n18763 ;
  assign n11874 = n8157 & n32178 ;
  assign n11451 = n740 & n11430 ;
  assign n11496 = n8195 & n11476 ;
  assign n18765 = n11451 | n11496 ;
  assign n18766 = n9052 & n32176 ;
  assign n18767 = n18765 | n18766 ;
  assign n18768 = n11874 | n18767 ;
  assign n18769 = x5 | n18768 ;
  assign n18770 = x5 & n18768 ;
  assign n34062 = ~n18770 ;
  assign n18771 = n18769 & n34062 ;
  assign n18772 = n18764 & n18771 ;
  assign n18773 = n18764 | n18771 ;
  assign n34063 = ~n18772 ;
  assign n18774 = n34063 & n18773 ;
  assign n34064 = ~n18307 ;
  assign n18775 = n34064 & n18488 ;
  assign n18776 = n18489 | n18775 ;
  assign n11469 = n8157 & n11463 ;
  assign n10677 = n8195 & n10656 ;
  assign n11488 = n740 & n11476 ;
  assign n18777 = n10677 | n11488 ;
  assign n18778 = n9052 & n11430 ;
  assign n18779 = n18777 | n18778 ;
  assign n18780 = n11469 | n18779 ;
  assign n18781 = x5 | n18780 ;
  assign n18782 = x5 & n18780 ;
  assign n34065 = ~n18782 ;
  assign n18783 = n18781 & n34065 ;
  assign n18785 = n18776 | n18783 ;
  assign n34066 = ~n18776 ;
  assign n18784 = n34066 & n18783 ;
  assign n34067 = ~n18783 ;
  assign n18786 = n18776 & n34067 ;
  assign n18787 = n18784 | n18786 ;
  assign n18486 = n18320 & n18485 ;
  assign n18788 = n18320 | n18485 ;
  assign n34068 = ~n18486 ;
  assign n18789 = n34068 & n18788 ;
  assign n11519 = n8157 & n11511 ;
  assign n10669 = n740 & n10656 ;
  assign n11043 = n8195 & n10679 ;
  assign n18790 = n10669 | n11043 ;
  assign n18791 = n9052 & n11452 ;
  assign n18792 = n18790 | n18791 ;
  assign n18793 = n11519 | n18792 ;
  assign n18794 = x5 | n18793 ;
  assign n18795 = x5 & n18793 ;
  assign n34069 = ~n18795 ;
  assign n18796 = n18794 & n34069 ;
  assign n18797 = n18789 & n18796 ;
  assign n18798 = n18789 | n18796 ;
  assign n34070 = ~n18797 ;
  assign n18799 = n34070 & n18798 ;
  assign n18483 = n18481 & n18482 ;
  assign n18800 = n18481 | n18482 ;
  assign n34071 = ~n18483 ;
  assign n18801 = n34071 & n18800 ;
  assign n11040 = n8157 & n11030 ;
  assign n10694 = n8195 & n10681 ;
  assign n11053 = n740 & n10679 ;
  assign n18802 = n10694 | n11053 ;
  assign n18803 = n9052 & n10656 ;
  assign n18804 = n18802 | n18803 ;
  assign n18805 = n11040 | n18804 ;
  assign n18806 = x5 | n18805 ;
  assign n18807 = x5 & n18805 ;
  assign n34072 = ~n18807 ;
  assign n18808 = n18806 & n34072 ;
  assign n18810 = n18801 | n18808 ;
  assign n18479 = n18344 & n18478 ;
  assign n18811 = n18344 | n18478 ;
  assign n34073 = ~n18479 ;
  assign n18812 = n34073 & n18811 ;
  assign n11546 = n8157 & n11536 ;
  assign n10701 = n740 & n10681 ;
  assign n10711 = n8195 & n10703 ;
  assign n18813 = n10701 | n10711 ;
  assign n18814 = n9052 & n10679 ;
  assign n18815 = n18813 | n18814 ;
  assign n18816 = n11546 | n18815 ;
  assign n18817 = x5 | n18816 ;
  assign n18818 = x5 & n18816 ;
  assign n34074 = ~n18818 ;
  assign n18819 = n18817 & n34074 ;
  assign n18821 = n18812 | n18819 ;
  assign n18820 = n18812 & n18819 ;
  assign n34075 = ~n18820 ;
  assign n18822 = n34075 & n18821 ;
  assign n13168 = n8157 & n13157 ;
  assign n10707 = n740 & n10703 ;
  assign n10742 = n8195 & n10727 ;
  assign n18823 = n10707 | n10742 ;
  assign n18824 = n9052 & n10681 ;
  assign n18825 = n18823 | n18824 ;
  assign n18826 = n13168 | n18825 ;
  assign n18827 = x5 | n18826 ;
  assign n18828 = x5 & n18826 ;
  assign n34076 = ~n18828 ;
  assign n18829 = n18827 & n34076 ;
  assign n18473 = n18368 & n18472 ;
  assign n18830 = n18368 | n18472 ;
  assign n34077 = ~n18473 ;
  assign n18831 = n34077 & n18830 ;
  assign n13192 = n8157 & n13182 ;
  assign n10747 = n740 & n10727 ;
  assign n10770 = n8195 & n31999 ;
  assign n18832 = n10747 | n10770 ;
  assign n18833 = n9052 & n13151 ;
  assign n18834 = n18832 | n18833 ;
  assign n18835 = n13192 | n18834 ;
  assign n18836 = x5 | n18835 ;
  assign n18837 = x5 & n18835 ;
  assign n34078 = ~n18837 ;
  assign n18838 = n18836 & n34078 ;
  assign n18840 = n18831 | n18838 ;
  assign n34079 = ~n18831 ;
  assign n18839 = n34079 & n18838 ;
  assign n34080 = ~n18838 ;
  assign n18841 = n18831 & n34080 ;
  assign n18842 = n18839 | n18841 ;
  assign n18470 = n18380 & n18469 ;
  assign n18843 = n18380 | n18469 ;
  assign n34081 = ~n18470 ;
  assign n18844 = n34081 & n18843 ;
  assign n11697 = n8157 & n32125 ;
  assign n10762 = n740 & n31999 ;
  assign n10775 = n8195 & n10773 ;
  assign n18845 = n10762 | n10775 ;
  assign n18846 = n9052 & n10727 ;
  assign n18847 = n18845 | n18846 ;
  assign n18848 = n11697 | n18847 ;
  assign n18849 = x5 | n18848 ;
  assign n18850 = x5 & n18848 ;
  assign n34082 = ~n18850 ;
  assign n18851 = n18849 & n34082 ;
  assign n18852 = n18844 & n18851 ;
  assign n18853 = n18844 | n18851 ;
  assign n34083 = ~n18852 ;
  assign n18854 = n34083 & n18853 ;
  assign n13233 = n8157 & n32477 ;
  assign n10793 = n740 & n10773 ;
  assign n10815 = n8195 & n31998 ;
  assign n18855 = n10793 | n10815 ;
  assign n18856 = n9052 & n32478 ;
  assign n18857 = n18855 | n18856 ;
  assign n18858 = n13233 | n18857 ;
  assign n34084 = ~n18858 ;
  assign n18859 = x5 & n34084 ;
  assign n18860 = n30053 & n18858 ;
  assign n18861 = n18859 | n18860 ;
  assign n34085 = ~n18393 ;
  assign n18862 = n34085 & n18467 ;
  assign n18863 = n18468 | n18862 ;
  assign n18864 = n18861 | n18863 ;
  assign n18865 = n18861 & n18863 ;
  assign n34086 = ~n18865 ;
  assign n18866 = n18864 & n34086 ;
  assign n34087 = ~n18408 ;
  assign n18465 = n34087 & n18464 ;
  assign n34088 = ~n18464 ;
  assign n18867 = n18408 & n34088 ;
  assign n18868 = n18465 | n18867 ;
  assign n13290 = n8157 & n32482 ;
  assign n10816 = n740 & n31998 ;
  assign n10838 = n8195 & n10818 ;
  assign n18869 = n10816 | n10838 ;
  assign n18870 = n9052 & n13292 ;
  assign n18871 = n18869 | n18870 ;
  assign n18872 = n13290 | n18871 ;
  assign n18873 = x5 | n18872 ;
  assign n18874 = x5 & n18872 ;
  assign n34089 = ~n18874 ;
  assign n18875 = n18873 & n34089 ;
  assign n18877 = n18868 | n18875 ;
  assign n18876 = n18868 & n18875 ;
  assign n34090 = ~n18876 ;
  assign n18878 = n34090 & n18877 ;
  assign n13328 = n8157 & n32488 ;
  assign n10839 = n740 & n10818 ;
  assign n10851 = n8195 & n10841 ;
  assign n18879 = n10839 | n10851 ;
  assign n18880 = n9052 & n31998 ;
  assign n18881 = n18879 | n18880 ;
  assign n18882 = n13328 | n18881 ;
  assign n34091 = ~n18882 ;
  assign n18883 = x5 & n34091 ;
  assign n18884 = n30053 & n18882 ;
  assign n18885 = n18883 | n18884 ;
  assign n13393 = n8157 & n13382 ;
  assign n10857 = n740 & n10841 ;
  assign n10867 = n8195 & n10865 ;
  assign n18886 = n10857 | n10867 ;
  assign n18887 = n9052 & n10818 ;
  assign n18888 = n18886 | n18887 ;
  assign n18889 = n13393 | n18888 ;
  assign n18890 = x5 | n18889 ;
  assign n18891 = x5 & n18889 ;
  assign n34092 = ~n18891 ;
  assign n18892 = n18890 & n34092 ;
  assign n34093 = ~n18459 ;
  assign n18893 = n18458 & n34093 ;
  assign n18894 = n18460 | n18893 ;
  assign n18896 = n18892 & n18894 ;
  assign n34094 = ~n18894 ;
  assign n18895 = n18892 & n34094 ;
  assign n34095 = ~n18892 ;
  assign n18897 = n34095 & n18894 ;
  assign n18898 = n18895 | n18897 ;
  assign n13465 = n8157 & n13456 ;
  assign n10879 = n740 & n10865 ;
  assign n10900 = n8195 & n10892 ;
  assign n18899 = n10879 | n10900 ;
  assign n18900 = n9052 & n10841 ;
  assign n18901 = n18899 | n18900 ;
  assign n18902 = n13465 | n18901 ;
  assign n34096 = ~n18902 ;
  assign n18903 = x5 & n34096 ;
  assign n18904 = n30053 & n18902 ;
  assign n18905 = n18903 | n18904 ;
  assign n34097 = ~n18435 ;
  assign n18437 = n10992 & n34097 ;
  assign n18434 = x8 & n18433 ;
  assign n34098 = ~x9 ;
  assign n18907 = n34098 & n18434 ;
  assign n34099 = ~n18434 ;
  assign n18906 = x9 & n34099 ;
  assign n18908 = n10992 | n18906 ;
  assign n18909 = n18907 | n18908 ;
  assign n34100 = ~n18437 ;
  assign n18910 = n34100 & n18909 ;
  assign n34101 = ~n18444 ;
  assign n18911 = n34101 & n18910 ;
  assign n34102 = ~n18910 ;
  assign n18912 = n18444 & n34102 ;
  assign n18913 = n18911 | n18912 ;
  assign n18915 = n18905 | n18913 ;
  assign n34103 = ~n18905 ;
  assign n18914 = n34103 & n18913 ;
  assign n34104 = ~n18913 ;
  assign n18916 = n18905 & n34104 ;
  assign n18917 = n18914 | n18916 ;
  assign n18918 = x8 & n18426 ;
  assign n18919 = n18432 & n18918 ;
  assign n18920 = n18432 | n18918 ;
  assign n34105 = ~n18919 ;
  assign n18921 = n34105 & n18920 ;
  assign n13531 = n8157 & n32502 ;
  assign n10908 = n740 & n10892 ;
  assign n10937 = n8195 & n32503 ;
  assign n18922 = n10908 | n10937 ;
  assign n18923 = n9052 & n10865 ;
  assign n18924 = n18922 | n18923 ;
  assign n18925 = n13531 | n18924 ;
  assign n18926 = x5 | n18925 ;
  assign n18927 = x5 & n18925 ;
  assign n34106 = ~n18927 ;
  assign n18928 = n18926 & n34106 ;
  assign n18930 = n18921 | n18928 ;
  assign n18929 = n18921 & n18928 ;
  assign n34107 = ~n18929 ;
  assign n18931 = n34107 & n18930 ;
  assign n18932 = n9969 & n32507 ;
  assign n14868 = n8157 & n14859 ;
  assign n18933 = n9052 & n31995 ;
  assign n18934 = n740 & n32507 ;
  assign n18935 = n18933 | n18934 ;
  assign n18936 = n14868 | n18935 ;
  assign n18937 = n18932 | n18936 ;
  assign n10946 = n9052 & n10940 ;
  assign n18938 = n740 & n31995 ;
  assign n18939 = n8195 & n32507 ;
  assign n18940 = n18938 | n18939 ;
  assign n18941 = n10946 | n18940 ;
  assign n18942 = n8157 & n13637 ;
  assign n18943 = n18941 | n18942 ;
  assign n18944 = n18937 | n18943 ;
  assign n34108 = ~n18944 ;
  assign n18946 = x5 & n34108 ;
  assign n18947 = n18420 | n18946 ;
  assign n13701 = n8157 & n13690 ;
  assign n10970 = n740 & n10940 ;
  assign n10985 = n8195 & n31995 ;
  assign n18949 = n10970 | n10985 ;
  assign n18950 = n9052 & n32503 ;
  assign n18951 = n18949 | n18950 ;
  assign n18952 = n13701 | n18951 ;
  assign n34109 = ~n18952 ;
  assign n18953 = x5 & n34109 ;
  assign n18954 = n30053 & n18952 ;
  assign n18955 = n18953 | n18954 ;
  assign n18956 = n18947 & n18955 ;
  assign n18957 = n18421 & n18425 ;
  assign n34110 = ~n18957 ;
  assign n18958 = n18426 & n34110 ;
  assign n18960 = n18956 | n18958 ;
  assign n13766 = n8157 & n13756 ;
  assign n10931 = n740 & n32503 ;
  assign n10971 = n8195 & n10940 ;
  assign n18961 = n10931 | n10971 ;
  assign n18962 = n9052 & n10892 ;
  assign n18963 = n18961 | n18962 ;
  assign n18964 = n13766 | n18963 ;
  assign n18965 = x5 | n18964 ;
  assign n18966 = x5 & n18964 ;
  assign n34111 = ~n18966 ;
  assign n18967 = n18965 & n34111 ;
  assign n18959 = n18956 & n18958 ;
  assign n34112 = ~n18959 ;
  assign n18968 = n34112 & n18960 ;
  assign n34113 = ~n18967 ;
  assign n18969 = n34113 & n18968 ;
  assign n34114 = ~n18969 ;
  assign n18971 = n18960 & n34114 ;
  assign n34115 = ~n18971 ;
  assign n18973 = n18931 & n34115 ;
  assign n34116 = ~n18973 ;
  assign n18974 = n18930 & n34116 ;
  assign n34117 = ~n18974 ;
  assign n18976 = n18917 & n34117 ;
  assign n34118 = ~n18976 ;
  assign n18977 = n18915 & n34118 ;
  assign n18978 = n18898 & n18977 ;
  assign n18979 = n18896 | n18978 ;
  assign n18981 = n18885 & n18979 ;
  assign n18462 = n18419 & n18461 ;
  assign n18982 = n18419 | n18461 ;
  assign n34119 = ~n18462 ;
  assign n18983 = n34119 & n18982 ;
  assign n18980 = n18885 | n18979 ;
  assign n34120 = ~n18981 ;
  assign n18984 = n18980 & n34120 ;
  assign n18985 = n18983 & n18984 ;
  assign n18986 = n18981 | n18985 ;
  assign n34121 = ~n18986 ;
  assign n18988 = n18878 & n34121 ;
  assign n34122 = ~n18988 ;
  assign n18989 = n18877 & n34122 ;
  assign n34123 = ~n18989 ;
  assign n18991 = n18866 & n34123 ;
  assign n34124 = ~n18991 ;
  assign n18992 = n18864 & n34124 ;
  assign n18993 = n18854 & n18992 ;
  assign n18994 = n18852 | n18993 ;
  assign n34125 = ~n18994 ;
  assign n18995 = n18842 & n34125 ;
  assign n34126 = ~n18995 ;
  assign n18996 = n18840 & n34126 ;
  assign n18998 = n18829 | n18996 ;
  assign n18476 = n18356 & n18475 ;
  assign n18999 = n18356 | n18475 ;
  assign n34127 = ~n18476 ;
  assign n19000 = n34127 & n18999 ;
  assign n18997 = n18829 & n18996 ;
  assign n34128 = ~n18997 ;
  assign n19001 = n34128 & n18998 ;
  assign n34129 = ~n19000 ;
  assign n19002 = n34129 & n19001 ;
  assign n34130 = ~n19002 ;
  assign n19003 = n18998 & n34130 ;
  assign n34131 = ~n19003 ;
  assign n19005 = n18822 & n34131 ;
  assign n34132 = ~n19005 ;
  assign n19006 = n18821 & n34132 ;
  assign n18809 = n18801 & n18808 ;
  assign n34133 = ~n18809 ;
  assign n19007 = n34133 & n18810 ;
  assign n34134 = ~n19006 ;
  assign n19008 = n34134 & n19007 ;
  assign n34135 = ~n19008 ;
  assign n19009 = n18810 & n34135 ;
  assign n19010 = n18799 & n19009 ;
  assign n19011 = n18797 | n19010 ;
  assign n34136 = ~n19011 ;
  assign n19012 = n18787 & n34136 ;
  assign n34137 = ~n19012 ;
  assign n19013 = n18785 & n34137 ;
  assign n19014 = n18774 & n19013 ;
  assign n19015 = n18772 | n19014 ;
  assign n19017 = n18762 & n19015 ;
  assign n18495 = n18284 | n18494 ;
  assign n19018 = n18284 & n18494 ;
  assign n34138 = ~n19018 ;
  assign n19019 = n18495 & n34138 ;
  assign n19016 = n18762 | n19015 ;
  assign n34139 = ~n19017 ;
  assign n19020 = n19016 & n34139 ;
  assign n19021 = n19019 & n19020 ;
  assign n19022 = n19017 | n19021 ;
  assign n19023 = n18755 | n19022 ;
  assign n12202 = n8157 & n32255 ;
  assign n11860 = n8195 & n32176 ;
  assign n12181 = n740 & n12161 ;
  assign n19024 = n11860 | n12181 ;
  assign n19025 = n9052 & n32253 ;
  assign n19026 = n19024 | n19025 ;
  assign n19027 = n12202 | n19026 ;
  assign n19028 = x5 | n19027 ;
  assign n19029 = x5 & n19027 ;
  assign n34140 = ~n19029 ;
  assign n19030 = n19028 & n34140 ;
  assign n19031 = n18755 & n19022 ;
  assign n34141 = ~n19031 ;
  assign n19032 = n19023 & n34141 ;
  assign n34142 = ~n19030 ;
  assign n19034 = n34142 & n19032 ;
  assign n34143 = ~n19034 ;
  assign n19035 = n19023 & n34143 ;
  assign n18753 = n18745 & n18752 ;
  assign n34144 = ~n18753 ;
  assign n19036 = n34144 & n18754 ;
  assign n34145 = ~n19035 ;
  assign n19037 = n34145 & n19036 ;
  assign n34146 = ~n19037 ;
  assign n19038 = n18754 & n34146 ;
  assign n34147 = ~n19038 ;
  assign n19040 = n18743 & n34147 ;
  assign n34148 = ~n19040 ;
  assign n19041 = n18741 & n34148 ;
  assign n34149 = ~n19041 ;
  assign n19042 = n18731 & n34149 ;
  assign n34150 = ~n19042 ;
  assign n19043 = n18729 & n34150 ;
  assign n19045 = n18718 | n19043 ;
  assign n34151 = ~n18224 ;
  assign n19046 = n34151 & n18510 ;
  assign n19047 = n18511 | n19046 ;
  assign n19044 = n18718 & n19043 ;
  assign n34152 = ~n19044 ;
  assign n19048 = n34152 & n19045 ;
  assign n34153 = ~n19047 ;
  assign n19049 = n34153 & n19048 ;
  assign n34154 = ~n19049 ;
  assign n19050 = n19045 & n34154 ;
  assign n19052 = n18711 | n19050 ;
  assign n13857 = n8157 & n32557 ;
  assign n12551 = n8195 & n32354 ;
  assign n13080 = n740 & n13077 ;
  assign n19053 = n12551 | n13080 ;
  assign n19054 = n9052 & n32456 ;
  assign n19055 = n19053 | n19054 ;
  assign n19056 = n13857 | n19055 ;
  assign n19057 = x5 | n19056 ;
  assign n19058 = x5 & n19056 ;
  assign n34155 = ~n19058 ;
  assign n19059 = n19057 & n34155 ;
  assign n19051 = n18711 & n19050 ;
  assign n34156 = ~n19051 ;
  assign n19060 = n34156 & n19052 ;
  assign n34157 = ~n19059 ;
  assign n19062 = n34157 & n19060 ;
  assign n34158 = ~n19062 ;
  assign n19063 = n19052 & n34158 ;
  assign n19064 = n18708 | n19063 ;
  assign n19065 = n18709 & n19064 ;
  assign n18697 = n18689 & n18696 ;
  assign n34159 = ~n18697 ;
  assign n19066 = n34159 & n18698 ;
  assign n34160 = ~n19065 ;
  assign n19068 = n34160 & n19066 ;
  assign n34161 = ~n19068 ;
  assign n19069 = n18698 & n34161 ;
  assign n19071 = n18687 | n19069 ;
  assign n34162 = ~n18685 ;
  assign n19072 = n34162 & n19071 ;
  assign n19073 = n18674 | n19072 ;
  assign n34163 = ~n18672 ;
  assign n19074 = n34163 & n19073 ;
  assign n34164 = ~n19074 ;
  assign n19076 = n18661 & n34164 ;
  assign n34165 = ~n19076 ;
  assign n19077 = n18660 & n34165 ;
  assign n19079 = n18649 | n19077 ;
  assign n34166 = ~n18648 ;
  assign n19080 = n34166 & n19079 ;
  assign n19082 = n18637 | n19080 ;
  assign n34167 = ~n18636 ;
  assign n19083 = n34167 & n19082 ;
  assign n34168 = ~n19083 ;
  assign n19084 = n18625 & n34168 ;
  assign n34169 = ~n19084 ;
  assign n19085 = n18624 & n34169 ;
  assign n34170 = ~n19085 ;
  assign n19087 = n18613 & n34170 ;
  assign n34171 = ~n19087 ;
  assign n19088 = n18612 & n34171 ;
  assign n34172 = ~n19088 ;
  assign n19090 = n18601 & n34172 ;
  assign n34173 = ~n19090 ;
  assign n19091 = n18600 & n34173 ;
  assign n34174 = ~n19091 ;
  assign n19093 = n18589 & n34174 ;
  assign n34175 = ~n19093 ;
  assign n19094 = n18587 & n34175 ;
  assign n19096 = n18576 | n19094 ;
  assign n19097 = n18576 & n19094 ;
  assign n19092 = n18589 | n19091 ;
  assign n19098 = n18589 & n19091 ;
  assign n34176 = ~n19098 ;
  assign n19099 = n19092 & n34176 ;
  assign n19086 = n18613 & n19085 ;
  assign n19100 = n18613 | n19085 ;
  assign n34177 = ~n19086 ;
  assign n19101 = n34177 & n19100 ;
  assign n15229 = n10105 & n15221 ;
  assign n15255 = n10126 & n32890 ;
  assign n19102 = n15229 | n15255 ;
  assign n19103 = n9562 & n15526 ;
  assign n19104 = n19102 | n19103 ;
  assign n19105 = n30049 & n19104 ;
  assign n15164 = n733 | n15158 ;
  assign n19106 = x2 & n15164 ;
  assign n34178 = ~n19104 ;
  assign n19107 = n34178 & n19106 ;
  assign n19108 = n19105 | n19107 ;
  assign n19110 = n19101 | n19108 ;
  assign n34179 = ~n19101 ;
  assign n19109 = n34179 & n19108 ;
  assign n34180 = ~n19108 ;
  assign n19111 = n19101 & n34180 ;
  assign n19112 = n19109 | n19111 ;
  assign n15272 = n9562 & n32889 ;
  assign n15070 = n9552 & n32856 ;
  assign n15160 = n10126 & n32876 ;
  assign n19113 = n15070 | n15160 ;
  assign n19114 = n10105 & n32890 ;
  assign n19115 = n19113 | n19114 ;
  assign n19116 = n15272 | n19115 ;
  assign n34181 = ~n19116 ;
  assign n19117 = x2 & n34181 ;
  assign n19118 = n30049 & n19116 ;
  assign n19119 = n19117 | n19118 ;
  assign n19075 = n18661 & n19074 ;
  assign n19120 = n18661 | n19074 ;
  assign n34182 = ~n19075 ;
  assign n19121 = n34182 & n19120 ;
  assign n14516 = n9552 & n32706 ;
  assign n15295 = n9562 & n15288 ;
  assign n19122 = n10126 & n32707 ;
  assign n19123 = n10105 & n15081 ;
  assign n19124 = n19122 | n19123 ;
  assign n19125 = n15295 | n19124 ;
  assign n34183 = ~n19125 ;
  assign n19126 = x2 & n34183 ;
  assign n19127 = n30049 & n19125 ;
  assign n19128 = n19126 | n19127 ;
  assign n34184 = ~n14516 ;
  assign n19129 = n34184 & n19128 ;
  assign n19131 = n19121 | n19129 ;
  assign n19130 = n19121 & n19129 ;
  assign n34185 = ~n19130 ;
  assign n19132 = n34185 & n19131 ;
  assign n19133 = n18674 & n19072 ;
  assign n34186 = ~n19133 ;
  assign n19134 = n19073 & n34186 ;
  assign n14537 = n9552 & n14536 ;
  assign n14578 = n9562 & n14570 ;
  assign n19135 = n10105 & n32707 ;
  assign n19136 = n10126 & n32706 ;
  assign n19137 = n19135 | n19136 ;
  assign n19138 = n14578 | n19137 ;
  assign n34187 = ~n19138 ;
  assign n19139 = x2 & n34187 ;
  assign n19140 = n30049 & n19138 ;
  assign n19141 = n19139 | n19140 ;
  assign n34188 = ~n14537 ;
  assign n19142 = n34188 & n19141 ;
  assign n34189 = ~n19134 ;
  assign n19143 = n34189 & n19142 ;
  assign n34190 = ~n19142 ;
  assign n19144 = n19134 & n34190 ;
  assign n19145 = n19143 | n19144 ;
  assign n19067 = n19065 & n19066 ;
  assign n19146 = n19065 | n19066 ;
  assign n34191 = ~n19067 ;
  assign n19147 = n34191 & n19146 ;
  assign n19061 = n19059 & n19060 ;
  assign n19148 = n19059 | n19060 ;
  assign n34192 = ~n19061 ;
  assign n19149 = n34192 & n19148 ;
  assign n14288 = n9562 & n14283 ;
  assign n13047 = n9552 & n13027 ;
  assign n14164 = n10126 & n14147 ;
  assign n19150 = n13047 | n14164 ;
  assign n19151 = n10105 & n14295 ;
  assign n19152 = n19150 | n19151 ;
  assign n19153 = n14288 | n19152 ;
  assign n19154 = x2 | n19153 ;
  assign n19156 = x2 & n19153 ;
  assign n34193 = ~n19156 ;
  assign n19157 = n19154 & n34193 ;
  assign n19158 = n19149 | n19157 ;
  assign n34194 = ~n19153 ;
  assign n19155 = x2 & n34194 ;
  assign n19159 = n30049 & n19153 ;
  assign n19160 = n19155 | n19159 ;
  assign n19161 = n19149 & n19160 ;
  assign n34195 = ~n19048 ;
  assign n19162 = n19047 & n34195 ;
  assign n19163 = n19049 | n19162 ;
  assign n13059 = n9552 & n32456 ;
  assign n14664 = n9562 & n14655 ;
  assign n19164 = n10126 & n13027 ;
  assign n19165 = n10105 & n14147 ;
  assign n19166 = n19164 | n19165 ;
  assign n19167 = n14664 | n19166 ;
  assign n34196 = ~n19167 ;
  assign n19168 = x2 & n34196 ;
  assign n19169 = n30049 & n19167 ;
  assign n19170 = n19168 | n19169 ;
  assign n34197 = ~n13059 ;
  assign n19171 = n34197 & n19170 ;
  assign n19172 = n19163 | n19171 ;
  assign n19173 = n19163 & n19171 ;
  assign n34198 = ~n18731 ;
  assign n19174 = n34198 & n19041 ;
  assign n19175 = n19042 | n19174 ;
  assign n34199 = ~n18743 ;
  assign n19039 = n34199 & n19038 ;
  assign n19176 = n19039 | n19040 ;
  assign n12557 = n9552 & n32354 ;
  assign n13853 = n9562 & n32557 ;
  assign n19177 = n10105 & n32456 ;
  assign n19178 = n10126 & n13077 ;
  assign n19179 = n19177 | n19178 ;
  assign n19180 = n13853 | n19179 ;
  assign n34200 = ~n19180 ;
  assign n19181 = x2 & n34200 ;
  assign n19182 = n30049 & n19180 ;
  assign n19183 = n19181 | n19182 ;
  assign n34201 = ~n12557 ;
  assign n19184 = n34201 & n19183 ;
  assign n19185 = n19176 | n19184 ;
  assign n19500 = n19176 & n19184 ;
  assign n34202 = ~n19036 ;
  assign n19186 = n19035 & n34202 ;
  assign n19187 = n19037 | n19186 ;
  assign n34203 = ~n19032 ;
  assign n19033 = n19030 & n34203 ;
  assign n19188 = n19033 | n19034 ;
  assign n12553 = n10105 & n32354 ;
  assign n12575 = n10126 & n12570 ;
  assign n19189 = n12553 | n12575 ;
  assign n19190 = n9562 & n32356 ;
  assign n19191 = n19189 | n19190 ;
  assign n19192 = x2 & n19191 ;
  assign n19193 = n31643 & n12595 ;
  assign n34204 = ~n19193 ;
  assign n19194 = x2 & n34204 ;
  assign n19195 = n19191 | n19194 ;
  assign n34205 = ~n19192 ;
  assign n19196 = n34205 & n19195 ;
  assign n19198 = n19188 & n19196 ;
  assign n19197 = n19188 | n19196 ;
  assign n19199 = n19019 | n19020 ;
  assign n34206 = ~n19021 ;
  assign n19200 = n34206 & n19199 ;
  assign n12592 = n10105 & n12570 ;
  assign n12615 = n10126 & n12595 ;
  assign n19201 = n12592 | n12615 ;
  assign n19202 = n9562 & n12681 ;
  assign n19203 = n19201 | n19202 ;
  assign n19204 = n30049 & n19203 ;
  assign n12146 = n733 | n12136 ;
  assign n19205 = x2 & n12146 ;
  assign n34207 = ~n19203 ;
  assign n19206 = n34207 & n19205 ;
  assign n19207 = n19204 | n19206 ;
  assign n19208 = n19200 & n19207 ;
  assign n19483 = n19200 | n19207 ;
  assign n19209 = n18774 | n19013 ;
  assign n34208 = ~n19014 ;
  assign n19210 = n34208 & n19209 ;
  assign n34209 = ~n18787 ;
  assign n19211 = n34209 & n19011 ;
  assign n19212 = n19012 | n19211 ;
  assign n12203 = n9562 & n32255 ;
  assign n11854 = n9552 & n32176 ;
  assign n12174 = n10126 & n12161 ;
  assign n19213 = n11854 | n12174 ;
  assign n19214 = n10105 & n32253 ;
  assign n19215 = n19213 | n19214 ;
  assign n19216 = n12203 | n19215 ;
  assign n19217 = x2 | n19216 ;
  assign n19218 = x2 & n19216 ;
  assign n34210 = ~n19218 ;
  assign n19219 = n19217 & n34210 ;
  assign n19220 = n19212 & n19219 ;
  assign n19452 = n18799 | n19009 ;
  assign n34211 = ~n19010 ;
  assign n19453 = n34211 & n19452 ;
  assign n11443 = n9552 & n11430 ;
  assign n12665 = n9562 & n32362 ;
  assign n19454 = n10126 & n32176 ;
  assign n19455 = n10105 & n12161 ;
  assign n19456 = n19454 | n19455 ;
  assign n19457 = n12665 | n19456 ;
  assign n34212 = ~n19457 ;
  assign n19458 = x2 & n34212 ;
  assign n19459 = n30049 & n19457 ;
  assign n19460 = n19458 | n19459 ;
  assign n34213 = ~n11443 ;
  assign n19461 = n34213 & n19460 ;
  assign n19462 = n19453 & n19461 ;
  assign n19466 = n19220 | n19462 ;
  assign n11497 = n9552 & n11476 ;
  assign n11880 = n9562 & n32178 ;
  assign n19221 = n10126 & n11430 ;
  assign n19222 = n10105 & n32176 ;
  assign n19223 = n19221 | n19222 ;
  assign n19224 = n11880 | n19223 ;
  assign n34214 = ~n19224 ;
  assign n19225 = x2 & n34214 ;
  assign n19226 = n30049 & n19224 ;
  assign n19227 = n19225 | n19226 ;
  assign n34215 = ~n11497 ;
  assign n19228 = n34215 & n19227 ;
  assign n19004 = n18822 & n19003 ;
  assign n19229 = n18822 | n19003 ;
  assign n34216 = ~n19004 ;
  assign n19230 = n34216 & n19229 ;
  assign n11060 = n9552 & n10679 ;
  assign n11522 = n9562 & n11511 ;
  assign n19231 = n10126 & n10656 ;
  assign n19232 = n10105 & n11452 ;
  assign n19233 = n19231 | n19232 ;
  assign n19234 = n11522 | n19233 ;
  assign n34217 = ~n19234 ;
  assign n19235 = x2 & n34217 ;
  assign n19236 = n30049 & n19234 ;
  assign n19237 = n19235 | n19236 ;
  assign n34218 = ~n11060 ;
  assign n19238 = n34218 & n19237 ;
  assign n34219 = ~n18842 ;
  assign n19239 = n34219 & n18994 ;
  assign n19240 = n18995 | n19239 ;
  assign n19241 = n18854 | n18992 ;
  assign n34220 = ~n18993 ;
  assign n19242 = n34220 & n19241 ;
  assign n10718 = n9552 & n10703 ;
  assign n11547 = n9562 & n11536 ;
  assign n19243 = n10105 & n10679 ;
  assign n19244 = n10126 & n10681 ;
  assign n19245 = n19243 | n19244 ;
  assign n19246 = n11547 | n19245 ;
  assign n34221 = ~n19246 ;
  assign n19247 = x2 & n34221 ;
  assign n19248 = n30049 & n19246 ;
  assign n19249 = n19247 | n19248 ;
  assign n34222 = ~n10718 ;
  assign n19250 = n34222 & n19249 ;
  assign n19251 = n19242 & n19250 ;
  assign n19413 = n19242 | n19250 ;
  assign n18990 = n18866 & n18989 ;
  assign n19252 = n18866 | n18989 ;
  assign n34223 = ~n18990 ;
  assign n19253 = n34223 & n19252 ;
  assign n13160 = n9562 & n13157 ;
  assign n10715 = n10126 & n10703 ;
  assign n10748 = n9552 & n10727 ;
  assign n19254 = n10715 | n10748 ;
  assign n19255 = n10105 & n10681 ;
  assign n19256 = n19254 | n19255 ;
  assign n19257 = n13160 | n19256 ;
  assign n34224 = ~n19257 ;
  assign n19258 = x2 & n34224 ;
  assign n19259 = n30049 & n19257 ;
  assign n19260 = n19258 | n19259 ;
  assign n19262 = n19253 & n19260 ;
  assign n19261 = n19253 | n19260 ;
  assign n18987 = n18878 | n18986 ;
  assign n19263 = n18878 & n18986 ;
  assign n34225 = ~n19263 ;
  assign n19264 = n18987 & n34225 ;
  assign n13193 = n9562 & n13182 ;
  assign n19265 = n10105 & n13151 ;
  assign n19266 = n10126 & n10727 ;
  assign n19267 = n19265 | n19266 ;
  assign n19268 = n13193 | n19267 ;
  assign n19269 = x2 | n19268 ;
  assign n19270 = x2 & n19268 ;
  assign n34226 = ~n19270 ;
  assign n19271 = n19269 & n34226 ;
  assign n19272 = n9552 & n32478 ;
  assign n34227 = ~n19272 ;
  assign n19273 = n19271 & n34227 ;
  assign n19275 = n19264 & n19273 ;
  assign n19274 = n19264 | n19273 ;
  assign n19276 = n18983 | n18984 ;
  assign n34228 = ~n18985 ;
  assign n19277 = n34228 & n19276 ;
  assign n11696 = n9562 & n32125 ;
  assign n19278 = n10105 & n10727 ;
  assign n19279 = n10126 & n32478 ;
  assign n19280 = n19278 | n19279 ;
  assign n19281 = n11696 | n19280 ;
  assign n19282 = x2 | n19281 ;
  assign n19283 = x2 & n19281 ;
  assign n34229 = ~n19283 ;
  assign n19284 = n19282 & n34229 ;
  assign n19285 = n9552 & n13292 ;
  assign n34230 = ~n19285 ;
  assign n19286 = n19284 & n34230 ;
  assign n19407 = n19277 | n19286 ;
  assign n19408 = n19274 & n19407 ;
  assign n19287 = n19277 & n19286 ;
  assign n19288 = n18898 | n18977 ;
  assign n34231 = ~n18978 ;
  assign n19289 = n34231 & n19288 ;
  assign n10811 = n9552 & n31998 ;
  assign n13239 = n9562 & n32477 ;
  assign n19290 = n10105 & n32478 ;
  assign n19291 = n10126 & n13292 ;
  assign n19292 = n19290 | n19291 ;
  assign n19293 = n13239 | n19292 ;
  assign n34232 = ~n19293 ;
  assign n19294 = x2 & n34232 ;
  assign n19295 = n30049 & n19293 ;
  assign n19296 = n19294 | n19295 ;
  assign n34233 = ~n10811 ;
  assign n19297 = n34233 & n19296 ;
  assign n19299 = n19289 | n19297 ;
  assign n13280 = n9562 & n32482 ;
  assign n19394 = n10105 & n13292 ;
  assign n19395 = n10126 & n31998 ;
  assign n19396 = n19394 | n19395 ;
  assign n19397 = n13280 | n19396 ;
  assign n19398 = n30049 & n19397 ;
  assign n10828 = n31643 & n10818 ;
  assign n34234 = ~n10828 ;
  assign n19399 = x2 & n34234 ;
  assign n34235 = ~n19397 ;
  assign n19400 = n34235 & n19399 ;
  assign n19401 = n19398 | n19400 ;
  assign n18975 = n18917 & n18974 ;
  assign n19300 = n18917 | n18974 ;
  assign n34236 = ~n18975 ;
  assign n19301 = n34236 & n19300 ;
  assign n10883 = n9552 & n10865 ;
  assign n13387 = n9562 & n13382 ;
  assign n19302 = n10105 & n10818 ;
  assign n19303 = n10126 & n10841 ;
  assign n19304 = n19302 | n19303 ;
  assign n19305 = n13387 | n19304 ;
  assign n34237 = ~n19305 ;
  assign n19306 = x2 & n34237 ;
  assign n19307 = n30049 & n19305 ;
  assign n19308 = n19306 | n19307 ;
  assign n34238 = ~n10883 ;
  assign n19309 = n34238 & n19308 ;
  assign n34239 = ~n18946 ;
  assign n18948 = n10992 & n34239 ;
  assign n18945 = x5 & n18944 ;
  assign n34240 = ~x6 ;
  assign n19311 = n34240 & n18945 ;
  assign n34241 = ~n18945 ;
  assign n19310 = x6 & n34241 ;
  assign n19312 = n10992 | n19310 ;
  assign n19313 = n19311 | n19312 ;
  assign n34242 = ~n18948 ;
  assign n19314 = n34242 & n19313 ;
  assign n34243 = ~n18955 ;
  assign n19315 = n34243 & n19314 ;
  assign n34244 = ~n19314 ;
  assign n19316 = n18955 & n34244 ;
  assign n19317 = n19315 | n19316 ;
  assign n19318 = x5 & n18937 ;
  assign n19319 = n18943 & n19318 ;
  assign n19320 = n18943 | n19318 ;
  assign n34245 = ~n19319 ;
  assign n19321 = n34245 & n19320 ;
  assign n13528 = n9562 & n32502 ;
  assign n10896 = n10126 & n10892 ;
  assign n10938 = n9552 & n32503 ;
  assign n19322 = n10896 | n10938 ;
  assign n19323 = n10105 & n10865 ;
  assign n19324 = n19322 | n19323 ;
  assign n19325 = n13528 | n19324 ;
  assign n19326 = x2 | n19325 ;
  assign n19327 = x2 & n19325 ;
  assign n34246 = ~n19327 ;
  assign n19328 = n19326 & n34246 ;
  assign n19329 = n19321 & n19328 ;
  assign n19358 = n19321 | n19328 ;
  assign n19330 = n18932 & n18936 ;
  assign n34247 = ~n19330 ;
  assign n19331 = n18937 & n34247 ;
  assign n10952 = n9552 & n10940 ;
  assign n13767 = n9562 & n13756 ;
  assign n19332 = n10105 & n10892 ;
  assign n19333 = n10126 & n32503 ;
  assign n19334 = n19332 | n19333 ;
  assign n19335 = n13767 | n19334 ;
  assign n34248 = ~n19335 ;
  assign n19336 = x2 & n34248 ;
  assign n19337 = n30049 & n19335 ;
  assign n19338 = n19336 | n19337 ;
  assign n34249 = ~n10952 ;
  assign n19339 = n34249 & n19338 ;
  assign n19341 = n19331 & n19339 ;
  assign n19340 = n19331 | n19339 ;
  assign n13692 = n9562 & n13690 ;
  assign n10955 = n10126 & n10940 ;
  assign n10986 = n9552 & n31995 ;
  assign n19342 = n10955 | n10986 ;
  assign n19343 = n10105 & n32503 ;
  assign n19344 = n19342 | n19343 ;
  assign n19345 = n13692 | n19344 ;
  assign n19349 = x3 & n32507 ;
  assign n34250 = ~n19349 ;
  assign n19350 = x2 & n34250 ;
  assign n10972 = x0 & n10940 ;
  assign n19346 = x1 | n9562 ;
  assign n19347 = n31995 & n19346 ;
  assign n19348 = n10972 | n19347 ;
  assign n19351 = n10992 & n19348 ;
  assign n34251 = ~n19351 ;
  assign n19352 = n19350 & n34251 ;
  assign n19353 = n19345 | n19352 ;
  assign n19354 = n30049 & n19349 ;
  assign n34252 = ~n19354 ;
  assign n19355 = n19345 & n34252 ;
  assign n34253 = ~n19355 ;
  assign n19356 = n19353 & n34253 ;
  assign n19357 = n19340 & n19356 ;
  assign n19359 = n19341 | n19357 ;
  assign n19360 = n19358 & n19359 ;
  assign n19361 = n19329 | n19360 ;
  assign n19362 = n19317 & n19361 ;
  assign n10862 = n10105 & n10841 ;
  assign n10887 = n10126 & n10865 ;
  assign n19363 = n10862 | n10887 ;
  assign n19364 = n9562 & n13456 ;
  assign n19365 = n19363 | n19364 ;
  assign n19366 = x2 & n19365 ;
  assign n19367 = n9552 & n10892 ;
  assign n19368 = x2 | n19365 ;
  assign n34254 = ~n19367 ;
  assign n19369 = n34254 & n19368 ;
  assign n34255 = ~n19366 ;
  assign n19370 = n34255 & n19369 ;
  assign n19371 = n19317 | n19361 ;
  assign n19372 = n19370 & n19371 ;
  assign n19373 = n19362 | n19372 ;
  assign n19375 = n19309 | n19373 ;
  assign n19374 = n19309 & n19373 ;
  assign n18970 = n18967 & n18968 ;
  assign n19376 = n18967 | n18968 ;
  assign n34256 = ~n18970 ;
  assign n19377 = n34256 & n19376 ;
  assign n19378 = n19374 | n19377 ;
  assign n19379 = n19375 & n19378 ;
  assign n13327 = n9562 & n32488 ;
  assign n10840 = n10126 & n10818 ;
  assign n10863 = n9552 & n10841 ;
  assign n19380 = n10840 | n10863 ;
  assign n19381 = n10105 & n31998 ;
  assign n19382 = n19380 | n19381 ;
  assign n19383 = n13327 | n19382 ;
  assign n19384 = x2 | n19383 ;
  assign n19385 = x2 & n19383 ;
  assign n34257 = ~n19385 ;
  assign n19386 = n19384 & n34257 ;
  assign n19387 = n19379 & n19386 ;
  assign n18972 = n18931 & n18971 ;
  assign n19388 = n18931 | n18971 ;
  assign n34258 = ~n18972 ;
  assign n19389 = n34258 & n19388 ;
  assign n19390 = n19387 | n19389 ;
  assign n19391 = n19379 | n19386 ;
  assign n19392 = n19390 & n19391 ;
  assign n19402 = n19301 | n19392 ;
  assign n19403 = n19401 & n19402 ;
  assign n19298 = n19289 & n19297 ;
  assign n19393 = n19301 & n19392 ;
  assign n19404 = n19298 | n19393 ;
  assign n19405 = n19403 | n19404 ;
  assign n19406 = n19299 & n19405 ;
  assign n19409 = n19287 | n19406 ;
  assign n19410 = n19408 & n19409 ;
  assign n19411 = n19275 | n19410 ;
  assign n19412 = n19261 & n19411 ;
  assign n19414 = n19262 | n19412 ;
  assign n19415 = n19413 & n19414 ;
  assign n19416 = n19251 | n19415 ;
  assign n19417 = n19240 & n19416 ;
  assign n10673 = n10105 & n10656 ;
  assign n11062 = n10126 & n10679 ;
  assign n19418 = n10673 | n11062 ;
  assign n19419 = n9562 & n11030 ;
  assign n19420 = n19418 | n19419 ;
  assign n19421 = x2 & n19420 ;
  assign n19422 = n9552 & n10681 ;
  assign n19423 = x2 | n19420 ;
  assign n34259 = ~n19422 ;
  assign n19424 = n34259 & n19423 ;
  assign n34260 = ~n19421 ;
  assign n19425 = n34260 & n19424 ;
  assign n19426 = n19240 | n19416 ;
  assign n19427 = n19425 & n19426 ;
  assign n19428 = n19417 | n19427 ;
  assign n19430 = n19238 | n19428 ;
  assign n19429 = n19238 & n19428 ;
  assign n34261 = ~n19001 ;
  assign n19431 = n19000 & n34261 ;
  assign n19432 = n19002 | n19431 ;
  assign n19433 = n19429 | n19432 ;
  assign n19434 = n19430 & n19433 ;
  assign n19435 = n19230 & n19434 ;
  assign n11464 = n9562 & n11463 ;
  assign n19436 = n10105 & n11430 ;
  assign n19437 = n10126 & n11452 ;
  assign n19438 = n19436 | n19437 ;
  assign n19439 = n11464 | n19438 ;
  assign n19440 = x2 & n19439 ;
  assign n19441 = n9552 & n10656 ;
  assign n19442 = x2 | n19439 ;
  assign n34262 = ~n19441 ;
  assign n19443 = n34262 & n19442 ;
  assign n34263 = ~n19440 ;
  assign n19444 = n34263 & n19443 ;
  assign n19445 = n19230 | n19434 ;
  assign n19446 = n19444 & n19445 ;
  assign n19447 = n19435 | n19446 ;
  assign n19448 = n19228 & n19447 ;
  assign n34264 = ~n19007 ;
  assign n19449 = n19006 & n34264 ;
  assign n19450 = n19008 | n19449 ;
  assign n19451 = n19448 | n19450 ;
  assign n19463 = n19228 | n19447 ;
  assign n19464 = n19453 | n19461 ;
  assign n19465 = n19463 & n19464 ;
  assign n19467 = n19451 & n19465 ;
  assign n19468 = n19466 | n19467 ;
  assign n19469 = n19212 | n19219 ;
  assign n19470 = n19468 & n19469 ;
  assign n19471 = n19210 | n19470 ;
  assign n13832 = n9562 & n32550 ;
  assign n19472 = n10126 & n32253 ;
  assign n19473 = n10105 & n12595 ;
  assign n19474 = n19472 | n19473 ;
  assign n19475 = n13832 | n19474 ;
  assign n19476 = x2 | n19475 ;
  assign n19477 = x2 & n19475 ;
  assign n34265 = ~n19477 ;
  assign n19478 = n19476 & n34265 ;
  assign n19479 = n9552 & n12161 ;
  assign n34266 = ~n19479 ;
  assign n19480 = n19478 & n34266 ;
  assign n19481 = n19471 & n19480 ;
  assign n19482 = n19210 & n19470 ;
  assign n19484 = n19481 | n19482 ;
  assign n19485 = n19483 & n19484 ;
  assign n19486 = n19208 | n19485 ;
  assign n19487 = n19197 & n19486 ;
  assign n19488 = n19198 | n19487 ;
  assign n19490 = n19187 | n19488 ;
  assign n19489 = n19187 & n19488 ;
  assign n14255 = n9562 & n32641 ;
  assign n19491 = n10126 & n32354 ;
  assign n19492 = n10105 & n13077 ;
  assign n19493 = n19491 | n19492 ;
  assign n19494 = n14255 | n19493 ;
  assign n19495 = n30049 & n19494 ;
  assign n12578 = n31643 & n12570 ;
  assign n34267 = ~n12578 ;
  assign n19496 = x2 & n34267 ;
  assign n34268 = ~n19494 ;
  assign n19497 = n34268 & n19496 ;
  assign n19498 = n19495 | n19497 ;
  assign n19499 = n19489 | n19498 ;
  assign n19501 = n19490 & n19499 ;
  assign n19502 = n19500 | n19501 ;
  assign n19503 = n19185 & n19502 ;
  assign n19505 = n19175 | n19503 ;
  assign n19504 = n19175 & n19503 ;
  assign n13113 = n9562 & n32455 ;
  assign n19506 = n10105 & n13027 ;
  assign n19507 = n10126 & n32456 ;
  assign n19508 = n19506 | n19507 ;
  assign n19509 = n13113 | n19508 ;
  assign n19510 = n30049 & n19509 ;
  assign n13094 = n31643 & n13077 ;
  assign n34269 = ~n13094 ;
  assign n19511 = x2 & n34269 ;
  assign n34270 = ~n19509 ;
  assign n19512 = n34270 & n19511 ;
  assign n19513 = n19510 | n19512 ;
  assign n19514 = n19504 | n19513 ;
  assign n19515 = n19505 & n19514 ;
  assign n19516 = n19173 | n19515 ;
  assign n19517 = n19172 & n19516 ;
  assign n19518 = n19161 | n19517 ;
  assign n19519 = n19158 & n19518 ;
  assign n34271 = ~n18708 ;
  assign n19520 = n34271 & n18709 ;
  assign n34272 = ~n19520 ;
  assign n19521 = n19063 & n34272 ;
  assign n34273 = ~n19063 ;
  assign n19522 = n34273 & n19520 ;
  assign n19523 = n19521 | n19522 ;
  assign n19525 = n19519 & n19523 ;
  assign n19524 = n19519 | n19523 ;
  assign n14166 = n9552 & n14147 ;
  assign n14191 = n9562 & n14183 ;
  assign n19526 = n10105 & n14196 ;
  assign n19527 = n10126 & n14295 ;
  assign n19528 = n19526 | n19527 ;
  assign n19529 = n14191 | n19528 ;
  assign n19530 = x2 | n19529 ;
  assign n34274 = ~n14166 ;
  assign n19531 = n34274 & n19530 ;
  assign n19532 = x2 & n19529 ;
  assign n34275 = ~n19532 ;
  assign n19533 = n19531 & n34275 ;
  assign n19534 = n19524 & n19533 ;
  assign n19535 = n19525 | n19534 ;
  assign n19536 = n19147 & n19535 ;
  assign n14138 = n9552 & n14124 ;
  assign n14973 = n9562 & n14965 ;
  assign n19537 = n10126 & n14196 ;
  assign n19538 = n10105 & n14536 ;
  assign n19539 = n19537 | n19538 ;
  assign n19540 = n14973 | n19539 ;
  assign n34276 = ~n19540 ;
  assign n19541 = x2 & n34276 ;
  assign n19542 = n30049 & n19540 ;
  assign n19543 = n19541 | n19542 ;
  assign n34277 = ~n14138 ;
  assign n19544 = n34277 & n19543 ;
  assign n19545 = n19147 | n19535 ;
  assign n19546 = n19544 & n19545 ;
  assign n19547 = n19536 | n19546 ;
  assign n14117 = n9552 & n14101 ;
  assign n14684 = n9562 & n32735 ;
  assign n19548 = n10105 & n32706 ;
  assign n19549 = n10126 & n14536 ;
  assign n19550 = n19548 | n19549 ;
  assign n19551 = n14684 | n19550 ;
  assign n34278 = ~n19551 ;
  assign n19552 = x2 & n34278 ;
  assign n19553 = n30049 & n19551 ;
  assign n19554 = n19552 | n19553 ;
  assign n34279 = ~n14117 ;
  assign n19555 = n34279 & n19554 ;
  assign n19556 = n19547 & n19555 ;
  assign n34280 = ~n18687 ;
  assign n19070 = n34280 & n19069 ;
  assign n34281 = ~n19069 ;
  assign n19557 = n18687 & n34281 ;
  assign n19558 = n19070 | n19557 ;
  assign n19559 = n19547 | n19555 ;
  assign n34282 = ~n19556 ;
  assign n19560 = n34282 & n19559 ;
  assign n34283 = ~n19558 ;
  assign n19561 = n34283 & n19560 ;
  assign n19562 = n19556 | n19561 ;
  assign n34284 = ~n19145 ;
  assign n19564 = n34284 & n19562 ;
  assign n19565 = n19143 | n19564 ;
  assign n34285 = ~n19565 ;
  assign n19567 = n19132 & n34285 ;
  assign n34286 = ~n19567 ;
  assign n19568 = n19131 & n34286 ;
  assign n14506 = n9552 & n32707 ;
  assign n15120 = n9562 & n15111 ;
  assign n19569 = n10105 & n32856 ;
  assign n19570 = n10126 & n15081 ;
  assign n19571 = n19569 | n19570 ;
  assign n19572 = n15120 | n19571 ;
  assign n34287 = ~n19572 ;
  assign n19573 = x2 & n34287 ;
  assign n19574 = n30049 & n19572 ;
  assign n19575 = n19573 | n19574 ;
  assign n34288 = ~n14506 ;
  assign n19576 = n34288 & n19575 ;
  assign n19578 = n19568 & n19576 ;
  assign n19078 = n18649 & n19077 ;
  assign n34289 = ~n19078 ;
  assign n19579 = n34289 & n19079 ;
  assign n19580 = n19568 | n19576 ;
  assign n34290 = ~n19579 ;
  assign n19581 = n34290 & n19580 ;
  assign n19582 = n19578 | n19581 ;
  assign n15087 = n9552 & n15081 ;
  assign n15191 = n9562 & n32875 ;
  assign n19583 = n10126 & n32856 ;
  assign n19584 = n10105 & n32876 ;
  assign n19585 = n19583 | n19584 ;
  assign n19586 = n15191 | n19585 ;
  assign n34291 = ~n19586 ;
  assign n19587 = x2 & n34291 ;
  assign n19588 = n30049 & n19586 ;
  assign n19589 = n19587 | n19588 ;
  assign n34292 = ~n15087 ;
  assign n19590 = n34292 & n19589 ;
  assign n19591 = n19582 & n19590 ;
  assign n34293 = ~n18637 ;
  assign n19081 = n34293 & n19080 ;
  assign n34294 = ~n19080 ;
  assign n19592 = n18637 & n34294 ;
  assign n19593 = n19081 | n19592 ;
  assign n19594 = n19582 | n19590 ;
  assign n34295 = ~n19591 ;
  assign n19595 = n34295 & n19594 ;
  assign n34296 = ~n19593 ;
  assign n19596 = n34296 & n19595 ;
  assign n19597 = n19591 | n19596 ;
  assign n19599 = n19119 & n19597 ;
  assign n34297 = ~n18625 ;
  assign n19600 = n34297 & n19083 ;
  assign n19601 = n19084 | n19600 ;
  assign n19598 = n19119 | n19597 ;
  assign n34298 = ~n19599 ;
  assign n19602 = n19598 & n34298 ;
  assign n19603 = n19601 & n19602 ;
  assign n19604 = n19599 | n19603 ;
  assign n34299 = ~n19604 ;
  assign n19605 = n19112 & n34299 ;
  assign n34300 = ~n19605 ;
  assign n19606 = n19110 & n34300 ;
  assign n15225 = n10126 & n15221 ;
  assign n19607 = n10105 | n15225 ;
  assign n19608 = x0 & n15516 ;
  assign n19609 = n19607 | n19608 ;
  assign n19610 = x2 & n19609 ;
  assign n19611 = n733 | n15252 ;
  assign n19612 = x2 & n19611 ;
  assign n19613 = n19609 | n19612 ;
  assign n34301 = ~n19610 ;
  assign n19614 = n34301 & n19613 ;
  assign n19616 = n19606 & n19614 ;
  assign n19089 = n18601 & n19088 ;
  assign n19617 = n18601 | n19088 ;
  assign n34302 = ~n19089 ;
  assign n19618 = n34302 & n19617 ;
  assign n34303 = ~n19614 ;
  assign n19615 = n19606 & n34303 ;
  assign n34304 = ~n19606 ;
  assign n19619 = n34304 & n19614 ;
  assign n19620 = n19615 | n19619 ;
  assign n19621 = n19618 & n19620 ;
  assign n19622 = n19616 | n19621 ;
  assign n19624 = n19099 & n19622 ;
  assign n19623 = n19099 | n19622 ;
  assign n34305 = ~n19624 ;
  assign n19625 = n19623 & n34305 ;
  assign n15236 = n9552 & n32883 ;
  assign n19626 = n734 | n15236 ;
  assign n19628 = n19625 & n19626 ;
  assign n19629 = n19624 | n19628 ;
  assign n19630 = n19097 | n19629 ;
  assign n19631 = n19096 & n19630 ;
  assign n34306 = ~n18574 ;
  assign n19632 = n34306 & n19631 ;
  assign n19634 = n18573 | n19632 ;
  assign n34307 = ~n19634 ;
  assign n19635 = n18555 & n34307 ;
  assign n34308 = ~n19635 ;
  assign n19637 = n18554 & n34308 ;
  assign n19640 = n18038 | n19637 ;
  assign n34309 = ~n18036 ;
  assign n19641 = n34309 & n19640 ;
  assign n19642 = n17545 | n19641 ;
  assign n34310 = ~n17543 ;
  assign n19643 = n34310 & n19642 ;
  assign n34311 = ~n19643 ;
  assign n19646 = n17088 & n34311 ;
  assign n34312 = ~n19646 ;
  assign n19647 = n17086 & n34312 ;
  assign n19648 = n16658 | n19647 ;
  assign n34313 = ~n16657 ;
  assign n19649 = n34313 & n19648 ;
  assign n19652 = n16260 | n19649 ;
  assign n34314 = ~n16258 ;
  assign n19653 = n34314 & n19652 ;
  assign n19654 = n15894 | n19653 ;
  assign n34315 = ~n15893 ;
  assign n19655 = n34315 & n19654 ;
  assign n34316 = ~n15561 ;
  assign n19656 = n34316 & n19655 ;
  assign n34317 = ~n19655 ;
  assign n19658 = n15561 & n34317 ;
  assign n19659 = n19656 | n19658 ;
  assign n19681 = n15894 & n19653 ;
  assign n34318 = ~n19681 ;
  assign n19682 = n19654 & n34318 ;
  assign n34319 = ~n16260 ;
  assign n19650 = n34319 & n19649 ;
  assign n34320 = ~n19649 ;
  assign n19704 = n16260 & n34320 ;
  assign n19705 = n19650 | n19704 ;
  assign n19728 = n16658 & n19647 ;
  assign n34321 = ~n19728 ;
  assign n19729 = n19648 & n34321 ;
  assign n19644 = n17088 & n19643 ;
  assign n19751 = n17088 | n19643 ;
  assign n34322 = ~n19644 ;
  assign n19752 = n34322 & n19751 ;
  assign n34323 = ~n17545 ;
  assign n19774 = n34323 & n19641 ;
  assign n34324 = ~n19641 ;
  assign n19775 = n17545 & n34324 ;
  assign n19776 = n19774 | n19775 ;
  assign n34325 = ~n18038 ;
  assign n19638 = n34325 & n19637 ;
  assign n34326 = ~n19637 ;
  assign n19799 = n18038 & n34326 ;
  assign n19800 = n19638 | n19799 ;
  assign n19636 = n18555 | n19634 ;
  assign n19823 = n18555 & n19634 ;
  assign n34327 = ~n19823 ;
  assign n19824 = n19636 & n34327 ;
  assign n34328 = ~n19094 ;
  assign n19095 = n18576 & n34328 ;
  assign n34329 = ~n18576 ;
  assign n20063 = n34329 & n19094 ;
  assign n20064 = n19095 | n20063 ;
  assign n20065 = n19629 & n20064 ;
  assign n20066 = n19629 | n20064 ;
  assign n34330 = ~n20065 ;
  assign n20067 = n34330 & n20066 ;
  assign n19627 = n19625 | n19626 ;
  assign n34331 = ~n19628 ;
  assign n19846 = n19627 & n34331 ;
  assign n19869 = n19618 | n19620 ;
  assign n34332 = ~n19621 ;
  assign n19870 = n34332 & n19869 ;
  assign n34333 = ~n19112 ;
  assign n19892 = n34333 & n19604 ;
  assign n19893 = n19605 | n19892 ;
  assign n19916 = n19601 | n19602 ;
  assign n34334 = ~n19603 ;
  assign n19917 = n34334 & n19916 ;
  assign n34335 = ~n19595 ;
  assign n19941 = n19593 & n34335 ;
  assign n19942 = n19596 | n19941 ;
  assign n34336 = ~n19568 ;
  assign n19577 = n34336 & n19576 ;
  assign n34337 = ~n19576 ;
  assign n19964 = n19568 & n34337 ;
  assign n19965 = n19577 | n19964 ;
  assign n19966 = n19579 & n19965 ;
  assign n19967 = n19579 | n19965 ;
  assign n34338 = ~n19966 ;
  assign n19968 = n34338 & n19967 ;
  assign n34339 = ~n19132 ;
  assign n19566 = n34339 & n19565 ;
  assign n19991 = n19566 | n19567 ;
  assign n34340 = ~n19562 ;
  assign n19563 = n19145 & n34340 ;
  assign n20022 = n19563 | n19564 ;
  assign n34341 = ~n19560 ;
  assign n20037 = n19558 & n34341 ;
  assign n20038 = n19561 | n20037 ;
  assign n20052 = n20022 | n20038 ;
  assign n34342 = ~n19991 ;
  assign n20054 = n34342 & n20052 ;
  assign n20056 = n19968 | n20054 ;
  assign n20057 = n19942 & n20056 ;
  assign n34343 = ~n20057 ;
  assign n20059 = n19917 & n34343 ;
  assign n20060 = n19893 | n20059 ;
  assign n20062 = n19870 & n20060 ;
  assign n20090 = n19846 | n20062 ;
  assign n20091 = n20067 & n20090 ;
  assign n34344 = ~n19631 ;
  assign n20092 = n18574 & n34344 ;
  assign n20093 = n19632 | n20092 ;
  assign n34345 = ~n20091 ;
  assign n20116 = n34345 & n20093 ;
  assign n34346 = ~n20116 ;
  assign n20118 = n19824 & n34346 ;
  assign n34347 = ~n20118 ;
  assign n20119 = n19800 & n34347 ;
  assign n20121 = n19776 | n20119 ;
  assign n34348 = ~n19752 ;
  assign n20122 = n34348 & n20121 ;
  assign n20124 = n19729 | n20122 ;
  assign n20125 = n19705 & n20124 ;
  assign n34349 = ~n19682 ;
  assign n20126 = n34349 & n20125 ;
  assign n34350 = ~n20022 ;
  assign n20024 = n19991 & n34350 ;
  assign n34351 = ~n20024 ;
  assign n20127 = n19968 & n34351 ;
  assign n20128 = n19942 | n20127 ;
  assign n34352 = ~n19917 ;
  assign n20129 = n34352 & n20128 ;
  assign n34353 = ~n20129 ;
  assign n20130 = n19893 & n34353 ;
  assign n20131 = n19870 | n20130 ;
  assign n20132 = n19846 & n20131 ;
  assign n20133 = n20067 | n20132 ;
  assign n34354 = ~n20093 ;
  assign n20135 = n34354 & n20133 ;
  assign n20136 = n19824 | n20135 ;
  assign n34355 = ~n19800 ;
  assign n20137 = n34355 & n20136 ;
  assign n34356 = ~n20137 ;
  assign n20138 = n19776 & n34356 ;
  assign n34357 = ~n20138 ;
  assign n20140 = n19752 & n34357 ;
  assign n34358 = ~n20140 ;
  assign n20141 = n19729 & n34358 ;
  assign n20142 = n19705 | n20141 ;
  assign n34359 = ~n20142 ;
  assign n20143 = n19682 & n34359 ;
  assign n20144 = n20126 | n20143 ;
  assign n34360 = ~n19659 ;
  assign n20145 = n34360 & n20144 ;
  assign n34361 = ~n20144 ;
  assign n20146 = n19659 & n34361 ;
  assign n20147 = n20145 | n20146 ;
  assign n34362 = ~n20147 ;
  assign n20149 = n37300 & n34362 ;
  assign n19695 = n5144 & n34349 ;
  assign n34363 = ~n19705 ;
  assign n19713 = n5166 & n34363 ;
  assign n20161 = n19695 | n19713 ;
  assign n19657 = n15561 & n19655 ;
  assign n20159 = n15561 | n19655 ;
  assign n34364 = ~n19657 ;
  assign n20160 = n34364 & n20159 ;
  assign n34365 = ~n20160 ;
  assign n20162 = n5191 & n34365 ;
  assign n20163 = n20161 | n20162 ;
  assign n20164 = n20149 | n20163 ;
  assign n34366 = ~n20164 ;
  assign n20165 = x17 & n34366 ;
  assign n20166 = n30580 & n20164 ;
  assign n20167 = n20165 | n20166 ;
  assign n34367 = ~n20038 ;
  assign n20168 = n108 & n34367 ;
  assign n20050 = n891 & n34367 ;
  assign n20047 = n34350 & n20038 ;
  assign n20169 = n20022 & n34367 ;
  assign n20170 = n20047 | n20169 ;
  assign n20171 = n895 & n20170 ;
  assign n20182 = n894 & n34350 ;
  assign n20183 = n2849 & n34367 ;
  assign n20184 = n20182 | n20183 ;
  assign n20185 = n20171 | n20184 ;
  assign n20186 = n20050 | n20185 ;
  assign n20187 = x29 & n20186 ;
  assign n20000 = n894 & n19991 ;
  assign n20192 = n2849 & n34350 ;
  assign n20193 = n2861 & n34367 ;
  assign n20194 = n20192 | n20193 ;
  assign n20195 = n20000 | n20194 ;
  assign n20048 = n19991 & n20047 ;
  assign n20188 = n19991 | n20047 ;
  assign n34368 = ~n20048 ;
  assign n20189 = n34368 & n20188 ;
  assign n20196 = n895 & n20189 ;
  assign n20197 = n20195 | n20196 ;
  assign n20199 = n20187 | n20197 ;
  assign n34369 = ~n20199 ;
  assign n20200 = x29 & n34369 ;
  assign n20202 = n20168 | n20200 ;
  assign n20180 = n19991 & n20022 ;
  assign n20203 = n19991 | n20052 ;
  assign n34370 = ~n20180 ;
  assign n20204 = n34370 & n20203 ;
  assign n20205 = n19968 | n20204 ;
  assign n20206 = n19968 & n20204 ;
  assign n34371 = ~n20206 ;
  assign n20207 = n20205 & n34371 ;
  assign n20208 = n895 & n20207 ;
  assign n20016 = n2849 & n19991 ;
  assign n20031 = n2861 & n34350 ;
  assign n20218 = n20016 | n20031 ;
  assign n34372 = ~n19968 ;
  assign n20219 = n894 & n34372 ;
  assign n20220 = n20218 | n20219 ;
  assign n20221 = n20208 | n20220 ;
  assign n34373 = ~n20221 ;
  assign n20222 = x29 & n34373 ;
  assign n20223 = n30024 & n20221 ;
  assign n20224 = n20222 | n20223 ;
  assign n20225 = n20202 & n20224 ;
  assign n20049 = n108 & n20047 ;
  assign n34374 = ~n20052 ;
  assign n20053 = n6562 & n34374 ;
  assign n20227 = n20049 | n20053 ;
  assign n20181 = n6561 & n20022 ;
  assign n20226 = n3329 | n20181 ;
  assign n20228 = n34367 & n20226 ;
  assign n20229 = n20227 | n20228 ;
  assign n20230 = n2472 | n5613 ;
  assign n20231 = n12064 | n12749 ;
  assign n20232 = n20230 | n20231 ;
  assign n20233 = n659 | n858 ;
  assign n20234 = n2517 | n3016 ;
  assign n20235 = n20233 | n20234 ;
  assign n20236 = n214 | n245 ;
  assign n20237 = n368 | n622 ;
  assign n20238 = n20236 | n20237 ;
  assign n20239 = n1853 | n20238 ;
  assign n20240 = n20235 | n20239 ;
  assign n20241 = n282 | n395 ;
  assign n20242 = n401 | n407 ;
  assign n20243 = n20241 | n20242 ;
  assign n20244 = n1764 | n20243 ;
  assign n34375 = ~n20244 ;
  assign n20245 = n2557 & n34375 ;
  assign n34376 = ~n20240 ;
  assign n20246 = n34376 & n20245 ;
  assign n34377 = ~n20232 ;
  assign n20247 = n34377 & n20246 ;
  assign n20248 = n2282 | n2746 ;
  assign n20249 = n3040 | n20248 ;
  assign n20250 = n216 | n276 ;
  assign n20251 = n349 | n20250 ;
  assign n20252 = n2016 | n2030 ;
  assign n20253 = n20251 | n20252 ;
  assign n20254 = n1463 | n11230 ;
  assign n20255 = n20253 | n20254 ;
  assign n20256 = n20249 | n20255 ;
  assign n20257 = n1969 | n3743 ;
  assign n20258 = n13711 | n20257 ;
  assign n20259 = n1041 | n1177 ;
  assign n20260 = n12723 | n20259 ;
  assign n20261 = n478 | n823 ;
  assign n20262 = n11222 | n20261 ;
  assign n20263 = n372 | n529 ;
  assign n20264 = n150 | n20263 ;
  assign n20265 = n678 | n20264 ;
  assign n20266 = n20262 | n20265 ;
  assign n20267 = n20260 | n20266 ;
  assign n20268 = n20258 | n20267 ;
  assign n20269 = n20256 | n20268 ;
  assign n34378 = ~n20269 ;
  assign n20270 = n20247 & n34378 ;
  assign n34379 = ~n13414 ;
  assign n20271 = n34379 & n20270 ;
  assign n20272 = n20229 & n20271 ;
  assign n20273 = n20229 | n20271 ;
  assign n34380 = ~n20272 ;
  assign n20274 = n34380 & n20273 ;
  assign n20055 = n34372 & n20054 ;
  assign n20275 = n19968 & n20024 ;
  assign n20276 = n20055 | n20275 ;
  assign n34381 = ~n19942 ;
  assign n20277 = n34381 & n20276 ;
  assign n34382 = ~n20276 ;
  assign n20278 = n19942 & n34382 ;
  assign n20279 = n20277 | n20278 ;
  assign n34383 = ~n20279 ;
  assign n20282 = n895 & n34383 ;
  assign n19979 = n2849 & n34372 ;
  assign n19997 = n2861 & n19991 ;
  assign n20292 = n19979 | n19997 ;
  assign n20293 = n894 & n34381 ;
  assign n20294 = n20292 | n20293 ;
  assign n20295 = n20282 | n20294 ;
  assign n20296 = x29 | n20295 ;
  assign n20297 = x29 & n20295 ;
  assign n34384 = ~n20297 ;
  assign n20298 = n20296 & n34384 ;
  assign n34385 = ~n20274 ;
  assign n20299 = n34385 & n20298 ;
  assign n34386 = ~n20298 ;
  assign n20300 = n20274 & n34386 ;
  assign n20301 = n20299 | n20300 ;
  assign n34387 = ~n20301 ;
  assign n20302 = n20225 & n34387 ;
  assign n34388 = ~n20225 ;
  assign n20304 = n34388 & n20301 ;
  assign n20305 = n20302 | n20304 ;
  assign n34389 = ~n19893 ;
  assign n20306 = n34389 & n20059 ;
  assign n20307 = n19893 & n20129 ;
  assign n20308 = n20306 | n20307 ;
  assign n20309 = n19870 & n20308 ;
  assign n20310 = n19870 | n20308 ;
  assign n34390 = ~n20309 ;
  assign n20311 = n34390 & n20310 ;
  assign n20312 = n3791 & n20311 ;
  assign n19902 = n3802 & n19893 ;
  assign n19925 = n209 & n19917 ;
  assign n20323 = n19902 | n19925 ;
  assign n20324 = n3818 & n19870 ;
  assign n20325 = n20323 | n20324 ;
  assign n20326 = n20312 | n20325 ;
  assign n20327 = x26 | n20326 ;
  assign n20328 = x26 & n20326 ;
  assign n34391 = ~n20328 ;
  assign n20329 = n20327 & n34391 ;
  assign n34392 = ~n20329 ;
  assign n20331 = n20305 & n34392 ;
  assign n20330 = n20305 & n20329 ;
  assign n20332 = n20305 | n20329 ;
  assign n34393 = ~n20330 ;
  assign n20333 = n34393 & n20332 ;
  assign n20201 = n20168 & n20200 ;
  assign n34394 = ~n20201 ;
  assign n20334 = n34394 & n20202 ;
  assign n34395 = ~n20224 ;
  assign n20335 = n34395 & n20334 ;
  assign n34396 = ~n20334 ;
  assign n20336 = n20224 & n34396 ;
  assign n20337 = n20335 | n20336 ;
  assign n20058 = n19917 & n20057 ;
  assign n20338 = n19917 | n20128 ;
  assign n34397 = ~n20058 ;
  assign n20339 = n34397 & n20338 ;
  assign n34398 = ~n20339 ;
  assign n20340 = n19893 & n34398 ;
  assign n20341 = n34389 & n20339 ;
  assign n20342 = n20340 | n20341 ;
  assign n34399 = ~n20342 ;
  assign n20343 = n3791 & n34399 ;
  assign n19923 = n3802 & n19917 ;
  assign n19956 = n209 & n34381 ;
  assign n20353 = n19923 | n19956 ;
  assign n20354 = n3818 & n19893 ;
  assign n20355 = n20353 | n20354 ;
  assign n20356 = n20343 | n20355 ;
  assign n20357 = x26 | n20356 ;
  assign n20358 = x26 & n20356 ;
  assign n34400 = ~n20358 ;
  assign n20359 = n20357 & n34400 ;
  assign n20361 = n20337 | n20359 ;
  assign n20360 = n20337 & n20359 ;
  assign n34401 = ~n20360 ;
  assign n20362 = n34401 & n20361 ;
  assign n20198 = n20187 & n20197 ;
  assign n34402 = ~n20198 ;
  assign n20363 = n34402 & n20199 ;
  assign n20364 = x29 & n20050 ;
  assign n34403 = ~n20185 ;
  assign n20365 = n34403 & n20364 ;
  assign n34404 = ~n20364 ;
  assign n20366 = n20185 & n34404 ;
  assign n20367 = n20365 | n20366 ;
  assign n20285 = n3791 & n34383 ;
  assign n19978 = n3802 & n34372 ;
  assign n20015 = n209 & n19991 ;
  assign n20368 = n19978 | n20015 ;
  assign n20369 = n3818 & n34381 ;
  assign n20370 = n20368 | n20369 ;
  assign n20371 = n20285 | n20370 ;
  assign n20372 = x26 | n20371 ;
  assign n20373 = x26 & n20371 ;
  assign n34405 = ~n20373 ;
  assign n20374 = n20372 & n34405 ;
  assign n20376 = n20367 | n20374 ;
  assign n20377 = n260 & n34367 ;
  assign n20172 = n3791 & n20170 ;
  assign n20378 = n3818 & n34350 ;
  assign n20379 = n3802 & n34367 ;
  assign n20380 = n20378 | n20379 ;
  assign n20381 = n20172 | n20380 ;
  assign n20382 = n20377 | n20381 ;
  assign n20383 = x26 & n20382 ;
  assign n20004 = n3818 & n19991 ;
  assign n20384 = n3802 & n34350 ;
  assign n20385 = n209 & n34367 ;
  assign n20386 = n20384 | n20385 ;
  assign n20387 = n20004 | n20386 ;
  assign n20388 = n3791 & n20189 ;
  assign n20389 = n20387 | n20388 ;
  assign n20391 = n20383 | n20389 ;
  assign n34406 = ~n20391 ;
  assign n20392 = x26 & n34406 ;
  assign n20394 = n20050 | n20392 ;
  assign n20210 = n3791 & n20207 ;
  assign n20009 = n3802 & n19991 ;
  assign n20028 = n209 & n34350 ;
  assign n20395 = n20009 | n20028 ;
  assign n20396 = n3818 & n34372 ;
  assign n20397 = n20395 | n20396 ;
  assign n20398 = n20210 | n20397 ;
  assign n34407 = ~n20398 ;
  assign n20399 = x26 & n34407 ;
  assign n20400 = n30019 & n20398 ;
  assign n20401 = n20399 | n20400 ;
  assign n20402 = n20394 & n20401 ;
  assign n20375 = n20367 & n20374 ;
  assign n34408 = ~n20375 ;
  assign n20403 = n34408 & n20376 ;
  assign n34409 = ~n20402 ;
  assign n20404 = n34409 & n20403 ;
  assign n34410 = ~n20404 ;
  assign n20405 = n20376 & n34410 ;
  assign n20407 = n20363 | n20405 ;
  assign n34411 = ~n20056 ;
  assign n20291 = n19942 & n34411 ;
  assign n20408 = n34381 & n20127 ;
  assign n20409 = n20291 | n20408 ;
  assign n20410 = n19917 & n20409 ;
  assign n20411 = n19917 | n20409 ;
  assign n34412 = ~n20410 ;
  assign n20412 = n34412 & n20411 ;
  assign n20413 = n3791 & n20412 ;
  assign n19953 = n3802 & n34381 ;
  assign n19980 = n209 & n34372 ;
  assign n20423 = n19953 | n19980 ;
  assign n20424 = n3818 & n19917 ;
  assign n20425 = n20423 | n20424 ;
  assign n20426 = n20413 | n20425 ;
  assign n34413 = ~n20426 ;
  assign n20427 = x26 & n34413 ;
  assign n20428 = n30019 & n20426 ;
  assign n20429 = n20427 | n20428 ;
  assign n20406 = n20363 & n20405 ;
  assign n34414 = ~n20406 ;
  assign n20430 = n34414 & n20407 ;
  assign n34415 = ~n20429 ;
  assign n20431 = n34415 & n20430 ;
  assign n34416 = ~n20431 ;
  assign n20432 = n20407 & n34416 ;
  assign n34417 = ~n20432 ;
  assign n20434 = n20362 & n34417 ;
  assign n34418 = ~n20434 ;
  assign n20435 = n20361 & n34418 ;
  assign n20437 = n20333 | n20435 ;
  assign n34419 = ~n20331 ;
  assign n20438 = n34419 & n20437 ;
  assign n34420 = ~n20271 ;
  assign n20439 = n20229 & n34420 ;
  assign n20440 = n3504 | n4859 ;
  assign n20441 = n11600 | n20440 ;
  assign n20442 = n200 | n560 ;
  assign n20443 = n447 | n20442 ;
  assign n20444 = n1454 | n1626 ;
  assign n20445 = n20443 | n20444 ;
  assign n20446 = n20441 | n20445 ;
  assign n20447 = n12333 | n13886 ;
  assign n20448 = n20446 | n20447 ;
  assign n20449 = n401 | n978 ;
  assign n20450 = n233 | n20449 ;
  assign n20451 = n771 | n1100 ;
  assign n20452 = n20450 | n20451 ;
  assign n34421 = ~n20452 ;
  assign n20453 = n3292 & n34421 ;
  assign n34422 = ~n3760 ;
  assign n20454 = n34422 & n20453 ;
  assign n34423 = ~n20448 ;
  assign n20455 = n34423 & n20454 ;
  assign n20456 = n30449 & n20455 ;
  assign n20457 = n34379 & n20456 ;
  assign n20458 = n20439 & n20457 ;
  assign n20459 = n20439 | n20457 ;
  assign n34424 = ~n20458 ;
  assign n20460 = n34424 & n20459 ;
  assign n20190 = n889 & n20189 ;
  assign n20027 = n3329 & n34350 ;
  assign n20046 = n3311 & n34367 ;
  assign n20461 = n20027 | n20046 ;
  assign n20462 = n3343 & n19991 ;
  assign n20463 = n20461 | n20462 ;
  assign n20464 = n20190 | n20463 ;
  assign n20465 = n20460 | n20464 ;
  assign n20466 = n20460 & n20464 ;
  assign n34425 = ~n20466 ;
  assign n20467 = n20465 & n34425 ;
  assign n20414 = n895 & n20412 ;
  assign n19946 = n2849 & n34381 ;
  assign n19976 = n2861 & n34372 ;
  assign n20468 = n19946 | n19976 ;
  assign n20469 = n894 & n19917 ;
  assign n20470 = n20468 | n20469 ;
  assign n20471 = n20414 | n20470 ;
  assign n34426 = ~n20471 ;
  assign n20472 = x29 & n34426 ;
  assign n20473 = n30024 & n20471 ;
  assign n20474 = n20472 | n20473 ;
  assign n34427 = ~n20474 ;
  assign n20475 = n20467 & n34427 ;
  assign n34428 = ~n20467 ;
  assign n20476 = n34428 & n20474 ;
  assign n20477 = n20475 | n20476 ;
  assign n20303 = n20225 | n20301 ;
  assign n34429 = ~n20300 ;
  assign n20478 = n34429 & n20303 ;
  assign n34430 = ~n20477 ;
  assign n20479 = n34430 & n20478 ;
  assign n34431 = ~n20478 ;
  assign n20480 = n20477 & n34431 ;
  assign n20481 = n20479 | n20480 ;
  assign n34432 = ~n20060 ;
  assign n20061 = n19870 & n34432 ;
  assign n34433 = ~n19870 ;
  assign n20482 = n34433 & n20130 ;
  assign n20483 = n20061 | n20482 ;
  assign n20484 = n19846 & n20483 ;
  assign n20485 = n19846 | n20483 ;
  assign n34434 = ~n20484 ;
  assign n20486 = n34434 & n20485 ;
  assign n20487 = n3791 & n20486 ;
  assign n19879 = n3802 & n19870 ;
  assign n19901 = n209 & n19893 ;
  assign n20498 = n19879 | n19901 ;
  assign n20499 = n3818 & n19846 ;
  assign n20500 = n20498 | n20499 ;
  assign n20501 = n20487 | n20500 ;
  assign n34435 = ~n20501 ;
  assign n20502 = x26 & n34435 ;
  assign n20503 = n30019 & n20501 ;
  assign n20504 = n20502 | n20503 ;
  assign n34436 = ~n20504 ;
  assign n20505 = n20481 & n34436 ;
  assign n34437 = ~n20481 ;
  assign n20506 = n34437 & n20504 ;
  assign n20507 = n20505 | n20506 ;
  assign n34438 = ~n20507 ;
  assign n20508 = n20438 & n34438 ;
  assign n34439 = ~n20438 ;
  assign n20509 = n34439 & n20507 ;
  assign n20510 = n20508 | n20509 ;
  assign n20511 = n20116 | n20135 ;
  assign n34440 = ~n20511 ;
  assign n20512 = n19824 & n34440 ;
  assign n34441 = ~n19824 ;
  assign n20513 = n34441 & n20511 ;
  assign n20514 = n20512 | n20513 ;
  assign n34442 = ~n20514 ;
  assign n20515 = n4135 & n34442 ;
  assign n20079 = n4185 & n20067 ;
  assign n20105 = n4148 & n34354 ;
  assign n20528 = n20079 | n20105 ;
  assign n34443 = ~n18555 ;
  assign n20526 = n34443 & n19634 ;
  assign n20527 = n19635 | n20526 ;
  assign n20529 = n4165 & n20527 ;
  assign n20530 = n20528 | n20529 ;
  assign n20531 = n20515 | n20530 ;
  assign n20532 = x23 | n20531 ;
  assign n20533 = x23 & n20531 ;
  assign n34444 = ~n20533 ;
  assign n20534 = n20532 & n34444 ;
  assign n34445 = ~n20534 ;
  assign n20536 = n20510 & n34445 ;
  assign n20535 = n20510 & n20534 ;
  assign n20537 = n20510 | n20534 ;
  assign n34446 = ~n20535 ;
  assign n20538 = n34446 & n20537 ;
  assign n34447 = ~n20333 ;
  assign n20436 = n34447 & n20435 ;
  assign n34448 = ~n20435 ;
  assign n20539 = n20333 & n34448 ;
  assign n20540 = n20436 | n20539 ;
  assign n20541 = n34345 & n20133 ;
  assign n20542 = n34354 & n20541 ;
  assign n34449 = ~n20541 ;
  assign n20543 = n20093 & n34449 ;
  assign n20544 = n20542 | n20543 ;
  assign n34450 = ~n20544 ;
  assign n20545 = n4135 & n34450 ;
  assign n19857 = n4185 & n19846 ;
  assign n20081 = n4148 & n20067 ;
  assign n20558 = n19857 | n20081 ;
  assign n19633 = n18574 & n19631 ;
  assign n20556 = n18574 | n19631 ;
  assign n34451 = ~n19633 ;
  assign n20557 = n34451 & n20556 ;
  assign n34452 = ~n20557 ;
  assign n20559 = n4165 & n34452 ;
  assign n20560 = n20558 | n20559 ;
  assign n20561 = n20545 | n20560 ;
  assign n20562 = x23 | n20561 ;
  assign n20563 = x23 & n20561 ;
  assign n34453 = ~n20563 ;
  assign n20564 = n20562 & n34453 ;
  assign n34454 = ~n20564 ;
  assign n20566 = n20540 & n34454 ;
  assign n34455 = ~n20540 ;
  assign n20565 = n34455 & n20564 ;
  assign n20567 = n20565 | n20566 ;
  assign n20433 = n20362 & n20432 ;
  assign n20568 = n20362 | n20432 ;
  assign n34456 = ~n20433 ;
  assign n20569 = n34456 & n20568 ;
  assign n34457 = ~n20133 ;
  assign n20134 = n19846 & n34457 ;
  assign n34458 = ~n20130 ;
  assign n20574 = n19846 & n34458 ;
  assign n20575 = n19870 | n20574 ;
  assign n34459 = ~n20575 ;
  assign n20576 = n20067 & n34459 ;
  assign n20577 = n20134 | n20576 ;
  assign n34460 = ~n19846 ;
  assign n20570 = n34460 & n20060 ;
  assign n20571 = n20067 & n20570 ;
  assign n20572 = n20067 | n20570 ;
  assign n34461 = ~n20571 ;
  assign n20573 = n34461 & n20572 ;
  assign n20578 = n19870 & n20573 ;
  assign n20579 = n20577 | n20578 ;
  assign n20580 = n4135 & n20579 ;
  assign n19855 = n4148 & n19846 ;
  assign n19874 = n4185 & n19870 ;
  assign n20591 = n19855 | n19874 ;
  assign n20592 = n4165 & n20067 ;
  assign n20593 = n20591 | n20592 ;
  assign n20594 = n20580 | n20593 ;
  assign n20595 = x23 | n20594 ;
  assign n20596 = x23 & n20594 ;
  assign n34462 = ~n20596 ;
  assign n20597 = n20595 & n34462 ;
  assign n20599 = n20569 | n20597 ;
  assign n20598 = n20569 & n20597 ;
  assign n34463 = ~n20598 ;
  assign n20600 = n34463 & n20599 ;
  assign n34464 = ~n20430 ;
  assign n20601 = n20429 & n34464 ;
  assign n20602 = n20431 | n20601 ;
  assign n20488 = n4135 & n20486 ;
  assign n19876 = n4148 & n19870 ;
  assign n19900 = n4185 & n19893 ;
  assign n20603 = n19876 | n19900 ;
  assign n20604 = n4165 & n19846 ;
  assign n20605 = n20603 | n20604 ;
  assign n20606 = n20488 | n20605 ;
  assign n20607 = x23 | n20606 ;
  assign n20608 = x23 & n20606 ;
  assign n34465 = ~n20608 ;
  assign n20609 = n20607 & n34465 ;
  assign n20611 = n20602 | n20609 ;
  assign n20610 = n20602 & n20609 ;
  assign n34466 = ~n20610 ;
  assign n20612 = n34466 & n20611 ;
  assign n34467 = ~n20403 ;
  assign n20613 = n20402 & n34467 ;
  assign n20614 = n20404 | n20613 ;
  assign n20315 = n4135 & n20311 ;
  assign n19899 = n4148 & n19893 ;
  assign n19922 = n4185 & n19917 ;
  assign n20615 = n19899 | n19922 ;
  assign n20616 = n4165 & n19870 ;
  assign n20617 = n20615 | n20616 ;
  assign n20618 = n20315 | n20617 ;
  assign n20619 = x23 | n20618 ;
  assign n20620 = x23 & n20618 ;
  assign n34468 = ~n20620 ;
  assign n20621 = n20619 & n34468 ;
  assign n20623 = n20614 | n20621 ;
  assign n20622 = n20614 & n20621 ;
  assign n34469 = ~n20622 ;
  assign n20624 = n34469 & n20623 ;
  assign n34470 = ~n20050 ;
  assign n20393 = n34470 & n20392 ;
  assign n34471 = ~n20392 ;
  assign n20625 = n20050 & n34471 ;
  assign n20626 = n20393 | n20625 ;
  assign n34472 = ~n20401 ;
  assign n20627 = n34472 & n20626 ;
  assign n34473 = ~n20626 ;
  assign n20628 = n20401 & n34473 ;
  assign n20629 = n20627 | n20628 ;
  assign n20390 = n20383 & n20389 ;
  assign n34474 = ~n20390 ;
  assign n20630 = n34474 & n20391 ;
  assign n20045 = n4132 & n34367 ;
  assign n20173 = n4135 & n20170 ;
  assign n20631 = n4165 & n34350 ;
  assign n20632 = n4148 & n34367 ;
  assign n20633 = n20631 | n20632 ;
  assign n20634 = n20173 | n20633 ;
  assign n20635 = n20045 | n20634 ;
  assign n20636 = x23 & n20635 ;
  assign n20005 = n4165 & n19991 ;
  assign n20637 = n4148 & n34350 ;
  assign n20638 = n4185 & n34367 ;
  assign n20639 = n20637 | n20638 ;
  assign n20640 = n20005 | n20639 ;
  assign n20641 = n4135 & n20189 ;
  assign n20642 = n20640 | n20641 ;
  assign n20644 = n20636 | n20642 ;
  assign n34475 = ~n20644 ;
  assign n20645 = x23 & n34475 ;
  assign n20647 = n20377 | n20645 ;
  assign n20212 = n4135 & n20207 ;
  assign n20018 = n4148 & n19991 ;
  assign n20030 = n4185 & n34350 ;
  assign n20648 = n20018 | n20030 ;
  assign n20649 = n4165 & n34372 ;
  assign n20650 = n20648 | n20649 ;
  assign n20651 = n20212 | n20650 ;
  assign n34476 = ~n20651 ;
  assign n20652 = x23 & n34476 ;
  assign n20653 = n30030 & n20651 ;
  assign n20654 = n20652 | n20653 ;
  assign n20655 = n20647 & n20654 ;
  assign n20656 = x26 & n20377 ;
  assign n34477 = ~n20381 ;
  assign n20657 = n34477 & n20656 ;
  assign n34478 = ~n20656 ;
  assign n20658 = n20381 & n34478 ;
  assign n20659 = n20657 | n20658 ;
  assign n20660 = n20655 & n20659 ;
  assign n20286 = n4135 & n34383 ;
  assign n19983 = n4148 & n34372 ;
  assign n20007 = n4185 & n19991 ;
  assign n20661 = n19983 | n20007 ;
  assign n20662 = n4165 & n34381 ;
  assign n20663 = n20661 | n20662 ;
  assign n20664 = n20286 | n20663 ;
  assign n34479 = ~n20664 ;
  assign n20665 = x23 & n34479 ;
  assign n20666 = n30030 & n20664 ;
  assign n20667 = n20665 | n20666 ;
  assign n20668 = n20655 | n20659 ;
  assign n34480 = ~n20660 ;
  assign n20669 = n34480 & n20668 ;
  assign n20670 = n20667 & n20669 ;
  assign n20671 = n20660 | n20670 ;
  assign n20672 = n20630 | n20671 ;
  assign n20673 = n20630 & n20671 ;
  assign n34481 = ~n20673 ;
  assign n20674 = n20672 & n34481 ;
  assign n20415 = n4135 & n20412 ;
  assign n19944 = n4148 & n34381 ;
  assign n19975 = n4185 & n34372 ;
  assign n20675 = n19944 | n19975 ;
  assign n20676 = n4165 & n19917 ;
  assign n20677 = n20675 | n20676 ;
  assign n20678 = n20415 | n20677 ;
  assign n34482 = ~n20678 ;
  assign n20679 = x23 & n34482 ;
  assign n20680 = n30030 & n20678 ;
  assign n20681 = n20679 | n20680 ;
  assign n34483 = ~n20681 ;
  assign n20682 = n20674 & n34483 ;
  assign n34484 = ~n20682 ;
  assign n20683 = n20672 & n34484 ;
  assign n20685 = n20629 | n20683 ;
  assign n20344 = n4135 & n34399 ;
  assign n19921 = n4148 & n19917 ;
  assign n19951 = n4185 & n34381 ;
  assign n20686 = n19921 | n19951 ;
  assign n20687 = n4165 & n19893 ;
  assign n20688 = n20686 | n20687 ;
  assign n20689 = n20344 | n20688 ;
  assign n20690 = x23 | n20689 ;
  assign n20691 = x23 & n20689 ;
  assign n34485 = ~n20691 ;
  assign n20692 = n20690 & n34485 ;
  assign n20684 = n20629 & n20683 ;
  assign n34486 = ~n20684 ;
  assign n20693 = n34486 & n20685 ;
  assign n34487 = ~n20692 ;
  assign n20694 = n34487 & n20693 ;
  assign n34488 = ~n20694 ;
  assign n20695 = n20685 & n34488 ;
  assign n34489 = ~n20695 ;
  assign n20697 = n20624 & n34489 ;
  assign n34490 = ~n20697 ;
  assign n20698 = n20623 & n34490 ;
  assign n34491 = ~n20698 ;
  assign n20700 = n20612 & n34491 ;
  assign n34492 = ~n20700 ;
  assign n20701 = n20611 & n34492 ;
  assign n34493 = ~n20701 ;
  assign n20703 = n20600 & n34493 ;
  assign n34494 = ~n20703 ;
  assign n20704 = n20599 & n34494 ;
  assign n20706 = n20567 | n20704 ;
  assign n34495 = ~n20566 ;
  assign n20707 = n34495 & n20706 ;
  assign n20709 = n20538 | n20707 ;
  assign n34496 = ~n20536 ;
  assign n20710 = n34496 & n20709 ;
  assign n20581 = n3791 & n20579 ;
  assign n19852 = n3802 & n19846 ;
  assign n19875 = n209 & n19870 ;
  assign n20711 = n19852 | n19875 ;
  assign n20712 = n3818 & n20067 ;
  assign n20713 = n20711 | n20712 ;
  assign n20714 = n20581 | n20713 ;
  assign n20715 = x26 | n20714 ;
  assign n20716 = x26 & n20714 ;
  assign n34497 = ~n20716 ;
  assign n20717 = n20715 & n34497 ;
  assign n34498 = ~n20457 ;
  assign n20718 = n20439 & n34498 ;
  assign n34499 = ~n20460 ;
  assign n20719 = n34499 & n20464 ;
  assign n20720 = n20718 | n20719 ;
  assign n20721 = n611 | n1010 ;
  assign n20722 = n2985 | n20721 ;
  assign n20723 = n689 | n2224 ;
  assign n20724 = n417 | n1787 ;
  assign n20725 = n696 | n20724 ;
  assign n20726 = n20723 | n20725 ;
  assign n20727 = n20722 | n20726 ;
  assign n20728 = n665 | n2955 ;
  assign n20729 = n3922 | n5598 ;
  assign n20730 = n20728 | n20729 ;
  assign n20731 = n1525 | n20730 ;
  assign n20732 = n20727 | n20731 ;
  assign n20733 = n3169 | n20732 ;
  assign n20734 = n3183 | n20733 ;
  assign n20735 = n1840 | n20734 ;
  assign n20736 = n3664 | n20735 ;
  assign n20737 = n20720 | n20736 ;
  assign n20738 = n20720 & n20736 ;
  assign n34500 = ~n20738 ;
  assign n20739 = n20737 & n34500 ;
  assign n20213 = n889 & n20207 ;
  assign n20002 = n3329 & n19991 ;
  assign n20032 = n3311 & n34350 ;
  assign n20740 = n20002 | n20032 ;
  assign n20741 = n3343 & n34372 ;
  assign n20742 = n20740 | n20741 ;
  assign n20743 = n20213 | n20742 ;
  assign n34501 = ~n20743 ;
  assign n20744 = n20739 & n34501 ;
  assign n34502 = ~n20739 ;
  assign n20745 = n34502 & n20743 ;
  assign n20746 = n20744 | n20745 ;
  assign n20347 = n895 & n34399 ;
  assign n19920 = n2849 & n19917 ;
  assign n19955 = n2861 & n34381 ;
  assign n20747 = n19920 | n19955 ;
  assign n20748 = n894 & n19893 ;
  assign n20749 = n20747 | n20748 ;
  assign n20750 = n20347 | n20749 ;
  assign n20751 = x29 | n20750 ;
  assign n20752 = x29 & n20750 ;
  assign n34503 = ~n20752 ;
  assign n20753 = n20751 & n34503 ;
  assign n20754 = n20746 & n20753 ;
  assign n20755 = n20746 | n20753 ;
  assign n34504 = ~n20754 ;
  assign n20756 = n34504 & n20755 ;
  assign n20757 = n20477 | n20478 ;
  assign n34505 = ~n20475 ;
  assign n20758 = n34505 & n20757 ;
  assign n20759 = n20756 & n20758 ;
  assign n20760 = n20756 | n20758 ;
  assign n34506 = ~n20759 ;
  assign n20761 = n34506 & n20760 ;
  assign n20762 = n20717 & n20761 ;
  assign n20763 = n20717 | n20761 ;
  assign n34507 = ~n20762 ;
  assign n20764 = n34507 & n20763 ;
  assign n20765 = n20438 | n20507 ;
  assign n34508 = ~n20505 ;
  assign n20766 = n34508 & n20765 ;
  assign n20767 = n20764 & n20766 ;
  assign n20768 = n20764 | n20766 ;
  assign n34509 = ~n20767 ;
  assign n20769 = n34509 & n20768 ;
  assign n20117 = n19824 & n20116 ;
  assign n20770 = n34441 & n20135 ;
  assign n20771 = n20117 | n20770 ;
  assign n20772 = n34355 & n20771 ;
  assign n34510 = ~n20771 ;
  assign n20773 = n19800 & n34510 ;
  assign n20774 = n20772 | n20773 ;
  assign n34511 = ~n20774 ;
  assign n20775 = n4135 & n34511 ;
  assign n19835 = n4148 & n19824 ;
  assign n20100 = n4185 & n34354 ;
  assign n20788 = n19835 | n20100 ;
  assign n19639 = n18038 & n19637 ;
  assign n34512 = ~n19639 ;
  assign n20786 = n34512 & n19640 ;
  assign n34513 = ~n20786 ;
  assign n20789 = n4165 & n34513 ;
  assign n20790 = n20788 | n20789 ;
  assign n20791 = n20775 | n20790 ;
  assign n20792 = x23 | n20791 ;
  assign n20793 = x23 & n20791 ;
  assign n34514 = ~n20793 ;
  assign n20794 = n20792 & n34514 ;
  assign n20795 = n20769 & n20794 ;
  assign n20796 = n20769 | n20794 ;
  assign n34515 = ~n20795 ;
  assign n20797 = n34515 & n20796 ;
  assign n20798 = n20710 & n20797 ;
  assign n20799 = n20710 | n20797 ;
  assign n34516 = ~n20798 ;
  assign n20800 = n34516 & n20799 ;
  assign n20139 = n19752 & n20138 ;
  assign n20801 = n19752 | n20121 ;
  assign n34517 = ~n20139 ;
  assign n20802 = n34517 & n20801 ;
  assign n20803 = n19729 | n20802 ;
  assign n20804 = n19729 & n20802 ;
  assign n34518 = ~n20804 ;
  assign n20805 = n20803 & n34518 ;
  assign n20806 = n4686 & n20805 ;
  assign n19767 = n4706 & n19752 ;
  assign n34519 = ~n19776 ;
  assign n19778 = n4726 & n34519 ;
  assign n20817 = n19767 | n19778 ;
  assign n34520 = ~n19729 ;
  assign n20818 = n4748 & n34520 ;
  assign n20819 = n20817 | n20818 ;
  assign n20820 = n20806 | n20819 ;
  assign n20821 = x20 | n20820 ;
  assign n20822 = x20 & n20820 ;
  assign n34521 = ~n20822 ;
  assign n20823 = n20821 & n34521 ;
  assign n34522 = ~n20800 ;
  assign n20824 = n34522 & n20823 ;
  assign n34523 = ~n20823 ;
  assign n20825 = n20800 & n34523 ;
  assign n20826 = n20824 | n20825 ;
  assign n34524 = ~n20538 ;
  assign n20708 = n34524 & n20707 ;
  assign n34525 = ~n20707 ;
  assign n20827 = n20538 & n34525 ;
  assign n20828 = n20708 | n20827 ;
  assign n20120 = n34519 & n20119 ;
  assign n20829 = n19776 & n20137 ;
  assign n20830 = n20120 | n20829 ;
  assign n20831 = n19752 & n20830 ;
  assign n20832 = n19752 | n20830 ;
  assign n34526 = ~n20831 ;
  assign n20833 = n34526 & n20832 ;
  assign n20834 = n4686 & n20833 ;
  assign n19782 = n4706 & n34519 ;
  assign n19809 = n4726 & n34355 ;
  assign n20846 = n19782 | n19809 ;
  assign n34527 = ~n17088 ;
  assign n19645 = n34527 & n19643 ;
  assign n20845 = n19645 | n19646 ;
  assign n20847 = n4748 & n20845 ;
  assign n20848 = n20846 | n20847 ;
  assign n20849 = n20834 | n20848 ;
  assign n20850 = x20 | n20849 ;
  assign n20851 = x20 & n20849 ;
  assign n34528 = ~n20851 ;
  assign n20852 = n20850 & n34528 ;
  assign n34529 = ~n20852 ;
  assign n20854 = n20828 & n34529 ;
  assign n20853 = n20828 & n20852 ;
  assign n20855 = n20828 | n20852 ;
  assign n34530 = ~n20853 ;
  assign n20856 = n34530 & n20855 ;
  assign n34531 = ~n20567 ;
  assign n20705 = n34531 & n20704 ;
  assign n34532 = ~n20704 ;
  assign n20857 = n20567 & n34532 ;
  assign n20858 = n20705 | n20857 ;
  assign n20787 = n20118 & n20786 ;
  assign n20859 = n20136 | n20786 ;
  assign n34533 = ~n20787 ;
  assign n20860 = n34533 & n20859 ;
  assign n20861 = n19776 | n20860 ;
  assign n20862 = n19776 & n20860 ;
  assign n34534 = ~n20862 ;
  assign n20863 = n20861 & n34534 ;
  assign n20864 = n4686 & n20863 ;
  assign n19808 = n4706 & n34355 ;
  assign n19832 = n4726 & n19824 ;
  assign n20877 = n19808 | n19832 ;
  assign n20875 = n17545 & n19641 ;
  assign n34535 = ~n20875 ;
  assign n20876 = n19642 & n34535 ;
  assign n34536 = ~n20876 ;
  assign n20878 = n4748 & n34536 ;
  assign n20879 = n20877 | n20878 ;
  assign n20880 = n20864 | n20879 ;
  assign n20881 = x20 | n20880 ;
  assign n20882 = x20 & n20880 ;
  assign n34537 = ~n20882 ;
  assign n20883 = n20881 & n34537 ;
  assign n34538 = ~n20883 ;
  assign n20885 = n20858 & n34538 ;
  assign n20884 = n20858 & n20883 ;
  assign n20886 = n20858 | n20883 ;
  assign n34539 = ~n20884 ;
  assign n20887 = n34539 & n20886 ;
  assign n20702 = n20600 & n20701 ;
  assign n20888 = n20600 | n20701 ;
  assign n34540 = ~n20702 ;
  assign n20889 = n34540 & n20888 ;
  assign n20777 = n4686 & n34511 ;
  assign n19838 = n4706 & n19824 ;
  assign n20103 = n4726 & n34354 ;
  assign n20890 = n19838 | n20103 ;
  assign n20891 = n4748 & n34513 ;
  assign n20892 = n20890 | n20891 ;
  assign n20893 = n20777 | n20892 ;
  assign n20894 = x20 | n20893 ;
  assign n20895 = x20 & n20893 ;
  assign n34541 = ~n20895 ;
  assign n20896 = n20894 & n34541 ;
  assign n20898 = n20889 | n20896 ;
  assign n34542 = ~n20889 ;
  assign n20897 = n34542 & n20896 ;
  assign n34543 = ~n20896 ;
  assign n20899 = n20889 & n34543 ;
  assign n20900 = n20897 | n20899 ;
  assign n20699 = n20612 & n20698 ;
  assign n20901 = n20612 | n20698 ;
  assign n34544 = ~n20699 ;
  assign n20902 = n34544 & n20901 ;
  assign n20518 = n4686 & n34442 ;
  assign n20078 = n4726 & n20067 ;
  assign n20102 = n4706 & n34354 ;
  assign n20903 = n20078 | n20102 ;
  assign n20904 = n4748 & n20527 ;
  assign n20905 = n20903 | n20904 ;
  assign n20906 = n20518 | n20905 ;
  assign n20907 = x20 | n20906 ;
  assign n20908 = x20 & n20906 ;
  assign n34545 = ~n20908 ;
  assign n20909 = n20907 & n34545 ;
  assign n20911 = n20902 | n20909 ;
  assign n20910 = n20902 & n20909 ;
  assign n34546 = ~n20910 ;
  assign n20912 = n34546 & n20911 ;
  assign n20696 = n20624 & n20695 ;
  assign n20913 = n20624 | n20695 ;
  assign n34547 = ~n20696 ;
  assign n20914 = n34547 & n20913 ;
  assign n20546 = n4686 & n34450 ;
  assign n19851 = n4726 & n19846 ;
  assign n20076 = n4706 & n20067 ;
  assign n20915 = n19851 | n20076 ;
  assign n20916 = n4748 & n34452 ;
  assign n20917 = n20915 | n20916 ;
  assign n20918 = n20546 | n20917 ;
  assign n20919 = x20 | n20918 ;
  assign n20920 = x20 & n20918 ;
  assign n34548 = ~n20920 ;
  assign n20921 = n20919 & n34548 ;
  assign n20923 = n20914 | n20921 ;
  assign n20922 = n20914 & n20921 ;
  assign n34549 = ~n20922 ;
  assign n20924 = n34549 & n20923 ;
  assign n34550 = ~n20693 ;
  assign n20925 = n20692 & n34550 ;
  assign n20926 = n20694 | n20925 ;
  assign n20583 = n4686 & n20579 ;
  assign n19850 = n4706 & n19846 ;
  assign n19873 = n4726 & n19870 ;
  assign n20927 = n19850 | n19873 ;
  assign n20928 = n4748 & n20067 ;
  assign n20929 = n20927 | n20928 ;
  assign n20930 = n20583 | n20929 ;
  assign n20931 = x20 | n20930 ;
  assign n20932 = x20 & n20930 ;
  assign n34551 = ~n20932 ;
  assign n20933 = n20931 & n34551 ;
  assign n20935 = n20926 | n20933 ;
  assign n20934 = n20926 & n20933 ;
  assign n34552 = ~n20934 ;
  assign n20936 = n34552 & n20935 ;
  assign n34553 = ~n20674 ;
  assign n20937 = n34553 & n20681 ;
  assign n20938 = n20682 | n20937 ;
  assign n20489 = n4686 & n20486 ;
  assign n19872 = n4706 & n19870 ;
  assign n19905 = n4726 & n19893 ;
  assign n20939 = n19872 | n19905 ;
  assign n20940 = n4748 & n19846 ;
  assign n20941 = n20939 | n20940 ;
  assign n20942 = n20489 | n20941 ;
  assign n20943 = x20 | n20942 ;
  assign n20944 = x20 & n20942 ;
  assign n34554 = ~n20944 ;
  assign n20945 = n20943 & n34554 ;
  assign n20947 = n20938 | n20945 ;
  assign n34555 = ~n20938 ;
  assign n20946 = n34555 & n20945 ;
  assign n34556 = ~n20945 ;
  assign n20948 = n20938 & n34556 ;
  assign n20949 = n20946 | n20948 ;
  assign n20950 = n20667 | n20669 ;
  assign n34557 = ~n20670 ;
  assign n20951 = n34557 & n20950 ;
  assign n20316 = n4686 & n20311 ;
  assign n19898 = n4706 & n19893 ;
  assign n19919 = n4726 & n19917 ;
  assign n20952 = n19898 | n19919 ;
  assign n20953 = n4748 & n19870 ;
  assign n20954 = n20952 | n20953 ;
  assign n20955 = n20316 | n20954 ;
  assign n20956 = x20 | n20955 ;
  assign n20957 = x20 & n20955 ;
  assign n34558 = ~n20957 ;
  assign n20958 = n20956 & n34558 ;
  assign n20959 = n20951 & n20958 ;
  assign n20960 = n20951 | n20958 ;
  assign n34559 = ~n20959 ;
  assign n20961 = n34559 & n20960 ;
  assign n20349 = n4686 & n34399 ;
  assign n19928 = n4706 & n19917 ;
  assign n19948 = n4726 & n34381 ;
  assign n20962 = n19928 | n19948 ;
  assign n20963 = n4748 & n19893 ;
  assign n20964 = n20962 | n20963 ;
  assign n20965 = n20349 | n20964 ;
  assign n34560 = ~n20965 ;
  assign n20966 = x20 & n34560 ;
  assign n20967 = n30374 & n20965 ;
  assign n20968 = n20966 | n20967 ;
  assign n34561 = ~n20377 ;
  assign n20646 = n34561 & n20645 ;
  assign n34562 = ~n20645 ;
  assign n20969 = n20377 & n34562 ;
  assign n20970 = n20646 | n20969 ;
  assign n34563 = ~n20654 ;
  assign n20971 = n34563 & n20970 ;
  assign n34564 = ~n20970 ;
  assign n20972 = n20654 & n34564 ;
  assign n20973 = n20971 | n20972 ;
  assign n20974 = n20968 | n20973 ;
  assign n20975 = n20968 & n20973 ;
  assign n34565 = ~n20975 ;
  assign n20976 = n20974 & n34565 ;
  assign n20643 = n20636 & n20642 ;
  assign n34566 = ~n20643 ;
  assign n20977 = n34566 & n20644 ;
  assign n20044 = n4683 & n34367 ;
  assign n20174 = n4686 & n20170 ;
  assign n20978 = n4748 & n34350 ;
  assign n20979 = n4706 & n34367 ;
  assign n20980 = n20978 | n20979 ;
  assign n20981 = n20174 | n20980 ;
  assign n20982 = n20044 | n20981 ;
  assign n20983 = x20 & n20982 ;
  assign n20001 = n4748 & n19991 ;
  assign n20984 = n4706 & n34350 ;
  assign n20985 = n4726 & n34367 ;
  assign n20986 = n20984 | n20985 ;
  assign n20987 = n20001 | n20986 ;
  assign n20988 = n4686 & n20189 ;
  assign n20989 = n20987 | n20988 ;
  assign n20991 = n20983 | n20989 ;
  assign n34567 = ~n20991 ;
  assign n20992 = x20 & n34567 ;
  assign n20994 = n20045 | n20992 ;
  assign n20215 = n4686 & n20207 ;
  assign n20006 = n4706 & n19991 ;
  assign n20029 = n4726 & n34350 ;
  assign n20995 = n20006 | n20029 ;
  assign n20996 = n4748 & n34372 ;
  assign n20997 = n20995 | n20996 ;
  assign n20998 = n20215 | n20997 ;
  assign n34568 = ~n20998 ;
  assign n20999 = x20 & n34568 ;
  assign n21000 = n30374 & n20998 ;
  assign n21001 = n20999 | n21000 ;
  assign n21002 = n20994 & n21001 ;
  assign n21003 = x23 & n20045 ;
  assign n34569 = ~n20634 ;
  assign n21004 = n34569 & n21003 ;
  assign n34570 = ~n21003 ;
  assign n21005 = n20634 & n34570 ;
  assign n21006 = n21004 | n21005 ;
  assign n21007 = n21002 & n21006 ;
  assign n20287 = n4686 & n34383 ;
  assign n19971 = n4706 & n34372 ;
  assign n19999 = n4726 & n19991 ;
  assign n21008 = n19971 | n19999 ;
  assign n21009 = n4748 & n34381 ;
  assign n21010 = n21008 | n21009 ;
  assign n21011 = n20287 | n21010 ;
  assign n34571 = ~n21011 ;
  assign n21012 = x20 & n34571 ;
  assign n21013 = n30374 & n21011 ;
  assign n21014 = n21012 | n21013 ;
  assign n21015 = n21002 | n21006 ;
  assign n34572 = ~n21007 ;
  assign n21016 = n34572 & n21015 ;
  assign n21018 = n21014 & n21016 ;
  assign n21019 = n21007 | n21018 ;
  assign n21021 = n20977 | n21019 ;
  assign n34573 = ~n21019 ;
  assign n21020 = n20977 & n34573 ;
  assign n34574 = ~n20977 ;
  assign n21022 = n34574 & n21019 ;
  assign n21023 = n21020 | n21022 ;
  assign n20417 = n4686 & n20412 ;
  assign n19947 = n4706 & n34381 ;
  assign n19973 = n4726 & n34372 ;
  assign n21024 = n19947 | n19973 ;
  assign n21025 = n4748 & n19917 ;
  assign n21026 = n21024 | n21025 ;
  assign n21027 = n20417 | n21026 ;
  assign n34575 = ~n21027 ;
  assign n21028 = x20 & n34575 ;
  assign n21029 = n30374 & n21027 ;
  assign n21030 = n21028 | n21029 ;
  assign n34576 = ~n21030 ;
  assign n21032 = n21023 & n34576 ;
  assign n34577 = ~n21032 ;
  assign n21033 = n21021 & n34577 ;
  assign n34578 = ~n21033 ;
  assign n21035 = n20976 & n34578 ;
  assign n34579 = ~n21035 ;
  assign n21036 = n20974 & n34579 ;
  assign n21038 = n20961 & n21036 ;
  assign n21039 = n20959 | n21038 ;
  assign n34580 = ~n21039 ;
  assign n21040 = n20949 & n34580 ;
  assign n34581 = ~n21040 ;
  assign n21041 = n20947 & n34581 ;
  assign n34582 = ~n21041 ;
  assign n21043 = n20936 & n34582 ;
  assign n34583 = ~n21043 ;
  assign n21044 = n20935 & n34583 ;
  assign n34584 = ~n21044 ;
  assign n21046 = n20924 & n34584 ;
  assign n34585 = ~n21046 ;
  assign n21047 = n20923 & n34585 ;
  assign n34586 = ~n21047 ;
  assign n21049 = n20912 & n34586 ;
  assign n34587 = ~n21049 ;
  assign n21050 = n20911 & n34587 ;
  assign n34588 = ~n21050 ;
  assign n21052 = n20900 & n34588 ;
  assign n34589 = ~n21052 ;
  assign n21053 = n20898 & n34589 ;
  assign n21055 = n20887 | n21053 ;
  assign n34590 = ~n20885 ;
  assign n21056 = n34590 & n21055 ;
  assign n21058 = n20856 | n21056 ;
  assign n34591 = ~n20854 ;
  assign n21059 = n34591 & n21058 ;
  assign n34592 = ~n20826 ;
  assign n21060 = n34592 & n21059 ;
  assign n34593 = ~n21059 ;
  assign n21061 = n20826 & n34593 ;
  assign n21062 = n21060 | n21061 ;
  assign n19651 = n16260 & n19649 ;
  assign n34594 = ~n19651 ;
  assign n21063 = n34594 & n19652 ;
  assign n34595 = ~n20124 ;
  assign n21064 = n34595 & n21063 ;
  assign n34596 = ~n21063 ;
  assign n21065 = n20141 & n34596 ;
  assign n21066 = n21064 | n21065 ;
  assign n21067 = n34349 & n21066 ;
  assign n34597 = ~n21066 ;
  assign n21068 = n19682 & n34597 ;
  assign n21069 = n21067 | n21068 ;
  assign n34598 = ~n21069 ;
  assign n21070 = n37300 & n34598 ;
  assign n19707 = n5144 & n34363 ;
  assign n19736 = n5166 & n34520 ;
  assign n21081 = n19707 | n19736 ;
  assign n21082 = n5191 & n34349 ;
  assign n21083 = n21081 | n21082 ;
  assign n21084 = n21070 | n21083 ;
  assign n21085 = x17 | n21084 ;
  assign n21086 = x17 & n21084 ;
  assign n34599 = ~n21086 ;
  assign n21087 = n21085 & n34599 ;
  assign n34600 = ~n20887 ;
  assign n21054 = n34600 & n21053 ;
  assign n34601 = ~n21053 ;
  assign n21088 = n20887 & n34601 ;
  assign n21089 = n21054 | n21088 ;
  assign n20123 = n34520 & n20122 ;
  assign n21090 = n19729 & n20140 ;
  assign n21091 = n20123 | n21090 ;
  assign n21092 = n34363 & n21091 ;
  assign n34602 = ~n21091 ;
  assign n21093 = n19705 & n34602 ;
  assign n21094 = n21092 | n21093 ;
  assign n34603 = ~n21094 ;
  assign n21095 = n37300 & n34603 ;
  assign n19734 = n5144 & n34520 ;
  assign n19766 = n5166 & n19752 ;
  assign n21106 = n19734 | n19766 ;
  assign n21107 = n5191 & n34596 ;
  assign n21108 = n21106 | n21107 ;
  assign n21109 = n21095 | n21108 ;
  assign n21110 = x17 | n21109 ;
  assign n21111 = x17 & n21109 ;
  assign n34604 = ~n21111 ;
  assign n21112 = n21110 & n34604 ;
  assign n34605 = ~n21112 ;
  assign n21114 = n21089 & n34605 ;
  assign n21113 = n21089 & n21112 ;
  assign n21115 = n21089 | n21112 ;
  assign n34606 = ~n21113 ;
  assign n21116 = n34606 & n21115 ;
  assign n20807 = n37300 & n20805 ;
  assign n19765 = n5144 & n19752 ;
  assign n19784 = n5166 & n34519 ;
  assign n21117 = n19765 | n19784 ;
  assign n21118 = n5191 & n34520 ;
  assign n21119 = n21117 | n21118 ;
  assign n21120 = n20807 | n21119 ;
  assign n21121 = x17 | n21120 ;
  assign n21122 = x17 & n21120 ;
  assign n34607 = ~n21122 ;
  assign n21123 = n21121 & n34607 ;
  assign n21048 = n20912 & n21047 ;
  assign n21124 = n20912 | n21047 ;
  assign n34608 = ~n21048 ;
  assign n21125 = n34608 & n21124 ;
  assign n20835 = n37300 & n20833 ;
  assign n19781 = n5144 & n34519 ;
  assign n19807 = n5166 & n34355 ;
  assign n21126 = n19781 | n19807 ;
  assign n21127 = n5191 & n20845 ;
  assign n21128 = n21126 | n21127 ;
  assign n21129 = n20835 | n21128 ;
  assign n21130 = x17 | n21129 ;
  assign n21131 = x17 & n21129 ;
  assign n34609 = ~n21131 ;
  assign n21132 = n21130 & n34609 ;
  assign n21134 = n21125 | n21132 ;
  assign n34610 = ~n21125 ;
  assign n21133 = n34610 & n21132 ;
  assign n34611 = ~n21132 ;
  assign n21135 = n21125 & n34611 ;
  assign n21136 = n21133 | n21135 ;
  assign n21045 = n20924 & n21044 ;
  assign n21137 = n20924 | n21044 ;
  assign n34612 = ~n21045 ;
  assign n21138 = n34612 & n21137 ;
  assign n20865 = n37300 & n20863 ;
  assign n19812 = n5144 & n34355 ;
  assign n19830 = n5166 & n19824 ;
  assign n21139 = n19812 | n19830 ;
  assign n21140 = n5191 & n34536 ;
  assign n21141 = n21139 | n21140 ;
  assign n21142 = n20865 | n21141 ;
  assign n21143 = x17 | n21142 ;
  assign n21144 = x17 & n21142 ;
  assign n34613 = ~n21144 ;
  assign n21145 = n21143 & n34613 ;
  assign n21147 = n21138 | n21145 ;
  assign n34614 = ~n21138 ;
  assign n21146 = n34614 & n21145 ;
  assign n34615 = ~n21145 ;
  assign n21148 = n21138 & n34615 ;
  assign n21149 = n21146 | n21148 ;
  assign n21042 = n20936 & n21041 ;
  assign n21150 = n20936 | n21041 ;
  assign n34616 = ~n21042 ;
  assign n21151 = n34616 & n21150 ;
  assign n20776 = n37300 & n34511 ;
  assign n19837 = n5144 & n19824 ;
  assign n20098 = n5166 & n34354 ;
  assign n21152 = n19837 | n20098 ;
  assign n21153 = n5191 & n34513 ;
  assign n21154 = n21152 | n21153 ;
  assign n21155 = n20776 | n21154 ;
  assign n21156 = x17 | n21155 ;
  assign n21157 = x17 & n21155 ;
  assign n34617 = ~n21157 ;
  assign n21158 = n21156 & n34617 ;
  assign n21160 = n21151 | n21158 ;
  assign n34618 = ~n21151 ;
  assign n21159 = n34618 & n21158 ;
  assign n34619 = ~n21158 ;
  assign n21161 = n21151 & n34619 ;
  assign n21162 = n21159 | n21161 ;
  assign n34620 = ~n20949 ;
  assign n21163 = n34620 & n21039 ;
  assign n21164 = n21040 | n21163 ;
  assign n20519 = n37300 & n34442 ;
  assign n20073 = n5166 & n20067 ;
  assign n20097 = n5144 & n34354 ;
  assign n21165 = n20073 | n20097 ;
  assign n21166 = n5191 & n20527 ;
  assign n21167 = n21165 | n21166 ;
  assign n21168 = n20519 | n21167 ;
  assign n21169 = x17 | n21168 ;
  assign n21170 = x17 & n21168 ;
  assign n34621 = ~n21170 ;
  assign n21171 = n21169 & n34621 ;
  assign n21173 = n21164 | n21171 ;
  assign n21172 = n21164 & n21171 ;
  assign n34622 = ~n21172 ;
  assign n21174 = n34622 & n21173 ;
  assign n34623 = ~n20961 ;
  assign n21037 = n34623 & n21036 ;
  assign n34624 = ~n21036 ;
  assign n21175 = n20961 & n34624 ;
  assign n21176 = n21037 | n21175 ;
  assign n20548 = n37300 & n34450 ;
  assign n19853 = n5166 & n19846 ;
  assign n20072 = n5144 & n20067 ;
  assign n21177 = n19853 | n20072 ;
  assign n21178 = n5191 & n34452 ;
  assign n21179 = n21177 | n21178 ;
  assign n21180 = n20548 | n21179 ;
  assign n21181 = x17 | n21180 ;
  assign n21182 = x17 & n21180 ;
  assign n34625 = ~n21182 ;
  assign n21183 = n21181 & n34625 ;
  assign n21185 = n21176 | n21183 ;
  assign n21184 = n21176 & n21183 ;
  assign n34626 = ~n21184 ;
  assign n21186 = n34626 & n21185 ;
  assign n21034 = n20976 & n21033 ;
  assign n21187 = n20976 | n21033 ;
  assign n34627 = ~n21034 ;
  assign n21188 = n34627 & n21187 ;
  assign n20586 = n37300 & n20579 ;
  assign n19854 = n5144 & n19846 ;
  assign n19877 = n5166 & n19870 ;
  assign n21189 = n19854 | n19877 ;
  assign n21190 = n5191 & n20067 ;
  assign n21191 = n21189 | n21190 ;
  assign n21192 = n20586 | n21191 ;
  assign n21193 = x17 | n21192 ;
  assign n21194 = x17 & n21192 ;
  assign n34628 = ~n21194 ;
  assign n21195 = n21193 & n34628 ;
  assign n21197 = n21188 | n21195 ;
  assign n21196 = n21188 & n21195 ;
  assign n34629 = ~n21196 ;
  assign n21198 = n34629 & n21197 ;
  assign n21031 = n21023 | n21030 ;
  assign n21199 = n21023 & n21030 ;
  assign n34630 = ~n21199 ;
  assign n21200 = n21031 & n34630 ;
  assign n20490 = n37300 & n20486 ;
  assign n19884 = n5144 & n19870 ;
  assign n19897 = n5166 & n19893 ;
  assign n21201 = n19884 | n19897 ;
  assign n21202 = n5191 & n19846 ;
  assign n21203 = n21201 | n21202 ;
  assign n21204 = n20490 | n21203 ;
  assign n21205 = x17 | n21204 ;
  assign n21206 = x17 & n21204 ;
  assign n34631 = ~n21206 ;
  assign n21207 = n21205 & n34631 ;
  assign n21209 = n21200 | n21207 ;
  assign n34632 = ~n21200 ;
  assign n21208 = n34632 & n21207 ;
  assign n34633 = ~n21207 ;
  assign n21210 = n21200 & n34633 ;
  assign n21211 = n21208 | n21210 ;
  assign n34634 = ~n21014 ;
  assign n21017 = n34634 & n21016 ;
  assign n34635 = ~n21016 ;
  assign n21212 = n21014 & n34635 ;
  assign n21213 = n21017 | n21212 ;
  assign n20313 = n37300 & n20311 ;
  assign n19906 = n5144 & n19893 ;
  assign n19927 = n5166 & n19917 ;
  assign n21214 = n19906 | n19927 ;
  assign n21215 = n5191 & n19870 ;
  assign n21216 = n21214 | n21215 ;
  assign n21217 = n20313 | n21216 ;
  assign n21218 = x17 | n21217 ;
  assign n21219 = x17 & n21217 ;
  assign n34636 = ~n21219 ;
  assign n21220 = n21218 & n34636 ;
  assign n21221 = n21213 & n21220 ;
  assign n34637 = ~n20045 ;
  assign n20993 = n34637 & n20992 ;
  assign n34638 = ~n20992 ;
  assign n21222 = n20045 & n34638 ;
  assign n21223 = n20993 | n21222 ;
  assign n34639 = ~n21001 ;
  assign n21224 = n34639 & n21223 ;
  assign n34640 = ~n21223 ;
  assign n21225 = n21001 & n34640 ;
  assign n21226 = n21224 | n21225 ;
  assign n20990 = n20983 & n20989 ;
  assign n34641 = ~n20990 ;
  assign n21227 = n34641 & n20991 ;
  assign n21228 = x20 & n20044 ;
  assign n34642 = ~n20981 ;
  assign n21229 = n34642 & n21228 ;
  assign n34643 = ~n21228 ;
  assign n21230 = n20981 & n34643 ;
  assign n21231 = n21229 | n21230 ;
  assign n20289 = n37300 & n34383 ;
  assign n19969 = n5144 & n34372 ;
  assign n20008 = n5166 & n19991 ;
  assign n21232 = n19969 | n20008 ;
  assign n21233 = n5191 & n34381 ;
  assign n21234 = n21232 | n21233 ;
  assign n21235 = n20289 | n21234 ;
  assign n21236 = x17 | n21235 ;
  assign n21237 = x17 & n21235 ;
  assign n34644 = ~n21237 ;
  assign n21238 = n21236 & n34644 ;
  assign n21240 = n21231 | n21238 ;
  assign n20042 = n37297 & n34367 ;
  assign n20176 = n37300 & n20170 ;
  assign n21241 = n5191 & n34350 ;
  assign n21242 = n5144 & n34367 ;
  assign n21243 = n21241 | n21242 ;
  assign n21244 = n20176 | n21243 ;
  assign n21245 = n20042 | n21244 ;
  assign n21246 = x17 & n21245 ;
  assign n19998 = n5191 & n19991 ;
  assign n21247 = n5144 & n34350 ;
  assign n21248 = n5166 & n34367 ;
  assign n21249 = n21247 | n21248 ;
  assign n21250 = n19998 | n21249 ;
  assign n21251 = n37300 & n20189 ;
  assign n21252 = n21250 | n21251 ;
  assign n21254 = n21246 | n21252 ;
  assign n34645 = ~n21254 ;
  assign n21255 = x17 & n34645 ;
  assign n21257 = n20044 | n21255 ;
  assign n20216 = n37300 & n20207 ;
  assign n19996 = n5144 & n19991 ;
  assign n20026 = n5166 & n34350 ;
  assign n21258 = n19996 | n20026 ;
  assign n21259 = n5191 & n34372 ;
  assign n21260 = n21258 | n21259 ;
  assign n21261 = n20216 | n21260 ;
  assign n34646 = ~n21261 ;
  assign n21262 = x17 & n34646 ;
  assign n21263 = n30580 & n21261 ;
  assign n21264 = n21262 | n21263 ;
  assign n21265 = n21257 & n21264 ;
  assign n21239 = n21231 & n21238 ;
  assign n34647 = ~n21239 ;
  assign n21266 = n34647 & n21240 ;
  assign n34648 = ~n21265 ;
  assign n21267 = n34648 & n21266 ;
  assign n34649 = ~n21267 ;
  assign n21269 = n21240 & n34649 ;
  assign n21270 = n21227 & n21269 ;
  assign n20418 = n37300 & n20412 ;
  assign n19954 = n5144 & n34381 ;
  assign n19982 = n5166 & n34372 ;
  assign n21271 = n19954 | n19982 ;
  assign n21272 = n5191 & n19917 ;
  assign n21273 = n21271 | n21272 ;
  assign n21274 = n20418 | n21273 ;
  assign n34650 = ~n21274 ;
  assign n21275 = x17 & n34650 ;
  assign n21276 = n30580 & n21274 ;
  assign n21277 = n21275 | n21276 ;
  assign n21278 = n21227 | n21269 ;
  assign n34651 = ~n21270 ;
  assign n21279 = n34651 & n21278 ;
  assign n21281 = n21277 & n21279 ;
  assign n21282 = n21270 | n21281 ;
  assign n21283 = n21226 | n21282 ;
  assign n20348 = n37300 & n34399 ;
  assign n19918 = n5144 & n19917 ;
  assign n19945 = n5166 & n34381 ;
  assign n21284 = n19918 | n19945 ;
  assign n21285 = n5191 & n19893 ;
  assign n21286 = n21284 | n21285 ;
  assign n21287 = n20348 | n21286 ;
  assign n21288 = x17 | n21287 ;
  assign n21289 = x17 & n21287 ;
  assign n34652 = ~n21289 ;
  assign n21290 = n21288 & n34652 ;
  assign n21291 = n21226 & n21282 ;
  assign n34653 = ~n21291 ;
  assign n21292 = n21283 & n34653 ;
  assign n34654 = ~n21290 ;
  assign n21294 = n34654 & n21292 ;
  assign n34655 = ~n21294 ;
  assign n21295 = n21283 & n34655 ;
  assign n21296 = n21213 | n21220 ;
  assign n34656 = ~n21221 ;
  assign n21297 = n34656 & n21296 ;
  assign n21298 = n21295 & n21297 ;
  assign n21299 = n21221 | n21298 ;
  assign n34657 = ~n21299 ;
  assign n21300 = n21211 & n34657 ;
  assign n34658 = ~n21300 ;
  assign n21302 = n21209 & n34658 ;
  assign n34659 = ~n21302 ;
  assign n21304 = n21198 & n34659 ;
  assign n34660 = ~n21304 ;
  assign n21305 = n21197 & n34660 ;
  assign n34661 = ~n21305 ;
  assign n21307 = n21186 & n34661 ;
  assign n34662 = ~n21307 ;
  assign n21308 = n21185 & n34662 ;
  assign n34663 = ~n21308 ;
  assign n21310 = n21174 & n34663 ;
  assign n34664 = ~n21310 ;
  assign n21311 = n21173 & n34664 ;
  assign n34665 = ~n21311 ;
  assign n21313 = n21162 & n34665 ;
  assign n34666 = ~n21313 ;
  assign n21314 = n21160 & n34666 ;
  assign n34667 = ~n21314 ;
  assign n21316 = n21149 & n34667 ;
  assign n34668 = ~n21316 ;
  assign n21317 = n21147 & n34668 ;
  assign n34669 = ~n21317 ;
  assign n21319 = n21136 & n34669 ;
  assign n34670 = ~n21319 ;
  assign n21320 = n21134 & n34670 ;
  assign n21322 = n21123 & n21320 ;
  assign n21051 = n20900 & n21050 ;
  assign n21323 = n20900 | n21050 ;
  assign n34671 = ~n21051 ;
  assign n21324 = n34671 & n21323 ;
  assign n34672 = ~n21320 ;
  assign n21321 = n21123 & n34672 ;
  assign n34673 = ~n21123 ;
  assign n21325 = n34673 & n21320 ;
  assign n21326 = n21321 | n21325 ;
  assign n21327 = n21324 & n21326 ;
  assign n21328 = n21322 | n21327 ;
  assign n21329 = n21116 | n21328 ;
  assign n34674 = ~n21114 ;
  assign n21330 = n34674 & n21329 ;
  assign n21331 = n21087 & n21330 ;
  assign n34675 = ~n20856 ;
  assign n21057 = n34675 & n21056 ;
  assign n34676 = ~n21056 ;
  assign n21332 = n20856 & n34676 ;
  assign n21333 = n21057 | n21332 ;
  assign n21334 = n21087 | n21330 ;
  assign n34677 = ~n21331 ;
  assign n21335 = n34677 & n21334 ;
  assign n34678 = ~n21333 ;
  assign n21336 = n34678 & n21335 ;
  assign n21337 = n21331 | n21336 ;
  assign n21338 = n21062 | n21337 ;
  assign n21339 = n21062 & n21337 ;
  assign n34679 = ~n21339 ;
  assign n21340 = n21338 & n34679 ;
  assign n34680 = ~n20167 ;
  assign n21341 = n34680 & n21340 ;
  assign n34681 = ~n21340 ;
  assign n21342 = n20167 & n34681 ;
  assign n21343 = n21341 | n21342 ;
  assign n13116 = n3791 & n32455 ;
  assign n13070 = n3802 & n32456 ;
  assign n13096 = n209 & n13077 ;
  assign n21344 = n13070 | n13096 ;
  assign n21345 = n3818 & n13027 ;
  assign n21346 = n21344 | n21345 ;
  assign n21347 = n13116 | n21346 ;
  assign n34682 = ~n21347 ;
  assign n21348 = x26 & n34682 ;
  assign n21349 = n30019 & n21347 ;
  assign n21350 = n21348 | n21349 ;
  assign n21351 = n2244 | n2490 ;
  assign n21352 = n4591 | n21351 ;
  assign n21353 = n2937 | n21352 ;
  assign n21354 = n3651 | n21353 ;
  assign n21355 = n508 | n1091 ;
  assign n21356 = n377 | n21355 ;
  assign n21357 = n966 | n21356 ;
  assign n21358 = n2186 | n21357 ;
  assign n21359 = n212 | n704 ;
  assign n21360 = n336 | n21359 ;
  assign n21361 = n956 | n1099 ;
  assign n21362 = n21360 | n21361 ;
  assign n21363 = n11127 | n21362 ;
  assign n21364 = n21358 | n21363 ;
  assign n21365 = n21354 | n21364 ;
  assign n21366 = n1040 | n21365 ;
  assign n21367 = n3458 | n3918 ;
  assign n34683 = ~n21367 ;
  assign n21368 = n5051 & n34683 ;
  assign n34684 = ~n21366 ;
  assign n21369 = n34684 & n21368 ;
  assign n21370 = n15551 & n21369 ;
  assign n21371 = n15551 | n21369 ;
  assign n34685 = ~n21370 ;
  assign n21372 = n34685 & n21371 ;
  assign n21373 = n15355 & n21372 ;
  assign n21374 = n15355 | n21372 ;
  assign n34686 = ~n21373 ;
  assign n21375 = n34686 & n21374 ;
  assign n34687 = ~n15466 ;
  assign n21376 = n34687 & n15469 ;
  assign n21377 = n15465 | n21376 ;
  assign n21378 = n21375 | n21377 ;
  assign n21379 = n21375 & n21377 ;
  assign n34688 = ~n21379 ;
  assign n21380 = n21378 & n34688 ;
  assign n12204 = n889 & n32255 ;
  assign n11861 = n3311 & n32176 ;
  assign n12182 = n3329 & n12161 ;
  assign n21381 = n11861 | n12182 ;
  assign n21382 = n3343 & n32253 ;
  assign n21383 = n21381 | n21382 ;
  assign n21384 = n12204 | n21383 ;
  assign n21385 = n21380 | n21384 ;
  assign n21386 = n21380 & n21384 ;
  assign n34689 = ~n21386 ;
  assign n21387 = n21385 & n34689 ;
  assign n12639 = n895 & n32356 ;
  assign n12581 = n2849 & n12570 ;
  assign n12609 = n2861 & n12595 ;
  assign n21388 = n12581 | n12609 ;
  assign n21389 = n894 & n32354 ;
  assign n21390 = n21388 | n21389 ;
  assign n21391 = n12639 | n21390 ;
  assign n21392 = x29 | n21391 ;
  assign n21393 = x29 & n21391 ;
  assign n34690 = ~n21393 ;
  assign n21394 = n21392 & n34690 ;
  assign n21395 = n15450 | n15479 ;
  assign n34691 = ~n15477 ;
  assign n21396 = n34691 & n21395 ;
  assign n21397 = n21394 & n21396 ;
  assign n21398 = n21394 | n21396 ;
  assign n34692 = ~n21397 ;
  assign n21399 = n34692 & n21398 ;
  assign n34693 = ~n21387 ;
  assign n21400 = n34693 & n21399 ;
  assign n34694 = ~n21399 ;
  assign n21401 = n21387 & n34694 ;
  assign n21402 = n21400 | n21401 ;
  assign n21403 = n21350 | n21402 ;
  assign n21404 = n21350 & n21402 ;
  assign n34695 = ~n21404 ;
  assign n21405 = n21403 & n34695 ;
  assign n34696 = ~n15486 ;
  assign n21406 = n34696 & n15488 ;
  assign n34697 = ~n21405 ;
  assign n21407 = n34697 & n21406 ;
  assign n34698 = ~n21406 ;
  assign n21408 = n21405 & n34698 ;
  assign n21409 = n21407 | n21408 ;
  assign n14190 = n4135 & n14183 ;
  assign n14140 = n4148 & n14124 ;
  assign n14151 = n4185 & n14147 ;
  assign n21410 = n14140 | n14151 ;
  assign n21411 = n4165 & n14196 ;
  assign n21412 = n21410 | n21411 ;
  assign n21413 = n14190 | n21412 ;
  assign n34699 = ~n21413 ;
  assign n21414 = x23 & n34699 ;
  assign n21415 = n30030 & n21413 ;
  assign n21416 = n21414 | n21415 ;
  assign n21417 = n21409 | n21416 ;
  assign n21418 = n21409 & n21416 ;
  assign n34700 = ~n21418 ;
  assign n21419 = n21417 & n34700 ;
  assign n34701 = ~n15490 ;
  assign n21420 = n34701 & n15491 ;
  assign n34702 = ~n15494 ;
  assign n21421 = n15436 & n34702 ;
  assign n21422 = n21420 | n21421 ;
  assign n21423 = n21419 | n21422 ;
  assign n21424 = n21419 & n21422 ;
  assign n34703 = ~n21424 ;
  assign n21425 = n21423 & n34703 ;
  assign n14579 = n4686 & n14570 ;
  assign n14514 = n4706 & n32706 ;
  assign n14540 = n4726 & n14536 ;
  assign n21426 = n14514 | n14540 ;
  assign n21427 = n4748 & n32707 ;
  assign n21428 = n21426 | n21427 ;
  assign n21429 = n14579 | n21428 ;
  assign n34704 = ~n21429 ;
  assign n21430 = x20 & n34704 ;
  assign n21431 = n30374 & n21429 ;
  assign n21432 = n21430 | n21431 ;
  assign n21433 = n21425 | n21432 ;
  assign n21434 = n21425 & n21432 ;
  assign n34705 = ~n21434 ;
  assign n21435 = n21433 & n34705 ;
  assign n34706 = ~n15501 ;
  assign n21436 = n34706 & n15503 ;
  assign n34707 = ~n21435 ;
  assign n21437 = n34707 & n21436 ;
  assign n34708 = ~n21436 ;
  assign n21438 = n21435 & n34708 ;
  assign n21439 = n21437 | n21438 ;
  assign n34709 = ~n15507 ;
  assign n21440 = n15505 & n34709 ;
  assign n34710 = ~n21440 ;
  assign n21441 = n15511 & n34710 ;
  assign n34711 = ~n21441 ;
  assign n21443 = n21439 & n34711 ;
  assign n15192 = n37300 & n32875 ;
  assign n15059 = n5144 & n32856 ;
  assign n15093 = n5166 & n15081 ;
  assign n21444 = n15059 | n15093 ;
  assign n21445 = n5191 & n32876 ;
  assign n21446 = n21444 | n21445 ;
  assign n21447 = n15192 | n21446 ;
  assign n21448 = x17 | n21447 ;
  assign n21449 = x17 & n21447 ;
  assign n34712 = ~n21449 ;
  assign n21450 = n21448 & n34712 ;
  assign n34713 = ~n21439 ;
  assign n21442 = n34713 & n21441 ;
  assign n21451 = n21442 | n21443 ;
  assign n21452 = n21450 | n21451 ;
  assign n34714 = ~n21443 ;
  assign n21454 = n34714 & n21452 ;
  assign n21455 = x14 | n5992 ;
  assign n21456 = n15221 | n21455 ;
  assign n5993 = x14 & n5992 ;
  assign n21457 = x13 | n5932 ;
  assign n34715 = ~n21457 ;
  assign n21458 = n15221 & n34715 ;
  assign n21459 = n5993 | n21458 ;
  assign n34716 = ~n21459 ;
  assign n21460 = n21456 & n34716 ;
  assign n21462 = n21454 | n21460 ;
  assign n21461 = n21454 & n21460 ;
  assign n34717 = ~n21461 ;
  assign n21463 = n34717 & n21462 ;
  assign n15274 = n37300 & n32889 ;
  assign n15060 = n5166 & n32856 ;
  assign n15161 = n5144 & n32876 ;
  assign n21464 = n15060 | n15161 ;
  assign n21465 = n5191 & n32890 ;
  assign n21466 = n21464 | n21465 ;
  assign n21467 = n15274 | n21466 ;
  assign n34718 = ~n21467 ;
  assign n21468 = x17 & n34718 ;
  assign n21469 = n30580 & n21467 ;
  assign n21470 = n21468 | n21469 ;
  assign n15298 = n4686 & n15288 ;
  assign n14507 = n4706 & n32707 ;
  assign n14529 = n4726 & n32706 ;
  assign n21471 = n14507 | n14529 ;
  assign n21472 = n4748 & n15081 ;
  assign n21473 = n21471 | n21472 ;
  assign n21474 = n15298 | n21473 ;
  assign n34719 = ~n21474 ;
  assign n21475 = x20 & n34719 ;
  assign n21476 = n30374 & n21474 ;
  assign n21477 = n21475 | n21476 ;
  assign n34720 = ~n21409 ;
  assign n21478 = n34720 & n21416 ;
  assign n34721 = ~n21419 ;
  assign n21479 = n34721 & n21422 ;
  assign n21480 = n21478 | n21479 ;
  assign n14967 = n4135 & n14965 ;
  assign n14118 = n4148 & n14101 ;
  assign n14141 = n4185 & n14124 ;
  assign n21481 = n14118 | n14141 ;
  assign n21482 = n4165 & n14536 ;
  assign n21483 = n21481 | n21482 ;
  assign n21484 = n14967 | n21483 ;
  assign n34722 = ~n21484 ;
  assign n21485 = x23 & n34722 ;
  assign n21486 = n30030 & n21484 ;
  assign n21487 = n21485 | n21486 ;
  assign n14666 = n3791 & n14655 ;
  assign n13048 = n3802 & n13027 ;
  assign n13072 = n209 & n32456 ;
  assign n21488 = n13048 | n13072 ;
  assign n21489 = n3818 & n14147 ;
  assign n21490 = n21488 | n21489 ;
  assign n21491 = n14666 | n21490 ;
  assign n34723 = ~n21491 ;
  assign n21492 = x26 & n34723 ;
  assign n21493 = n30019 & n21491 ;
  assign n21494 = n21492 | n21493 ;
  assign n14265 = n895 & n32641 ;
  assign n12565 = n2849 & n32354 ;
  assign n12593 = n2861 & n12570 ;
  assign n21495 = n12565 | n12593 ;
  assign n21496 = n894 & n13077 ;
  assign n21497 = n21495 | n21496 ;
  assign n21498 = n14265 | n21497 ;
  assign n34724 = ~n21498 ;
  assign n21499 = x29 & n34724 ;
  assign n21500 = n30024 & n21498 ;
  assign n21501 = n21499 | n21500 ;
  assign n34725 = ~n21375 ;
  assign n21502 = n34725 & n21377 ;
  assign n34726 = ~n21380 ;
  assign n21503 = n34726 & n21384 ;
  assign n21504 = n21502 | n21503 ;
  assign n21505 = n32935 & n21372 ;
  assign n34727 = ~n21505 ;
  assign n21506 = n21371 & n34727 ;
  assign n21507 = n130 | n232 ;
  assign n21508 = n2915 | n21507 ;
  assign n21509 = n212 | n300 ;
  assign n21510 = n560 | n21509 ;
  assign n21511 = n428 | n4859 ;
  assign n21512 = n21510 | n21511 ;
  assign n21513 = n3143 | n3488 ;
  assign n21514 = n290 | n508 ;
  assign n21515 = n3650 | n21514 ;
  assign n21516 = n21513 | n21515 ;
  assign n21517 = n21512 | n21516 ;
  assign n21518 = n364 | n21517 ;
  assign n21519 = n2436 | n21518 ;
  assign n21520 = n4640 | n21519 ;
  assign n21521 = n21508 | n21520 ;
  assign n34728 = ~n21521 ;
  assign n21522 = n21506 & n34728 ;
  assign n34729 = ~n21506 ;
  assign n21523 = n34729 & n21521 ;
  assign n21524 = n21522 | n21523 ;
  assign n13831 = n889 & n32550 ;
  assign n12144 = n3329 & n32253 ;
  assign n12179 = n3311 & n12161 ;
  assign n21525 = n12144 | n12179 ;
  assign n21526 = n3343 & n12595 ;
  assign n21527 = n21525 | n21526 ;
  assign n21528 = n13831 | n21527 ;
  assign n21529 = n21524 | n21528 ;
  assign n21530 = n21524 & n21528 ;
  assign n34730 = ~n21530 ;
  assign n21531 = n21529 & n34730 ;
  assign n21532 = n21504 & n21531 ;
  assign n21533 = n21504 | n21531 ;
  assign n34731 = ~n21532 ;
  assign n21534 = n34731 & n21533 ;
  assign n34732 = ~n21501 ;
  assign n21535 = n34732 & n21534 ;
  assign n34733 = ~n21534 ;
  assign n21536 = n21501 & n34733 ;
  assign n21537 = n21535 | n21536 ;
  assign n21538 = n21397 | n21400 ;
  assign n21539 = n21537 | n21538 ;
  assign n21540 = n21537 & n21538 ;
  assign n34734 = ~n21540 ;
  assign n21541 = n21539 & n34734 ;
  assign n34735 = ~n21494 ;
  assign n21542 = n34735 & n21541 ;
  assign n34736 = ~n21541 ;
  assign n21543 = n21494 & n34736 ;
  assign n21544 = n21542 | n21543 ;
  assign n34737 = ~n21402 ;
  assign n21545 = n21350 & n34737 ;
  assign n21546 = n21407 | n21545 ;
  assign n34738 = ~n21546 ;
  assign n21547 = n21544 & n34738 ;
  assign n34739 = ~n21544 ;
  assign n21548 = n34739 & n21546 ;
  assign n21549 = n21547 | n21548 ;
  assign n34740 = ~n21487 ;
  assign n21550 = n34740 & n21549 ;
  assign n34741 = ~n21549 ;
  assign n21551 = n21487 & n34741 ;
  assign n21552 = n21550 | n21551 ;
  assign n21553 = n21480 | n21552 ;
  assign n21554 = n21480 & n21552 ;
  assign n34742 = ~n21554 ;
  assign n21555 = n21553 & n34742 ;
  assign n34743 = ~n21477 ;
  assign n21556 = n34743 & n21555 ;
  assign n34744 = ~n21555 ;
  assign n21557 = n21477 & n34744 ;
  assign n21558 = n21556 | n21557 ;
  assign n34745 = ~n21425 ;
  assign n21559 = n34745 & n21432 ;
  assign n21560 = n21437 | n21559 ;
  assign n21561 = n21558 | n21560 ;
  assign n21562 = n21558 & n21560 ;
  assign n34746 = ~n21562 ;
  assign n21563 = n21561 & n34746 ;
  assign n34747 = ~n21470 ;
  assign n21564 = n34747 & n21563 ;
  assign n34748 = ~n21563 ;
  assign n21565 = n21470 & n34748 ;
  assign n21566 = n21564 | n21565 ;
  assign n34749 = ~n21566 ;
  assign n21568 = n21463 & n34749 ;
  assign n34750 = ~n21568 ;
  assign n21569 = n21462 & n34750 ;
  assign n15121 = n4686 & n15111 ;
  assign n14508 = n4726 & n32707 ;
  assign n15089 = n4706 & n15081 ;
  assign n21570 = n14508 | n15089 ;
  assign n21571 = n4748 & n32856 ;
  assign n21572 = n21570 | n21571 ;
  assign n21573 = n15121 | n21572 ;
  assign n21574 = x20 | n21573 ;
  assign n21575 = x20 & n21573 ;
  assign n34751 = ~n21575 ;
  assign n21576 = n21574 & n34751 ;
  assign n14689 = n4135 & n32735 ;
  assign n14120 = n4185 & n14101 ;
  assign n14545 = n4148 & n14536 ;
  assign n21577 = n14120 | n14545 ;
  assign n21578 = n4165 & n32706 ;
  assign n21579 = n21577 | n21578 ;
  assign n21580 = n14689 | n21579 ;
  assign n21581 = x23 | n21580 ;
  assign n21582 = x23 & n21580 ;
  assign n34752 = ~n21582 ;
  assign n21583 = n21581 & n34752 ;
  assign n14293 = n3791 & n14283 ;
  assign n13031 = n209 & n13027 ;
  assign n14153 = n3802 & n14147 ;
  assign n21584 = n13031 | n14153 ;
  assign n21585 = n3818 & n14295 ;
  assign n21586 = n21584 | n21585 ;
  assign n21587 = n14293 | n21586 ;
  assign n34753 = ~n21587 ;
  assign n21588 = x26 & n34753 ;
  assign n21589 = n30019 & n21587 ;
  assign n21590 = n21588 | n21589 ;
  assign n21591 = n21506 | n21521 ;
  assign n21592 = n34730 & n21591 ;
  assign n21593 = n713 | n1775 ;
  assign n21594 = n1943 | n21593 ;
  assign n21595 = n1034 | n2347 ;
  assign n21596 = n21594 | n21595 ;
  assign n21597 = n20244 | n21596 ;
  assign n21598 = n2540 | n3525 ;
  assign n21599 = n4658 | n11227 ;
  assign n21600 = n21598 | n21599 ;
  assign n21601 = n3665 | n21600 ;
  assign n21602 = n21597 | n21601 ;
  assign n21603 = n425 | n1949 ;
  assign n21604 = n13408 | n21603 ;
  assign n21605 = n533 | n921 ;
  assign n21606 = n1784 | n21605 ;
  assign n21607 = n107 | n331 ;
  assign n21608 = n476 | n827 ;
  assign n21609 = n21607 | n21608 ;
  assign n21610 = n5854 | n21609 ;
  assign n21611 = n21606 | n21610 ;
  assign n21612 = n12965 | n21611 ;
  assign n21613 = n21604 | n21612 ;
  assign n21614 = n13433 | n21613 ;
  assign n21615 = n21602 | n21614 ;
  assign n21616 = n2001 | n21615 ;
  assign n34754 = ~n21616 ;
  assign n21617 = n21521 & n34754 ;
  assign n21618 = n34728 & n21616 ;
  assign n21619 = n21617 | n21618 ;
  assign n12691 = n889 & n12681 ;
  assign n12157 = n3311 & n32253 ;
  assign n12598 = n3329 & n12595 ;
  assign n21620 = n12157 | n12598 ;
  assign n21621 = n3343 & n12570 ;
  assign n21622 = n21620 | n21621 ;
  assign n21623 = n12691 | n21622 ;
  assign n34755 = ~n21623 ;
  assign n21624 = n21619 & n34755 ;
  assign n34756 = ~n21619 ;
  assign n21626 = n34756 & n21623 ;
  assign n21627 = n21624 | n21626 ;
  assign n21628 = n21592 | n21627 ;
  assign n21629 = n21592 & n21627 ;
  assign n34757 = ~n21629 ;
  assign n21630 = n21628 & n34757 ;
  assign n34758 = ~n21535 ;
  assign n21631 = n21533 & n34758 ;
  assign n21632 = n21630 & n21631 ;
  assign n21633 = n21630 | n21631 ;
  assign n34759 = ~n21632 ;
  assign n21634 = n34759 & n21633 ;
  assign n13858 = n895 & n32557 ;
  assign n12561 = n2861 & n32354 ;
  assign n13097 = n2849 & n13077 ;
  assign n21635 = n12561 | n13097 ;
  assign n21636 = n894 & n32456 ;
  assign n21637 = n21635 | n21636 ;
  assign n21638 = n13858 | n21637 ;
  assign n21639 = x29 | n21638 ;
  assign n21640 = x29 & n21638 ;
  assign n34760 = ~n21640 ;
  assign n21641 = n21639 & n34760 ;
  assign n21642 = n21634 & n21641 ;
  assign n21643 = n21634 | n21641 ;
  assign n34761 = ~n21642 ;
  assign n21644 = n34761 & n21643 ;
  assign n34762 = ~n21590 ;
  assign n21645 = n34762 & n21644 ;
  assign n34763 = ~n21644 ;
  assign n21646 = n21590 & n34763 ;
  assign n21647 = n21645 | n21646 ;
  assign n21648 = n21494 & n21541 ;
  assign n21649 = n21540 | n21648 ;
  assign n21650 = n21647 | n21649 ;
  assign n21651 = n21647 & n21649 ;
  assign n34764 = ~n21651 ;
  assign n21652 = n21650 & n34764 ;
  assign n21653 = n21583 & n21652 ;
  assign n21654 = n21583 | n21652 ;
  assign n34765 = ~n21653 ;
  assign n21655 = n34765 & n21654 ;
  assign n21656 = n21544 | n21546 ;
  assign n34766 = ~n21550 ;
  assign n21657 = n34766 & n21656 ;
  assign n21658 = n21655 & n21657 ;
  assign n21659 = n21655 | n21657 ;
  assign n34767 = ~n21658 ;
  assign n21660 = n34767 & n21659 ;
  assign n21661 = n21576 & n21660 ;
  assign n21662 = n21576 | n21660 ;
  assign n34768 = ~n21661 ;
  assign n21663 = n34768 & n21662 ;
  assign n15533 = n37300 & n15526 ;
  assign n15159 = n5166 & n32876 ;
  assign n15231 = n5191 & n15221 ;
  assign n21664 = n15159 | n15231 ;
  assign n21665 = n5144 & n32890 ;
  assign n21666 = n21664 | n21665 ;
  assign n21667 = n15533 | n21666 ;
  assign n21668 = x17 | n21667 ;
  assign n21669 = x17 & n21667 ;
  assign n34769 = ~n21669 ;
  assign n21670 = n21668 & n34769 ;
  assign n34770 = ~n21556 ;
  assign n21671 = n21553 & n34770 ;
  assign n21672 = n21670 & n21671 ;
  assign n21673 = n21670 | n21671 ;
  assign n34771 = ~n21672 ;
  assign n21674 = n34771 & n21673 ;
  assign n21675 = n21663 & n21674 ;
  assign n21677 = n21663 | n21674 ;
  assign n34772 = ~n21675 ;
  assign n21678 = n34772 & n21677 ;
  assign n34773 = ~n5993 ;
  assign n21679 = n34773 & n21457 ;
  assign n21680 = n21470 & n21563 ;
  assign n21681 = n21562 | n21680 ;
  assign n21682 = n21679 | n21681 ;
  assign n21683 = n21679 & n21681 ;
  assign n34774 = ~n21683 ;
  assign n21684 = n21682 & n34774 ;
  assign n34775 = ~n21678 ;
  assign n21685 = n34775 & n21684 ;
  assign n34776 = ~n21684 ;
  assign n21686 = n21678 & n34776 ;
  assign n21687 = n21685 | n21686 ;
  assign n34777 = ~n21687 ;
  assign n21688 = n21569 & n34777 ;
  assign n34778 = ~n21569 ;
  assign n21689 = n34778 & n21687 ;
  assign n21690 = n21688 | n21689 ;
  assign n21567 = n21463 & n21566 ;
  assign n21691 = n21463 | n21566 ;
  assign n34779 = ~n21567 ;
  assign n21692 = n34779 & n21691 ;
  assign n15523 = n5934 & n15516 ;
  assign n15238 = n5970 & n15221 ;
  assign n21693 = n6018 | n15238 ;
  assign n21694 = n5994 & n32890 ;
  assign n21695 = n21693 | n21694 ;
  assign n21696 = n15523 | n21695 ;
  assign n34780 = ~n21696 ;
  assign n21697 = x14 & n34780 ;
  assign n21698 = n30547 & n21696 ;
  assign n21699 = n21697 | n21698 ;
  assign n34781 = ~n15513 ;
  assign n21700 = n34781 & n15547 ;
  assign n21701 = n15545 | n21700 ;
  assign n21702 = n21699 | n21701 ;
  assign n34782 = ~n21451 ;
  assign n21453 = n21450 & n34782 ;
  assign n34783 = ~n21450 ;
  assign n21703 = n34783 & n21451 ;
  assign n21704 = n21453 | n21703 ;
  assign n21705 = n21699 & n21701 ;
  assign n34784 = ~n21705 ;
  assign n21706 = n21702 & n34784 ;
  assign n21707 = n21704 & n21706 ;
  assign n34785 = ~n21707 ;
  assign n21708 = n21702 & n34785 ;
  assign n21710 = n21692 | n21708 ;
  assign n34786 = ~n21692 ;
  assign n21709 = n34786 & n21708 ;
  assign n34787 = ~n21708 ;
  assign n21711 = n21692 & n34787 ;
  assign n21712 = n21709 | n21711 ;
  assign n21713 = n15550 & n32966 ;
  assign n34788 = ~n21713 ;
  assign n21714 = n15554 & n34788 ;
  assign n21715 = n21704 | n21706 ;
  assign n21716 = n34785 & n21715 ;
  assign n34789 = ~n21714 ;
  assign n21718 = n34789 & n21716 ;
  assign n21717 = n21714 & n21716 ;
  assign n21719 = n21714 | n21716 ;
  assign n34790 = ~n21717 ;
  assign n21720 = n34790 & n21719 ;
  assign n34791 = ~n15559 ;
  assign n21721 = n34791 & n20159 ;
  assign n21722 = n21720 | n21721 ;
  assign n34792 = ~n21718 ;
  assign n21723 = n34792 & n21722 ;
  assign n34793 = ~n21723 ;
  assign n21725 = n21712 & n34793 ;
  assign n34794 = ~n21725 ;
  assign n21726 = n21710 & n34794 ;
  assign n21727 = n21690 & n21726 ;
  assign n21728 = n21690 | n21726 ;
  assign n34795 = ~n21727 ;
  assign n21729 = n34795 & n21728 ;
  assign n21724 = n21712 & n21723 ;
  assign n21752 = n21712 | n21723 ;
  assign n34796 = ~n21724 ;
  assign n21753 = n34796 & n21752 ;
  assign n21754 = n21720 & n21721 ;
  assign n34797 = ~n21754 ;
  assign n21755 = n21722 & n34797 ;
  assign n21777 = n19682 | n20125 ;
  assign n21778 = n19659 & n21777 ;
  assign n21779 = n21755 | n21778 ;
  assign n34798 = ~n21753 ;
  assign n21780 = n34798 & n21779 ;
  assign n21782 = n19682 & n20142 ;
  assign n21784 = n19659 | n21782 ;
  assign n21785 = n21755 & n21784 ;
  assign n34799 = ~n21785 ;
  assign n21786 = n21753 & n34799 ;
  assign n21787 = n21780 | n21786 ;
  assign n34800 = ~n21787 ;
  assign n21788 = n21729 & n34800 ;
  assign n34801 = ~n21729 ;
  assign n21789 = n34801 & n21787 ;
  assign n21790 = n21788 | n21789 ;
  assign n34802 = ~n21790 ;
  assign n21791 = n5937 & n34802 ;
  assign n34803 = ~n21755 ;
  assign n21767 = n5994 & n34803 ;
  assign n21819 = n5970 & n21753 ;
  assign n21828 = n21767 | n21819 ;
  assign n34804 = ~n21726 ;
  assign n21802 = n21690 & n34804 ;
  assign n34805 = ~n21690 ;
  assign n21803 = n34805 & n21726 ;
  assign n21804 = n21802 | n21803 ;
  assign n21829 = n6018 & n21804 ;
  assign n21830 = n21828 | n21829 ;
  assign n21831 = n21791 | n21830 ;
  assign n21832 = x14 | n21831 ;
  assign n21833 = x14 & n21831 ;
  assign n34806 = ~n21833 ;
  assign n21834 = n21832 & n34806 ;
  assign n21835 = n21343 & n21834 ;
  assign n21836 = n21343 | n21834 ;
  assign n34807 = ~n21835 ;
  assign n21837 = n34807 & n21836 ;
  assign n34808 = ~n21335 ;
  assign n21838 = n21333 & n34808 ;
  assign n21839 = n21336 | n21838 ;
  assign n21783 = n34360 & n21782 ;
  assign n34809 = ~n21777 ;
  assign n21840 = n19659 & n34809 ;
  assign n21841 = n21783 | n21840 ;
  assign n34810 = ~n21841 ;
  assign n21843 = n21755 & n34810 ;
  assign n21818 = n21753 & n21778 ;
  assign n21844 = n21753 | n21778 ;
  assign n34811 = ~n21818 ;
  assign n21845 = n34811 & n21844 ;
  assign n21846 = n21843 & n21845 ;
  assign n21847 = n21843 | n21845 ;
  assign n34812 = ~n21846 ;
  assign n21848 = n34812 & n21847 ;
  assign n21849 = n5937 & n21848 ;
  assign n19665 = n5994 & n34360 ;
  assign n21763 = n5970 & n34803 ;
  assign n21859 = n19665 | n21763 ;
  assign n21860 = n6018 & n21753 ;
  assign n21861 = n21859 | n21860 ;
  assign n21862 = n21849 | n21861 ;
  assign n21863 = x14 | n21862 ;
  assign n21864 = x14 & n21862 ;
  assign n34813 = ~n21864 ;
  assign n21865 = n21863 & n34813 ;
  assign n34814 = ~n21839 ;
  assign n21866 = n34814 & n21865 ;
  assign n34815 = ~n21865 ;
  assign n21867 = n21839 & n34815 ;
  assign n21868 = n21866 | n21867 ;
  assign n21869 = n21116 & n21328 ;
  assign n34816 = ~n21869 ;
  assign n21870 = n21329 & n34816 ;
  assign n21842 = n34803 & n21841 ;
  assign n21871 = n21842 | n21843 ;
  assign n34817 = ~n21871 ;
  assign n21872 = n5937 & n34817 ;
  assign n19667 = n5970 & n34360 ;
  assign n19687 = n5994 & n34349 ;
  assign n21883 = n19667 | n19687 ;
  assign n21884 = n6018 & n34803 ;
  assign n21885 = n21883 | n21884 ;
  assign n21886 = n21872 | n21885 ;
  assign n21887 = x14 | n21886 ;
  assign n21888 = x14 & n21886 ;
  assign n34818 = ~n21888 ;
  assign n21889 = n21887 & n34818 ;
  assign n34819 = ~n21889 ;
  assign n21891 = n21870 & n34819 ;
  assign n34820 = ~n21870 ;
  assign n21890 = n34820 & n21889 ;
  assign n21892 = n21890 | n21891 ;
  assign n21893 = n21324 | n21326 ;
  assign n34821 = ~n21327 ;
  assign n21894 = n34821 & n21893 ;
  assign n20151 = n5937 & n34362 ;
  assign n19691 = n5970 & n34349 ;
  assign n19718 = n5994 & n34363 ;
  assign n21895 = n19691 | n19718 ;
  assign n21896 = n6018 & n34365 ;
  assign n21897 = n21895 | n21896 ;
  assign n21898 = n20151 | n21897 ;
  assign n21899 = x14 | n21898 ;
  assign n21900 = x14 & n21898 ;
  assign n34822 = ~n21900 ;
  assign n21901 = n21899 & n34822 ;
  assign n21903 = n21894 | n21901 ;
  assign n21318 = n21136 & n21317 ;
  assign n21904 = n21136 | n21317 ;
  assign n34823 = ~n21318 ;
  assign n21905 = n34823 & n21904 ;
  assign n21072 = n5937 & n34598 ;
  assign n19709 = n5970 & n34363 ;
  assign n19731 = n5994 & n34520 ;
  assign n21906 = n19709 | n19731 ;
  assign n21907 = n6018 & n34349 ;
  assign n21908 = n21906 | n21907 ;
  assign n21909 = n21072 | n21908 ;
  assign n21910 = x14 | n21909 ;
  assign n21911 = x14 & n21909 ;
  assign n34824 = ~n21911 ;
  assign n21912 = n21910 & n34824 ;
  assign n21914 = n21905 | n21912 ;
  assign n21913 = n21905 & n21912 ;
  assign n34825 = ~n21913 ;
  assign n21915 = n34825 & n21914 ;
  assign n21315 = n21149 & n21314 ;
  assign n21916 = n21149 | n21314 ;
  assign n34826 = ~n21315 ;
  assign n21917 = n34826 & n21916 ;
  assign n21097 = n5937 & n34603 ;
  assign n19733 = n5970 & n34520 ;
  assign n19764 = n5994 & n19752 ;
  assign n21918 = n19733 | n19764 ;
  assign n21919 = n6018 & n34596 ;
  assign n21920 = n21918 | n21919 ;
  assign n21921 = n21097 | n21920 ;
  assign n21922 = x14 | n21921 ;
  assign n21923 = x14 & n21921 ;
  assign n34827 = ~n21923 ;
  assign n21924 = n21922 & n34827 ;
  assign n21926 = n21917 | n21924 ;
  assign n34828 = ~n21917 ;
  assign n21925 = n34828 & n21924 ;
  assign n34829 = ~n21924 ;
  assign n21927 = n21917 & n34829 ;
  assign n21928 = n21925 | n21927 ;
  assign n20808 = n5937 & n20805 ;
  assign n19763 = n5970 & n19752 ;
  assign n19788 = n5994 & n34519 ;
  assign n21929 = n19763 | n19788 ;
  assign n21930 = n6018 & n34520 ;
  assign n21931 = n21929 | n21930 ;
  assign n21932 = n20808 | n21931 ;
  assign n34830 = ~n21932 ;
  assign n21933 = x14 & n34830 ;
  assign n21934 = n30547 & n21932 ;
  assign n21935 = n21933 | n21934 ;
  assign n34831 = ~n21162 ;
  assign n21312 = n34831 & n21311 ;
  assign n21936 = n21312 | n21313 ;
  assign n21938 = n21935 & n21936 ;
  assign n21309 = n21174 & n21308 ;
  assign n21939 = n21174 | n21308 ;
  assign n34832 = ~n21309 ;
  assign n21940 = n34832 & n21939 ;
  assign n20836 = n5937 & n20833 ;
  assign n19787 = n5970 & n34519 ;
  assign n19810 = n5994 & n34355 ;
  assign n21941 = n19787 | n19810 ;
  assign n21942 = n6018 & n20845 ;
  assign n21943 = n21941 | n21942 ;
  assign n21944 = n20836 | n21943 ;
  assign n21945 = x14 | n21944 ;
  assign n21946 = x14 & n21944 ;
  assign n34833 = ~n21946 ;
  assign n21947 = n21945 & n34833 ;
  assign n21949 = n21940 | n21947 ;
  assign n34834 = ~n21940 ;
  assign n21948 = n34834 & n21947 ;
  assign n34835 = ~n21947 ;
  assign n21950 = n21940 & n34835 ;
  assign n21951 = n21948 | n21950 ;
  assign n21306 = n21186 & n21305 ;
  assign n21952 = n21186 | n21305 ;
  assign n34836 = ~n21306 ;
  assign n21953 = n34836 & n21952 ;
  assign n20867 = n5937 & n20863 ;
  assign n19813 = n5970 & n34355 ;
  assign n19829 = n5994 & n19824 ;
  assign n21954 = n19813 | n19829 ;
  assign n21955 = n6018 & n34536 ;
  assign n21956 = n21954 | n21955 ;
  assign n21957 = n20867 | n21956 ;
  assign n21958 = x14 | n21957 ;
  assign n21959 = x14 & n21957 ;
  assign n34837 = ~n21959 ;
  assign n21960 = n21958 & n34837 ;
  assign n21962 = n21953 | n21960 ;
  assign n34838 = ~n21953 ;
  assign n21961 = n34838 & n21960 ;
  assign n34839 = ~n21960 ;
  assign n21963 = n21953 & n34839 ;
  assign n21964 = n21961 | n21963 ;
  assign n21303 = n21198 & n21302 ;
  assign n21965 = n21198 | n21302 ;
  assign n34840 = ~n21303 ;
  assign n21966 = n34840 & n21965 ;
  assign n20778 = n5937 & n34511 ;
  assign n19834 = n5970 & n19824 ;
  assign n20096 = n5994 & n34354 ;
  assign n21967 = n19834 | n20096 ;
  assign n21968 = n6018 & n34513 ;
  assign n21969 = n21967 | n21968 ;
  assign n21970 = n20778 | n21969 ;
  assign n21971 = x14 | n21970 ;
  assign n21972 = x14 & n21970 ;
  assign n34841 = ~n21972 ;
  assign n21973 = n21971 & n34841 ;
  assign n21975 = n21966 | n21973 ;
  assign n34842 = ~n21966 ;
  assign n21974 = n34842 & n21973 ;
  assign n34843 = ~n21973 ;
  assign n21976 = n21966 & n34843 ;
  assign n21977 = n21974 | n21976 ;
  assign n21301 = n21211 | n21299 ;
  assign n21978 = n21211 & n21299 ;
  assign n34844 = ~n21978 ;
  assign n21979 = n21301 & n34844 ;
  assign n20520 = n5937 & n34442 ;
  assign n20074 = n5994 & n20067 ;
  assign n20094 = n5970 & n34354 ;
  assign n21980 = n20074 | n20094 ;
  assign n21981 = n6018 & n20527 ;
  assign n21982 = n21980 | n21981 ;
  assign n21983 = n20520 | n21982 ;
  assign n21984 = x14 | n21983 ;
  assign n21985 = x14 & n21983 ;
  assign n34845 = ~n21985 ;
  assign n21986 = n21984 & n34845 ;
  assign n21988 = n21979 | n21986 ;
  assign n21987 = n21979 & n21986 ;
  assign n34846 = ~n21987 ;
  assign n21989 = n34846 & n21988 ;
  assign n21990 = n21295 | n21297 ;
  assign n34847 = ~n21298 ;
  assign n21991 = n34847 & n21990 ;
  assign n20550 = n5937 & n34450 ;
  assign n19848 = n5994 & n19846 ;
  assign n20070 = n5970 & n20067 ;
  assign n21992 = n19848 | n20070 ;
  assign n21993 = n6018 & n34452 ;
  assign n21994 = n21992 | n21993 ;
  assign n21995 = n20550 | n21994 ;
  assign n21996 = x14 | n21995 ;
  assign n21997 = x14 & n21995 ;
  assign n34848 = ~n21997 ;
  assign n21998 = n21996 & n34848 ;
  assign n22000 = n21991 | n21998 ;
  assign n21999 = n21991 & n21998 ;
  assign n34849 = ~n21999 ;
  assign n22001 = n34849 & n22000 ;
  assign n21293 = n21290 & n21292 ;
  assign n22002 = n21290 | n21292 ;
  assign n34850 = ~n21293 ;
  assign n22003 = n34850 & n22002 ;
  assign n20587 = n5937 & n20579 ;
  assign n19847 = n5970 & n19846 ;
  assign n19871 = n5994 & n19870 ;
  assign n22004 = n19847 | n19871 ;
  assign n22005 = n6018 & n20067 ;
  assign n22006 = n22004 | n22005 ;
  assign n22007 = n20587 | n22006 ;
  assign n22008 = x14 | n22007 ;
  assign n22009 = x14 & n22007 ;
  assign n34851 = ~n22009 ;
  assign n22010 = n22008 & n34851 ;
  assign n22012 = n22003 | n22010 ;
  assign n22011 = n22003 & n22010 ;
  assign n34852 = ~n22011 ;
  assign n22013 = n34852 & n22012 ;
  assign n34853 = ~n21277 ;
  assign n21280 = n34853 & n21279 ;
  assign n34854 = ~n21279 ;
  assign n22014 = n21277 & n34854 ;
  assign n22015 = n21280 | n22014 ;
  assign n20491 = n5937 & n20486 ;
  assign n19880 = n5970 & n19870 ;
  assign n19904 = n5994 & n19893 ;
  assign n22016 = n19880 | n19904 ;
  assign n22017 = n6018 & n19846 ;
  assign n22018 = n22016 | n22017 ;
  assign n22019 = n20491 | n22018 ;
  assign n22020 = x14 | n22019 ;
  assign n22021 = x14 & n22019 ;
  assign n34855 = ~n22021 ;
  assign n22022 = n22020 & n34855 ;
  assign n22024 = n22015 | n22022 ;
  assign n21268 = n21265 & n21266 ;
  assign n22025 = n21265 | n21266 ;
  assign n34856 = ~n21268 ;
  assign n22026 = n34856 & n22025 ;
  assign n20317 = n5937 & n20311 ;
  assign n19896 = n5970 & n19893 ;
  assign n19926 = n5994 & n19917 ;
  assign n22027 = n19896 | n19926 ;
  assign n22028 = n6018 & n19870 ;
  assign n22029 = n22027 | n22028 ;
  assign n22030 = n20317 | n22029 ;
  assign n22031 = x14 | n22030 ;
  assign n22032 = x14 & n22030 ;
  assign n34857 = ~n22032 ;
  assign n22033 = n22031 & n34857 ;
  assign n22035 = n22026 | n22033 ;
  assign n22034 = n22026 & n22033 ;
  assign n34858 = ~n22034 ;
  assign n22036 = n34858 & n22035 ;
  assign n34859 = ~n20044 ;
  assign n21256 = n34859 & n21255 ;
  assign n34860 = ~n21255 ;
  assign n22037 = n20044 & n34860 ;
  assign n22038 = n21256 | n22037 ;
  assign n34861 = ~n21264 ;
  assign n22039 = n34861 & n22038 ;
  assign n34862 = ~n22038 ;
  assign n22040 = n21264 & n34862 ;
  assign n22041 = n22039 | n22040 ;
  assign n20345 = n5937 & n34399 ;
  assign n19931 = n5970 & n19917 ;
  assign n19943 = n5994 & n34381 ;
  assign n22042 = n19931 | n19943 ;
  assign n22043 = n6018 & n19893 ;
  assign n22044 = n22042 | n22043 ;
  assign n22045 = n20345 | n22044 ;
  assign n22046 = x14 | n22045 ;
  assign n22047 = x14 & n22045 ;
  assign n34863 = ~n22047 ;
  assign n22048 = n22046 & n34863 ;
  assign n22050 = n22041 | n22048 ;
  assign n22049 = n22041 & n22048 ;
  assign n34864 = ~n22049 ;
  assign n22051 = n34864 & n22050 ;
  assign n21253 = n21246 & n21252 ;
  assign n34865 = ~n21253 ;
  assign n22052 = n34865 & n21254 ;
  assign n20040 = n5934 & n34367 ;
  assign n20177 = n5937 & n20170 ;
  assign n22053 = n6018 & n34350 ;
  assign n22054 = n5970 & n34367 ;
  assign n22055 = n22053 | n22054 ;
  assign n22056 = n20177 | n22055 ;
  assign n22057 = n20040 | n22056 ;
  assign n22058 = x14 & n22057 ;
  assign n20191 = n5937 & n20189 ;
  assign n20025 = n5970 & n34350 ;
  assign n20051 = n5994 & n34367 ;
  assign n22059 = n20025 | n20051 ;
  assign n22060 = n6018 & n19991 ;
  assign n22061 = n22059 | n22060 ;
  assign n22062 = n20191 | n22061 ;
  assign n22064 = n22058 | n22062 ;
  assign n34866 = ~n22064 ;
  assign n22065 = x14 & n34866 ;
  assign n22067 = n20042 | n22065 ;
  assign n20214 = n5937 & n20207 ;
  assign n19995 = n5970 & n19991 ;
  assign n20023 = n5994 & n34350 ;
  assign n22068 = n19995 | n20023 ;
  assign n22069 = n6018 & n34372 ;
  assign n22070 = n22068 | n22069 ;
  assign n22071 = n20214 | n22070 ;
  assign n34867 = ~n22071 ;
  assign n22072 = x14 & n34867 ;
  assign n22073 = n30547 & n22071 ;
  assign n22074 = n22072 | n22073 ;
  assign n22075 = n22067 & n22074 ;
  assign n22076 = x17 & n20042 ;
  assign n34868 = ~n21244 ;
  assign n22077 = n34868 & n22076 ;
  assign n34869 = ~n22076 ;
  assign n22078 = n21244 & n34869 ;
  assign n22079 = n22077 | n22078 ;
  assign n22080 = n22075 & n22079 ;
  assign n20283 = n5937 & n34383 ;
  assign n19985 = n5970 & n34372 ;
  assign n19994 = n5994 & n19991 ;
  assign n22081 = n19985 | n19994 ;
  assign n22082 = n6018 & n34381 ;
  assign n22083 = n22081 | n22082 ;
  assign n22084 = n20283 | n22083 ;
  assign n22085 = x14 | n22084 ;
  assign n22086 = x14 & n22084 ;
  assign n34870 = ~n22086 ;
  assign n22087 = n22085 & n34870 ;
  assign n22088 = n22075 | n22079 ;
  assign n34871 = ~n22080 ;
  assign n22089 = n34871 & n22088 ;
  assign n22090 = n22087 & n22089 ;
  assign n22091 = n22080 | n22090 ;
  assign n22093 = n22052 & n22091 ;
  assign n20419 = n5937 & n20412 ;
  assign n19952 = n5970 & n34381 ;
  assign n19986 = n5994 & n34372 ;
  assign n22094 = n19952 | n19986 ;
  assign n22095 = n6018 & n19917 ;
  assign n22096 = n22094 | n22095 ;
  assign n22097 = n20419 | n22096 ;
  assign n34872 = ~n22097 ;
  assign n22098 = x14 & n34872 ;
  assign n22099 = n30547 & n22097 ;
  assign n22100 = n22098 | n22099 ;
  assign n22092 = n22052 | n22091 ;
  assign n34873 = ~n22093 ;
  assign n22101 = n22092 & n34873 ;
  assign n22102 = n22100 & n22101 ;
  assign n22104 = n22093 | n22102 ;
  assign n34874 = ~n22104 ;
  assign n22106 = n22051 & n34874 ;
  assign n34875 = ~n22106 ;
  assign n22107 = n22050 & n34875 ;
  assign n34876 = ~n22107 ;
  assign n22109 = n22036 & n34876 ;
  assign n34877 = ~n22109 ;
  assign n22110 = n22035 & n34877 ;
  assign n22023 = n22015 & n22022 ;
  assign n34878 = ~n22023 ;
  assign n22111 = n34878 & n22024 ;
  assign n34879 = ~n22110 ;
  assign n22113 = n34879 & n22111 ;
  assign n34880 = ~n22113 ;
  assign n22114 = n22024 & n34880 ;
  assign n34881 = ~n22114 ;
  assign n22116 = n22013 & n34881 ;
  assign n34882 = ~n22116 ;
  assign n22117 = n22012 & n34882 ;
  assign n34883 = ~n22117 ;
  assign n22119 = n22001 & n34883 ;
  assign n34884 = ~n22119 ;
  assign n22120 = n22000 & n34884 ;
  assign n34885 = ~n22120 ;
  assign n22122 = n21989 & n34885 ;
  assign n34886 = ~n22122 ;
  assign n22123 = n21988 & n34886 ;
  assign n34887 = ~n22123 ;
  assign n22125 = n21977 & n34887 ;
  assign n34888 = ~n22125 ;
  assign n22126 = n21975 & n34888 ;
  assign n34889 = ~n22126 ;
  assign n22128 = n21964 & n34889 ;
  assign n34890 = ~n22128 ;
  assign n22129 = n21962 & n34890 ;
  assign n34891 = ~n22129 ;
  assign n22131 = n21951 & n34891 ;
  assign n34892 = ~n22131 ;
  assign n22132 = n21949 & n34892 ;
  assign n21937 = n21935 | n21936 ;
  assign n34893 = ~n21938 ;
  assign n22133 = n21937 & n34893 ;
  assign n22135 = n22132 & n22133 ;
  assign n22136 = n21938 | n22135 ;
  assign n34894 = ~n22136 ;
  assign n22137 = n21928 & n34894 ;
  assign n34895 = ~n22137 ;
  assign n22138 = n21926 & n34895 ;
  assign n34896 = ~n22138 ;
  assign n22140 = n21915 & n34896 ;
  assign n34897 = ~n22140 ;
  assign n22141 = n21914 & n34897 ;
  assign n21902 = n21894 & n21901 ;
  assign n34898 = ~n21902 ;
  assign n22142 = n34898 & n21903 ;
  assign n34899 = ~n22141 ;
  assign n22143 = n34899 & n22142 ;
  assign n34900 = ~n22143 ;
  assign n22144 = n21903 & n34900 ;
  assign n22146 = n21892 | n22144 ;
  assign n34901 = ~n21891 ;
  assign n22147 = n34901 & n22146 ;
  assign n34902 = ~n21868 ;
  assign n22149 = n34902 & n22147 ;
  assign n22150 = n21866 | n22149 ;
  assign n34903 = ~n21837 ;
  assign n22151 = n34903 & n22150 ;
  assign n34904 = ~n22150 ;
  assign n22152 = n21837 & n34904 ;
  assign n22153 = n22151 | n22152 ;
  assign n15122 = n4135 & n15111 ;
  assign n14509 = n4185 & n32707 ;
  assign n15084 = n4148 & n15081 ;
  assign n22154 = n14509 | n15084 ;
  assign n22155 = n4165 & n32856 ;
  assign n22156 = n22154 | n22155 ;
  assign n22157 = n15122 | n22156 ;
  assign n34905 = ~n22157 ;
  assign n22158 = x23 & n34905 ;
  assign n22159 = n30030 & n22157 ;
  assign n22160 = n22158 | n22159 ;
  assign n14691 = n3791 & n32735 ;
  assign n14113 = n209 & n14101 ;
  assign n14552 = n3802 & n14536 ;
  assign n22161 = n14113 | n14552 ;
  assign n22162 = n3818 & n32706 ;
  assign n22163 = n22161 | n22162 ;
  assign n22164 = n14691 | n22163 ;
  assign n22165 = x26 | n22164 ;
  assign n22166 = x26 & n22164 ;
  assign n34906 = ~n22166 ;
  assign n22167 = n22165 & n34906 ;
  assign n14289 = n895 & n14283 ;
  assign n13042 = n2861 & n13027 ;
  assign n14154 = n2849 & n14147 ;
  assign n22168 = n13042 | n14154 ;
  assign n22169 = n894 & n14295 ;
  assign n22170 = n22168 | n22169 ;
  assign n22171 = n14289 | n22170 ;
  assign n22172 = x29 | n22171 ;
  assign n22173 = x29 & n22171 ;
  assign n34907 = ~n22173 ;
  assign n22174 = n22172 & n34907 ;
  assign n22175 = n538 | n540 ;
  assign n22176 = n684 | n22175 ;
  assign n22177 = n11208 | n22176 ;
  assign n22178 = n12725 | n22177 ;
  assign n22179 = n80 | n202 ;
  assign n22180 = n651 | n841 ;
  assign n22181 = n22179 | n22180 ;
  assign n22182 = n239 | n290 ;
  assign n22183 = n22181 | n22182 ;
  assign n22184 = n83 | n400 ;
  assign n22185 = n124 | n22184 ;
  assign n22186 = n250 | n11600 ;
  assign n22187 = n22185 | n22186 ;
  assign n22188 = n4263 | n22187 ;
  assign n22189 = n22183 | n22188 ;
  assign n22190 = n22178 | n22189 ;
  assign n22191 = n11144 | n22190 ;
  assign n22192 = n704 | n2396 ;
  assign n22193 = n22191 | n22192 ;
  assign n22194 = n1115 | n2707 ;
  assign n22195 = n5816 | n22194 ;
  assign n22196 = n174 | n200 ;
  assign n22197 = n978 | n22196 ;
  assign n22198 = n920 | n1136 ;
  assign n22199 = n22197 | n22198 ;
  assign n22200 = n759 | n22199 ;
  assign n22201 = n22195 | n22200 ;
  assign n22202 = n1094 | n1870 ;
  assign n22203 = n412 | n470 ;
  assign n22204 = n1472 | n2411 ;
  assign n22205 = n22203 | n22204 ;
  assign n22206 = n22202 | n22205 ;
  assign n22207 = n378 | n1049 ;
  assign n22208 = n11933 | n22207 ;
  assign n22209 = n649 | n1041 ;
  assign n22210 = n22208 | n22209 ;
  assign n22211 = n3540 | n22210 ;
  assign n22212 = n22206 | n22211 ;
  assign n22213 = n22201 | n22212 ;
  assign n22214 = n2536 | n22213 ;
  assign n22215 = n22193 | n22214 ;
  assign n22216 = n380 | n405 ;
  assign n22217 = n1242 | n22216 ;
  assign n22218 = n3553 | n22217 ;
  assign n34908 = ~n22218 ;
  assign n22219 = n2556 & n34908 ;
  assign n22220 = n418 | n422 ;
  assign n22221 = n996 | n22220 ;
  assign n22222 = n614 | n1243 ;
  assign n22223 = n22221 | n22222 ;
  assign n22224 = n2394 | n2743 ;
  assign n22225 = n22223 | n22224 ;
  assign n22226 = n158 | n314 ;
  assign n22227 = n5378 | n13709 ;
  assign n22228 = n22226 | n22227 ;
  assign n22229 = n1500 | n2110 ;
  assign n22230 = n3031 | n4255 ;
  assign n22231 = n22229 | n22230 ;
  assign n22232 = n22228 | n22231 ;
  assign n22233 = n22225 | n22232 ;
  assign n34909 = ~n22233 ;
  assign n22234 = n22219 & n34909 ;
  assign n34910 = ~n3122 ;
  assign n22235 = n34910 & n22234 ;
  assign n34911 = ~n2293 ;
  assign n22236 = n34911 & n22235 ;
  assign n34912 = ~n12278 ;
  assign n22237 = n34912 & n22236 ;
  assign n34913 = ~n22215 ;
  assign n22238 = n34913 & n22237 ;
  assign n34914 = ~n22237 ;
  assign n22239 = n22215 & n34914 ;
  assign n22240 = n22238 | n22239 ;
  assign n22241 = n810 | n3950 ;
  assign n22242 = n12809 | n22241 ;
  assign n22243 = n312 | n474 ;
  assign n22244 = n250 | n22243 ;
  assign n22245 = n1483 | n22244 ;
  assign n22246 = n13439 | n22245 ;
  assign n22247 = n276 | n302 ;
  assign n22248 = n400 | n22247 ;
  assign n22249 = n11575 | n13725 ;
  assign n22250 = n22248 | n22249 ;
  assign n22251 = n11129 | n11739 ;
  assign n22252 = n22250 | n22251 ;
  assign n22253 = n22246 | n22252 ;
  assign n22254 = n22242 | n22253 ;
  assign n22255 = n600 | n22254 ;
  assign n34915 = ~n22255 ;
  assign n22256 = n1711 & n34915 ;
  assign n34916 = ~n5300 ;
  assign n22257 = n34916 & n22256 ;
  assign n22259 = n21679 | n22257 ;
  assign n22258 = n21679 & n22257 ;
  assign n34917 = ~n22258 ;
  assign n22260 = n34917 & n22259 ;
  assign n22261 = n21521 & n22260 ;
  assign n34918 = ~n22261 ;
  assign n22262 = n22259 & n34918 ;
  assign n22264 = n22215 | n22262 ;
  assign n22263 = n34913 & n22262 ;
  assign n34919 = ~n22262 ;
  assign n22265 = n22215 & n34919 ;
  assign n22266 = n22263 | n22265 ;
  assign n14261 = n889 & n32641 ;
  assign n12566 = n3329 & n32354 ;
  assign n12588 = n3311 & n12570 ;
  assign n22267 = n12566 | n12588 ;
  assign n22268 = n3343 & n13077 ;
  assign n22269 = n22267 | n22268 ;
  assign n22270 = n14261 | n22269 ;
  assign n22272 = n22266 & n22270 ;
  assign n34920 = ~n22272 ;
  assign n22273 = n22264 & n34920 ;
  assign n22274 = n22240 & n22273 ;
  assign n22275 = n22240 | n22273 ;
  assign n34921 = ~n22274 ;
  assign n22276 = n34921 & n22275 ;
  assign n13859 = n889 & n32557 ;
  assign n12564 = n3311 & n32354 ;
  assign n13095 = n3329 & n13077 ;
  assign n22277 = n12564 | n13095 ;
  assign n22278 = n3343 & n32456 ;
  assign n22279 = n22277 | n22278 ;
  assign n22280 = n13859 | n22279 ;
  assign n34922 = ~n22280 ;
  assign n22281 = n22276 & n34922 ;
  assign n34923 = ~n22276 ;
  assign n22282 = n34923 & n22280 ;
  assign n22283 = n22281 | n22282 ;
  assign n34924 = ~n22283 ;
  assign n22284 = n22174 & n34924 ;
  assign n34925 = ~n22174 ;
  assign n22285 = n34925 & n22283 ;
  assign n22286 = n22284 | n22285 ;
  assign n21625 = n21618 | n21623 ;
  assign n34926 = ~n21617 ;
  assign n22287 = n34926 & n21625 ;
  assign n12640 = n889 & n32356 ;
  assign n12573 = n3329 & n12570 ;
  assign n12616 = n3311 & n12595 ;
  assign n22288 = n12573 | n12616 ;
  assign n22289 = n3343 & n32354 ;
  assign n22290 = n22288 | n22289 ;
  assign n22291 = n12640 | n22290 ;
  assign n22293 = n22287 & n22291 ;
  assign n22294 = n21521 | n22260 ;
  assign n22295 = n34918 & n22294 ;
  assign n34927 = ~n22291 ;
  assign n22292 = n22287 & n34927 ;
  assign n34928 = ~n22287 ;
  assign n22296 = n34928 & n22291 ;
  assign n22297 = n22292 | n22296 ;
  assign n22298 = n22295 & n22297 ;
  assign n22299 = n22293 | n22298 ;
  assign n22271 = n22266 | n22270 ;
  assign n22300 = n22271 & n34920 ;
  assign n22302 = n22299 | n22300 ;
  assign n14662 = n895 & n14655 ;
  assign n13032 = n2849 & n13027 ;
  assign n13067 = n2861 & n32456 ;
  assign n22303 = n13032 | n13067 ;
  assign n22304 = n894 & n14147 ;
  assign n22305 = n22303 | n22304 ;
  assign n22306 = n14662 | n22305 ;
  assign n34929 = ~n22306 ;
  assign n22307 = x29 & n34929 ;
  assign n22308 = n30024 & n22306 ;
  assign n22309 = n22307 | n22308 ;
  assign n34930 = ~n22299 ;
  assign n22301 = n34930 & n22300 ;
  assign n34931 = ~n22300 ;
  assign n22310 = n22299 & n34931 ;
  assign n22311 = n22301 | n22310 ;
  assign n34932 = ~n22309 ;
  assign n22312 = n34932 & n22311 ;
  assign n34933 = ~n22312 ;
  assign n22313 = n22302 & n34933 ;
  assign n34934 = ~n22286 ;
  assign n22314 = n34934 & n22313 ;
  assign n34935 = ~n22313 ;
  assign n22315 = n22286 & n34935 ;
  assign n22316 = n22314 | n22315 ;
  assign n34936 = ~n22316 ;
  assign n22317 = n22167 & n34936 ;
  assign n34937 = ~n22167 ;
  assign n22318 = n34937 & n22316 ;
  assign n22319 = n22317 | n22318 ;
  assign n34938 = ~n22311 ;
  assign n22320 = n22309 & n34938 ;
  assign n22321 = n22312 | n22320 ;
  assign n13121 = n895 & n32455 ;
  assign n13073 = n2849 & n32456 ;
  assign n13087 = n2861 & n13077 ;
  assign n22322 = n13073 | n13087 ;
  assign n22323 = n894 & n13027 ;
  assign n22324 = n22322 | n22323 ;
  assign n22325 = n13121 | n22324 ;
  assign n34939 = ~n22325 ;
  assign n22326 = x29 & n34939 ;
  assign n22327 = n30024 & n22325 ;
  assign n22328 = n22326 | n22327 ;
  assign n22329 = n22295 | n22297 ;
  assign n34940 = ~n22298 ;
  assign n22330 = n34940 & n22329 ;
  assign n22332 = n22328 | n22330 ;
  assign n34941 = ~n22328 ;
  assign n22331 = n34941 & n22330 ;
  assign n34942 = ~n22330 ;
  assign n22333 = n22328 & n34942 ;
  assign n22334 = n22331 | n22333 ;
  assign n34943 = ~n21631 ;
  assign n22335 = n21630 & n34943 ;
  assign n22336 = n21629 | n22335 ;
  assign n22338 = n22334 & n22336 ;
  assign n34944 = ~n22338 ;
  assign n22339 = n22332 & n34944 ;
  assign n22341 = n22321 | n22339 ;
  assign n14974 = n3791 & n14965 ;
  assign n14116 = n3802 & n14101 ;
  assign n14143 = n209 & n14124 ;
  assign n22342 = n14116 | n14143 ;
  assign n22343 = n3818 & n14536 ;
  assign n22344 = n22342 | n22343 ;
  assign n22345 = n14974 | n22344 ;
  assign n34945 = ~n22345 ;
  assign n22346 = x26 & n34945 ;
  assign n22347 = n30019 & n22345 ;
  assign n22348 = n22346 | n22347 ;
  assign n34946 = ~n22321 ;
  assign n22340 = n34946 & n22339 ;
  assign n34947 = ~n22339 ;
  assign n22349 = n22321 & n34947 ;
  assign n22350 = n22340 | n22349 ;
  assign n34948 = ~n22348 ;
  assign n22351 = n34948 & n22350 ;
  assign n34949 = ~n22351 ;
  assign n22352 = n22341 & n34949 ;
  assign n34950 = ~n22319 ;
  assign n22353 = n34950 & n22352 ;
  assign n34951 = ~n22352 ;
  assign n22354 = n22319 & n34951 ;
  assign n22355 = n22353 | n22354 ;
  assign n22356 = n22160 | n22355 ;
  assign n22357 = n22160 & n22355 ;
  assign n34952 = ~n22357 ;
  assign n22358 = n22356 & n34952 ;
  assign n15534 = n4686 & n15526 ;
  assign n15167 = n4726 & n32876 ;
  assign n15239 = n4748 & n15221 ;
  assign n22359 = n15167 | n15239 ;
  assign n22360 = n4706 & n32890 ;
  assign n22361 = n22359 | n22360 ;
  assign n22362 = n15534 | n22361 ;
  assign n22363 = x20 | n22362 ;
  assign n22364 = x20 & n22362 ;
  assign n34953 = ~n22364 ;
  assign n22365 = n22363 & n34953 ;
  assign n34954 = ~n22350 ;
  assign n22366 = n22348 & n34954 ;
  assign n22367 = n22351 | n22366 ;
  assign n34955 = ~n22336 ;
  assign n22337 = n22334 & n34955 ;
  assign n34956 = ~n22334 ;
  assign n22368 = n34956 & n22336 ;
  assign n22369 = n22337 | n22368 ;
  assign n14193 = n3791 & n14183 ;
  assign n14139 = n3802 & n14124 ;
  assign n14167 = n209 & n14147 ;
  assign n22370 = n14139 | n14167 ;
  assign n22371 = n3818 & n14196 ;
  assign n22372 = n22370 | n22371 ;
  assign n22373 = n14193 | n22372 ;
  assign n34957 = ~n22373 ;
  assign n22374 = x26 & n34957 ;
  assign n22375 = n30019 & n22373 ;
  assign n22376 = n22374 | n22375 ;
  assign n34958 = ~n22369 ;
  assign n22378 = n34958 & n22376 ;
  assign n34959 = ~n22376 ;
  assign n22377 = n22369 & n34959 ;
  assign n22379 = n22377 | n22378 ;
  assign n34960 = ~n21645 ;
  assign n22380 = n21643 & n34960 ;
  assign n34961 = ~n22379 ;
  assign n22381 = n34961 & n22380 ;
  assign n22382 = n22378 | n22381 ;
  assign n22383 = n22367 | n22382 ;
  assign n15296 = n4135 & n15288 ;
  assign n14496 = n4148 & n32707 ;
  assign n14518 = n4185 & n32706 ;
  assign n22384 = n14496 | n14518 ;
  assign n22385 = n4165 & n15081 ;
  assign n22386 = n22384 | n22385 ;
  assign n22387 = n15296 | n22386 ;
  assign n34962 = ~n22387 ;
  assign n22388 = x23 & n34962 ;
  assign n22389 = n30030 & n22387 ;
  assign n22390 = n22388 | n22389 ;
  assign n22391 = n22367 & n22382 ;
  assign n34963 = ~n22391 ;
  assign n22392 = n22383 & n34963 ;
  assign n34964 = ~n22390 ;
  assign n22393 = n34964 & n22392 ;
  assign n34965 = ~n22393 ;
  assign n22394 = n22383 & n34965 ;
  assign n22395 = n22365 & n22394 ;
  assign n22396 = n22365 | n22394 ;
  assign n34966 = ~n22395 ;
  assign n22397 = n34966 & n22396 ;
  assign n22398 = n22358 & n22397 ;
  assign n22399 = n22358 | n22397 ;
  assign n34967 = ~n22398 ;
  assign n22400 = n34967 & n22399 ;
  assign n37296 = x16 | n37294 ;
  assign n5165 = x17 & n5164 ;
  assign n34968 = ~n5165 ;
  assign n22401 = n37296 & n34968 ;
  assign n34969 = ~n22392 ;
  assign n22403 = n22390 & n34969 ;
  assign n22404 = n22393 | n22403 ;
  assign n34970 = ~n22380 ;
  assign n22405 = n22379 & n34970 ;
  assign n22406 = n22381 | n22405 ;
  assign n14581 = n4135 & n14570 ;
  assign n14530 = n4148 & n32706 ;
  assign n14553 = n4185 & n14536 ;
  assign n22407 = n14530 | n14553 ;
  assign n22408 = n4165 & n32707 ;
  assign n22409 = n22407 | n22408 ;
  assign n22410 = n14581 | n22409 ;
  assign n34971 = ~n22410 ;
  assign n22411 = x23 & n34971 ;
  assign n22412 = n30030 & n22410 ;
  assign n22413 = n22411 | n22412 ;
  assign n34972 = ~n22413 ;
  assign n22415 = n22406 & n34972 ;
  assign n22414 = n22406 | n22413 ;
  assign n22416 = n22406 & n22413 ;
  assign n34973 = ~n22416 ;
  assign n22417 = n22414 & n34973 ;
  assign n34974 = ~n21583 ;
  assign n22418 = n34974 & n21652 ;
  assign n34975 = ~n22418 ;
  assign n22419 = n21650 & n34975 ;
  assign n22421 = n22417 | n22419 ;
  assign n34976 = ~n22415 ;
  assign n22422 = n34976 & n22421 ;
  assign n22424 = n22404 & n22422 ;
  assign n34977 = ~n22404 ;
  assign n22423 = n34977 & n22422 ;
  assign n34978 = ~n22422 ;
  assign n22425 = n22404 & n34978 ;
  assign n22426 = n22423 | n22425 ;
  assign n15273 = n4686 & n32889 ;
  assign n15071 = n4726 & n32856 ;
  assign n15168 = n4706 & n32876 ;
  assign n22427 = n15071 | n15168 ;
  assign n22428 = n4748 & n32890 ;
  assign n22429 = n22427 | n22428 ;
  assign n22430 = n15273 | n22429 ;
  assign n34979 = ~n22430 ;
  assign n22431 = x20 & n34979 ;
  assign n22432 = n30374 & n22430 ;
  assign n22433 = n22431 | n22432 ;
  assign n22435 = n22426 & n22433 ;
  assign n22436 = n22424 | n22435 ;
  assign n22437 = n22401 | n22436 ;
  assign n22438 = n22401 & n22436 ;
  assign n34980 = ~n22438 ;
  assign n22439 = n22437 & n34980 ;
  assign n22440 = n22400 & n22439 ;
  assign n22441 = n22400 | n22439 ;
  assign n34981 = ~n22440 ;
  assign n22442 = n34981 & n22441 ;
  assign n34982 = ~n22417 ;
  assign n22420 = n34982 & n22419 ;
  assign n34983 = ~n22419 ;
  assign n22443 = n22417 & n34983 ;
  assign n22444 = n22420 | n22443 ;
  assign n22445 = n21658 | n21661 ;
  assign n34984 = ~n22444 ;
  assign n22454 = n34984 & n22445 ;
  assign n15193 = n4686 & n32875 ;
  assign n15072 = n4706 & n32856 ;
  assign n15088 = n4726 & n15081 ;
  assign n22447 = n15072 | n15088 ;
  assign n22448 = n4748 & n32876 ;
  assign n22449 = n22447 | n22448 ;
  assign n22450 = n15193 | n22449 ;
  assign n34985 = ~n22450 ;
  assign n22451 = x20 & n34985 ;
  assign n22452 = n30374 & n22450 ;
  assign n22453 = n22451 | n22452 ;
  assign n34986 = ~n22445 ;
  assign n22446 = n22444 & n34986 ;
  assign n22455 = n22446 | n22454 ;
  assign n34987 = ~n22455 ;
  assign n22457 = n22453 & n34987 ;
  assign n22458 = n22454 | n22457 ;
  assign n15234 = x17 & n32883 ;
  assign n22459 = n5164 | n15234 ;
  assign n22460 = x16 & n15221 ;
  assign n22461 = n22459 | n22460 ;
  assign n22462 = n34968 & n22461 ;
  assign n22464 = n22458 | n22462 ;
  assign n34988 = ~n22433 ;
  assign n22434 = n22426 & n34988 ;
  assign n34989 = ~n22426 ;
  assign n22465 = n34989 & n22433 ;
  assign n22466 = n22434 | n22465 ;
  assign n22463 = n22458 & n22462 ;
  assign n34990 = ~n22463 ;
  assign n22467 = n34990 & n22464 ;
  assign n34991 = ~n22466 ;
  assign n22468 = n34991 & n22467 ;
  assign n34992 = ~n22468 ;
  assign n22469 = n22464 & n34992 ;
  assign n22470 = n22442 & n22469 ;
  assign n22471 = n22442 | n22469 ;
  assign n34993 = ~n22470 ;
  assign n22472 = n34993 & n22471 ;
  assign n34994 = ~n22467 ;
  assign n22473 = n22466 & n34994 ;
  assign n22474 = n22468 | n22473 ;
  assign n15524 = n37297 & n15516 ;
  assign n15240 = n5144 & n15221 ;
  assign n22475 = n5191 | n15240 ;
  assign n22476 = n5166 & n32890 ;
  assign n22477 = n22475 | n22476 ;
  assign n22478 = n15524 | n22477 ;
  assign n22479 = x17 | n22478 ;
  assign n22480 = x17 & n22478 ;
  assign n34995 = ~n22480 ;
  assign n22481 = n22479 & n34995 ;
  assign n34996 = ~n21663 ;
  assign n21676 = n34996 & n21674 ;
  assign n34997 = ~n21676 ;
  assign n22482 = n21673 & n34997 ;
  assign n22483 = n22481 & n22482 ;
  assign n22456 = n22453 | n22455 ;
  assign n22484 = n22453 & n22455 ;
  assign n34998 = ~n22484 ;
  assign n22485 = n22456 & n34998 ;
  assign n22486 = n22481 | n22482 ;
  assign n34999 = ~n22483 ;
  assign n22487 = n34999 & n22486 ;
  assign n35000 = ~n22485 ;
  assign n22488 = n35000 & n22487 ;
  assign n22489 = n22483 | n22488 ;
  assign n22490 = n22474 | n22489 ;
  assign n22491 = n22474 & n22489 ;
  assign n35001 = ~n22491 ;
  assign n22492 = n22490 & n35001 ;
  assign n35002 = ~n22487 ;
  assign n22493 = n22485 & n35002 ;
  assign n22494 = n22488 | n22493 ;
  assign n35003 = ~n21685 ;
  assign n22495 = n21682 & n35003 ;
  assign n35004 = ~n22495 ;
  assign n22497 = n22494 & n35004 ;
  assign n35005 = ~n22494 ;
  assign n22496 = n35005 & n22495 ;
  assign n22498 = n22496 | n22497 ;
  assign n22499 = n21569 | n21687 ;
  assign n35006 = ~n21802 ;
  assign n22500 = n35006 & n22499 ;
  assign n22502 = n22498 | n22500 ;
  assign n35007 = ~n22497 ;
  assign n22503 = n35007 & n22502 ;
  assign n35008 = ~n22503 ;
  assign n22505 = n22492 & n35008 ;
  assign n35009 = ~n22505 ;
  assign n22506 = n22490 & n35009 ;
  assign n35010 = ~n22472 ;
  assign n22507 = n35010 & n22506 ;
  assign n35011 = ~n22506 ;
  assign n22508 = n22472 & n35011 ;
  assign n22509 = n22507 | n22508 ;
  assign n22504 = n22492 & n22503 ;
  assign n22532 = n22492 | n22503 ;
  assign n35012 = ~n22504 ;
  assign n22533 = n35012 & n22532 ;
  assign n35013 = ~n22498 ;
  assign n22501 = n35013 & n22500 ;
  assign n35014 = ~n22500 ;
  assign n22534 = n22498 & n35014 ;
  assign n22535 = n22501 | n22534 ;
  assign n35015 = ~n21780 ;
  assign n22557 = n21729 & n35015 ;
  assign n35016 = ~n22557 ;
  assign n22558 = n22535 & n35016 ;
  assign n35017 = ~n22558 ;
  assign n22559 = n22533 & n35017 ;
  assign n22560 = n21729 | n21786 ;
  assign n35018 = ~n22535 ;
  assign n22561 = n35018 & n22560 ;
  assign n22562 = n22533 | n22561 ;
  assign n35019 = ~n22559 ;
  assign n22563 = n35019 & n22562 ;
  assign n35020 = ~n22509 ;
  assign n22564 = n35020 & n22563 ;
  assign n35021 = ~n22563 ;
  assign n22565 = n22509 & n35021 ;
  assign n22566 = n22564 | n22565 ;
  assign n35022 = ~n22566 ;
  assign n22567 = n6272 & n35022 ;
  assign n22537 = n6244 & n35018 ;
  assign n22591 = n6190 & n22533 ;
  assign n22601 = n22537 | n22591 ;
  assign n22602 = n6217 & n35020 ;
  assign n22603 = n22601 | n22602 ;
  assign n22604 = n22567 | n22603 ;
  assign n22605 = x11 | n22604 ;
  assign n22606 = x11 & n22604 ;
  assign n35023 = ~n22606 ;
  assign n22607 = n22605 & n35023 ;
  assign n22608 = n22153 & n22607 ;
  assign n22609 = n22153 | n22607 ;
  assign n35024 = ~n22608 ;
  assign n22610 = n35024 & n22609 ;
  assign n22148 = n21868 & n22147 ;
  assign n22611 = n21868 | n22147 ;
  assign n35025 = ~n22148 ;
  assign n22612 = n35025 & n22611 ;
  assign n21781 = n21729 & n21780 ;
  assign n22613 = n34801 & n21786 ;
  assign n22614 = n21781 | n22613 ;
  assign n35026 = ~n22614 ;
  assign n22616 = n22535 & n35026 ;
  assign n35027 = ~n22560 ;
  assign n22588 = n22533 & n35027 ;
  assign n35028 = ~n22533 ;
  assign n22617 = n35028 & n22560 ;
  assign n22618 = n22588 | n22617 ;
  assign n22619 = n22616 | n22618 ;
  assign n22620 = n22616 & n22618 ;
  assign n35029 = ~n22620 ;
  assign n22621 = n22619 & n35029 ;
  assign n35030 = ~n22621 ;
  assign n22622 = n6272 & n35030 ;
  assign n21739 = n6244 & n21729 ;
  assign n22546 = n6190 & n35018 ;
  assign n22632 = n21739 | n22546 ;
  assign n22633 = n6217 & n22533 ;
  assign n22634 = n22632 | n22633 ;
  assign n22635 = n22622 | n22634 ;
  assign n22636 = x11 | n22635 ;
  assign n22637 = x11 & n22635 ;
  assign n35031 = ~n22637 ;
  assign n22638 = n22636 & n35031 ;
  assign n35032 = ~n22638 ;
  assign n22640 = n22612 & n35032 ;
  assign n35033 = ~n21892 ;
  assign n22145 = n35033 & n22144 ;
  assign n35034 = ~n22144 ;
  assign n22641 = n21892 & n35034 ;
  assign n22642 = n22145 | n22641 ;
  assign n22615 = n35018 & n22614 ;
  assign n22643 = n22615 | n22616 ;
  assign n35035 = ~n22643 ;
  assign n22644 = n6272 & n35035 ;
  assign n21741 = n6190 & n21729 ;
  assign n21808 = n6244 & n21753 ;
  assign n22655 = n21741 | n21808 ;
  assign n22656 = n6217 & n35018 ;
  assign n22657 = n22655 | n22656 ;
  assign n22658 = n22644 | n22657 ;
  assign n22659 = x11 | n22658 ;
  assign n22660 = x11 & n22658 ;
  assign n35036 = ~n22660 ;
  assign n22661 = n22659 & n35036 ;
  assign n35037 = ~n22661 ;
  assign n22663 = n22642 & n35037 ;
  assign n35038 = ~n22642 ;
  assign n22662 = n35038 & n22661 ;
  assign n22664 = n22662 | n22663 ;
  assign n21792 = n6272 & n34802 ;
  assign n21765 = n6244 & n34803 ;
  assign n21813 = n6190 & n21753 ;
  assign n22665 = n21765 | n21813 ;
  assign n22666 = n6217 & n21804 ;
  assign n22667 = n22665 | n22666 ;
  assign n22668 = n21792 | n22667 ;
  assign n22669 = x11 | n22668 ;
  assign n22670 = x11 & n22668 ;
  assign n35039 = ~n22670 ;
  assign n22671 = n22669 & n35039 ;
  assign n35040 = ~n22142 ;
  assign n22672 = n22141 & n35040 ;
  assign n22673 = n22143 | n22672 ;
  assign n22675 = n22671 | n22673 ;
  assign n35041 = ~n22673 ;
  assign n22674 = n22671 & n35041 ;
  assign n35042 = ~n22671 ;
  assign n22676 = n35042 & n22673 ;
  assign n22677 = n22674 | n22676 ;
  assign n22139 = n21915 & n22138 ;
  assign n22678 = n21915 | n22138 ;
  assign n35043 = ~n22139 ;
  assign n22679 = n35043 & n22678 ;
  assign n21850 = n6272 & n21848 ;
  assign n19666 = n6244 & n34360 ;
  assign n21761 = n6190 & n34803 ;
  assign n22680 = n19666 | n21761 ;
  assign n22681 = n6217 & n21753 ;
  assign n22682 = n22680 | n22681 ;
  assign n22683 = n21850 | n22682 ;
  assign n22684 = x11 | n22683 ;
  assign n22685 = x11 & n22683 ;
  assign n35044 = ~n22685 ;
  assign n22686 = n22684 & n35044 ;
  assign n22688 = n22679 | n22686 ;
  assign n22687 = n22679 & n22686 ;
  assign n35045 = ~n22687 ;
  assign n22689 = n35045 & n22688 ;
  assign n21875 = n6272 & n34817 ;
  assign n19664 = n6190 & n34360 ;
  assign n19690 = n6244 & n34349 ;
  assign n22690 = n19664 | n19690 ;
  assign n22691 = n6217 & n34803 ;
  assign n22692 = n22690 | n22691 ;
  assign n22693 = n21875 | n22692 ;
  assign n35046 = ~n22693 ;
  assign n22694 = x11 & n35046 ;
  assign n22695 = n30180 & n22693 ;
  assign n22696 = n22694 | n22695 ;
  assign n35047 = ~n21928 ;
  assign n22697 = n35047 & n22136 ;
  assign n22698 = n22137 | n22697 ;
  assign n22699 = n22696 | n22698 ;
  assign n22700 = n22696 & n22698 ;
  assign n35048 = ~n22700 ;
  assign n22701 = n22699 & n35048 ;
  assign n35049 = ~n22132 ;
  assign n22134 = n35049 & n22133 ;
  assign n35050 = ~n22133 ;
  assign n22702 = n22132 & n35050 ;
  assign n22703 = n22134 | n22702 ;
  assign n20152 = n6272 & n34362 ;
  assign n19689 = n6190 & n34349 ;
  assign n19720 = n6244 & n34363 ;
  assign n22704 = n19689 | n19720 ;
  assign n22705 = n6217 & n34365 ;
  assign n22706 = n22704 | n22705 ;
  assign n22707 = n20152 | n22706 ;
  assign n22708 = x11 | n22707 ;
  assign n22709 = x11 & n22707 ;
  assign n35051 = ~n22709 ;
  assign n22710 = n22708 & n35051 ;
  assign n22712 = n22703 | n22710 ;
  assign n22711 = n22703 & n22710 ;
  assign n35052 = ~n22711 ;
  assign n22713 = n35052 & n22712 ;
  assign n35053 = ~n21951 ;
  assign n22130 = n35053 & n22129 ;
  assign n22714 = n22130 | n22131 ;
  assign n21073 = n6272 & n34598 ;
  assign n19714 = n6190 & n34363 ;
  assign n19738 = n6244 & n34520 ;
  assign n22715 = n19714 | n19738 ;
  assign n22716 = n6217 & n34349 ;
  assign n22717 = n22715 | n22716 ;
  assign n22718 = n21073 | n22717 ;
  assign n22719 = x11 | n22718 ;
  assign n22720 = x11 & n22718 ;
  assign n35054 = ~n22720 ;
  assign n22721 = n22719 & n35054 ;
  assign n22723 = n22714 | n22721 ;
  assign n35055 = ~n22714 ;
  assign n22722 = n35055 & n22721 ;
  assign n35056 = ~n22721 ;
  assign n22724 = n22714 & n35056 ;
  assign n22725 = n22722 | n22724 ;
  assign n22127 = n21964 & n22126 ;
  assign n22726 = n21964 | n22126 ;
  assign n35057 = ~n22127 ;
  assign n22727 = n35057 & n22726 ;
  assign n21096 = n6272 & n34603 ;
  assign n19732 = n6190 & n34520 ;
  assign n19760 = n6244 & n19752 ;
  assign n22728 = n19732 | n19760 ;
  assign n22729 = n6217 & n34596 ;
  assign n22730 = n22728 | n22729 ;
  assign n22731 = n21096 | n22730 ;
  assign n22732 = x11 | n22731 ;
  assign n22733 = x11 & n22731 ;
  assign n35058 = ~n22733 ;
  assign n22734 = n22732 & n35058 ;
  assign n22736 = n22727 | n22734 ;
  assign n35059 = ~n22727 ;
  assign n22735 = n35059 & n22734 ;
  assign n35060 = ~n22734 ;
  assign n22737 = n22727 & n35060 ;
  assign n22738 = n22735 | n22737 ;
  assign n22124 = n21977 & n22123 ;
  assign n22739 = n21977 | n22123 ;
  assign n35061 = ~n22124 ;
  assign n22740 = n35061 & n22739 ;
  assign n20809 = n6272 & n20805 ;
  assign n19762 = n6190 & n19752 ;
  assign n19780 = n6244 & n34519 ;
  assign n22741 = n19762 | n19780 ;
  assign n22742 = n6217 & n34520 ;
  assign n22743 = n22741 | n22742 ;
  assign n22744 = n20809 | n22743 ;
  assign n22745 = x11 | n22744 ;
  assign n22746 = x11 & n22744 ;
  assign n35062 = ~n22746 ;
  assign n22747 = n22745 & n35062 ;
  assign n22749 = n22740 | n22747 ;
  assign n22121 = n21989 & n22120 ;
  assign n22750 = n21989 | n22120 ;
  assign n35063 = ~n22121 ;
  assign n22751 = n35063 & n22750 ;
  assign n20837 = n6272 & n20833 ;
  assign n19779 = n6190 & n34519 ;
  assign n19814 = n6244 & n34355 ;
  assign n22752 = n19779 | n19814 ;
  assign n22753 = n6217 & n20845 ;
  assign n22754 = n22752 | n22753 ;
  assign n22755 = n20837 | n22754 ;
  assign n22756 = x11 | n22755 ;
  assign n22757 = x11 & n22755 ;
  assign n35064 = ~n22757 ;
  assign n22758 = n22756 & n35064 ;
  assign n22760 = n22751 | n22758 ;
  assign n22118 = n22001 & n22117 ;
  assign n22761 = n22001 | n22117 ;
  assign n35065 = ~n22118 ;
  assign n22762 = n35065 & n22761 ;
  assign n20868 = n6272 & n20863 ;
  assign n19806 = n6190 & n34355 ;
  assign n19828 = n6244 & n19824 ;
  assign n22763 = n19806 | n19828 ;
  assign n22764 = n6217 & n34536 ;
  assign n22765 = n22763 | n22764 ;
  assign n22766 = n20868 | n22765 ;
  assign n22767 = x11 | n22766 ;
  assign n22768 = x11 & n22766 ;
  assign n35066 = ~n22768 ;
  assign n22769 = n22767 & n35066 ;
  assign n22771 = n22762 | n22769 ;
  assign n22770 = n22762 & n22769 ;
  assign n35067 = ~n22770 ;
  assign n22772 = n35067 & n22771 ;
  assign n22115 = n22013 & n22114 ;
  assign n22773 = n22013 | n22114 ;
  assign n35068 = ~n22115 ;
  assign n22774 = n35068 & n22773 ;
  assign n20779 = n6272 & n34511 ;
  assign n19826 = n6190 & n19824 ;
  assign n20104 = n6244 & n34354 ;
  assign n22775 = n19826 | n20104 ;
  assign n22776 = n6217 & n34513 ;
  assign n22777 = n22775 | n22776 ;
  assign n22778 = n20779 | n22777 ;
  assign n22779 = x11 | n22778 ;
  assign n22780 = x11 & n22778 ;
  assign n35069 = ~n22780 ;
  assign n22781 = n22779 & n35069 ;
  assign n22783 = n22774 | n22781 ;
  assign n35070 = ~n22774 ;
  assign n22782 = n35070 & n22781 ;
  assign n35071 = ~n22781 ;
  assign n22784 = n22774 & n35071 ;
  assign n22785 = n22782 | n22784 ;
  assign n20516 = n6272 & n34442 ;
  assign n20075 = n6244 & n20067 ;
  assign n20099 = n6190 & n34354 ;
  assign n22786 = n20075 | n20099 ;
  assign n22787 = n6217 & n20527 ;
  assign n22788 = n22786 | n22787 ;
  assign n22789 = n20516 | n22788 ;
  assign n22790 = x11 | n22789 ;
  assign n22791 = x11 & n22789 ;
  assign n35072 = ~n22791 ;
  assign n22792 = n22790 & n35072 ;
  assign n22112 = n22110 & n22111 ;
  assign n22793 = n22110 | n22111 ;
  assign n35073 = ~n22112 ;
  assign n22794 = n35073 & n22793 ;
  assign n22796 = n22792 | n22794 ;
  assign n35074 = ~n22794 ;
  assign n22795 = n22792 & n35074 ;
  assign n35075 = ~n22792 ;
  assign n22797 = n35075 & n22794 ;
  assign n22798 = n22795 | n22797 ;
  assign n20547 = n6272 & n34450 ;
  assign n19861 = n6244 & n19846 ;
  assign n20068 = n6190 & n20067 ;
  assign n22799 = n19861 | n20068 ;
  assign n22800 = n6217 & n34452 ;
  assign n22801 = n22799 | n22800 ;
  assign n22802 = n20547 | n22801 ;
  assign n22803 = x11 | n22802 ;
  assign n22804 = x11 & n22802 ;
  assign n35076 = ~n22804 ;
  assign n22805 = n22803 & n35076 ;
  assign n22105 = n22051 | n22104 ;
  assign n22806 = n22051 & n22104 ;
  assign n35077 = ~n22806 ;
  assign n22807 = n22105 & n35077 ;
  assign n20588 = n6272 & n20579 ;
  assign n19849 = n6190 & n19846 ;
  assign n19886 = n6244 & n19870 ;
  assign n22808 = n19849 | n19886 ;
  assign n22809 = n6217 & n20067 ;
  assign n22810 = n22808 | n22809 ;
  assign n22811 = n20588 | n22810 ;
  assign n22812 = x11 | n22811 ;
  assign n22813 = x11 & n22811 ;
  assign n35078 = ~n22813 ;
  assign n22814 = n22812 & n35078 ;
  assign n22816 = n22807 | n22814 ;
  assign n35079 = ~n22807 ;
  assign n22815 = n35079 & n22814 ;
  assign n35080 = ~n22814 ;
  assign n22817 = n22807 & n35080 ;
  assign n22818 = n22815 | n22817 ;
  assign n35081 = ~n22100 ;
  assign n22103 = n35081 & n22101 ;
  assign n35082 = ~n22101 ;
  assign n22819 = n22100 & n35082 ;
  assign n22820 = n22103 | n22819 ;
  assign n20492 = n6272 & n20486 ;
  assign n19888 = n6190 & n19870 ;
  assign n19894 = n6244 & n19893 ;
  assign n22821 = n19888 | n19894 ;
  assign n22822 = n6217 & n19846 ;
  assign n22823 = n22821 | n22822 ;
  assign n22824 = n20492 | n22823 ;
  assign n22825 = x11 | n22824 ;
  assign n22826 = x11 & n22824 ;
  assign n35083 = ~n22826 ;
  assign n22827 = n22825 & n35083 ;
  assign n22829 = n22820 | n22827 ;
  assign n22828 = n22820 & n22827 ;
  assign n35084 = ~n22828 ;
  assign n22830 = n35084 & n22829 ;
  assign n22831 = n22087 | n22089 ;
  assign n35085 = ~n22090 ;
  assign n22832 = n35085 & n22831 ;
  assign n20318 = n6272 & n20311 ;
  assign n19907 = n6190 & n19893 ;
  assign n19933 = n6244 & n19917 ;
  assign n22833 = n19907 | n19933 ;
  assign n22834 = n6217 & n19870 ;
  assign n22835 = n22833 | n22834 ;
  assign n22836 = n20318 | n22835 ;
  assign n22837 = x11 | n22836 ;
  assign n22838 = x11 & n22836 ;
  assign n35086 = ~n22838 ;
  assign n22839 = n22837 & n35086 ;
  assign n22840 = n22832 & n22839 ;
  assign n35087 = ~n20042 ;
  assign n22066 = n35087 & n22065 ;
  assign n35088 = ~n22065 ;
  assign n22841 = n20042 & n35088 ;
  assign n22842 = n22066 | n22841 ;
  assign n35089 = ~n22074 ;
  assign n22843 = n35089 & n22842 ;
  assign n35090 = ~n22842 ;
  assign n22844 = n22074 & n35090 ;
  assign n22845 = n22843 | n22844 ;
  assign n35091 = ~n22062 ;
  assign n22063 = n22058 & n35091 ;
  assign n35092 = ~n22058 ;
  assign n22846 = n35092 & n22062 ;
  assign n22847 = n22063 | n22846 ;
  assign n20041 = n6188 & n34367 ;
  assign n20175 = n6272 & n20170 ;
  assign n22848 = n6217 & n34350 ;
  assign n22849 = n6190 & n34367 ;
  assign n22850 = n22848 | n22849 ;
  assign n22851 = n20175 | n22850 ;
  assign n22852 = n20041 | n22851 ;
  assign n22853 = x11 & n22852 ;
  assign n20013 = n6217 & n19991 ;
  assign n22854 = n6190 & n34350 ;
  assign n22855 = n6244 & n34367 ;
  assign n22856 = n22854 | n22855 ;
  assign n22857 = n20013 | n22856 ;
  assign n22858 = n6272 & n20189 ;
  assign n22859 = n22857 | n22858 ;
  assign n22861 = n22853 | n22859 ;
  assign n35093 = ~n22861 ;
  assign n22862 = x11 & n35093 ;
  assign n22864 = n20040 | n22862 ;
  assign n20211 = n6272 & n20207 ;
  assign n20011 = n6190 & n19991 ;
  assign n20033 = n6244 & n34350 ;
  assign n22865 = n20011 | n20033 ;
  assign n22866 = n6217 & n34372 ;
  assign n22867 = n22865 | n22866 ;
  assign n22868 = n20211 | n22867 ;
  assign n35094 = ~n22868 ;
  assign n22869 = x11 & n35094 ;
  assign n22870 = n30180 & n22868 ;
  assign n22871 = n22869 | n22870 ;
  assign n22872 = n22864 & n22871 ;
  assign n22873 = x14 & n20040 ;
  assign n22874 = n22056 | n22873 ;
  assign n22875 = n22056 & n22873 ;
  assign n35095 = ~n22875 ;
  assign n22876 = n22874 & n35095 ;
  assign n22878 = n22872 | n22876 ;
  assign n22877 = n22872 & n22876 ;
  assign n35096 = ~n22877 ;
  assign n22879 = n35096 & n22878 ;
  assign n20288 = n6272 & n34383 ;
  assign n19987 = n6190 & n34372 ;
  assign n20012 = n6244 & n19991 ;
  assign n22880 = n19987 | n20012 ;
  assign n22881 = n6217 & n34381 ;
  assign n22882 = n22880 | n22881 ;
  assign n22883 = n20288 | n22882 ;
  assign n35097 = ~n22883 ;
  assign n22884 = x11 & n35097 ;
  assign n22885 = n30180 & n22883 ;
  assign n22886 = n22884 | n22885 ;
  assign n35098 = ~n22886 ;
  assign n22887 = n22879 & n35098 ;
  assign n35099 = ~n22887 ;
  assign n22888 = n22878 & n35099 ;
  assign n22890 = n22847 | n22888 ;
  assign n20420 = n6272 & n20412 ;
  assign n19960 = n6190 & n34381 ;
  assign n19977 = n6244 & n34372 ;
  assign n22891 = n19960 | n19977 ;
  assign n22892 = n6217 & n19917 ;
  assign n22893 = n22891 | n22892 ;
  assign n22894 = n20420 | n22893 ;
  assign n35100 = ~n22894 ;
  assign n22895 = x11 & n35100 ;
  assign n22896 = n30180 & n22894 ;
  assign n22897 = n22895 | n22896 ;
  assign n22889 = n22847 & n22888 ;
  assign n35101 = ~n22889 ;
  assign n22898 = n35101 & n22890 ;
  assign n35102 = ~n22897 ;
  assign n22899 = n35102 & n22898 ;
  assign n35103 = ~n22899 ;
  assign n22900 = n22890 & n35103 ;
  assign n22902 = n22845 | n22900 ;
  assign n20350 = n6272 & n34399 ;
  assign n19935 = n6190 & n19917 ;
  assign n19959 = n6244 & n34381 ;
  assign n22903 = n19935 | n19959 ;
  assign n22904 = n6217 & n19893 ;
  assign n22905 = n22903 | n22904 ;
  assign n22906 = n20350 | n22905 ;
  assign n22907 = x11 | n22906 ;
  assign n22908 = x11 & n22906 ;
  assign n35104 = ~n22908 ;
  assign n22909 = n22907 & n35104 ;
  assign n22901 = n22845 & n22900 ;
  assign n35105 = ~n22901 ;
  assign n22910 = n35105 & n22902 ;
  assign n35106 = ~n22909 ;
  assign n22911 = n35106 & n22910 ;
  assign n35107 = ~n22911 ;
  assign n22912 = n22902 & n35107 ;
  assign n22913 = n22832 | n22839 ;
  assign n35108 = ~n22840 ;
  assign n22914 = n35108 & n22913 ;
  assign n22915 = n22912 & n22914 ;
  assign n22916 = n22840 | n22915 ;
  assign n35109 = ~n22916 ;
  assign n22918 = n22830 & n35109 ;
  assign n35110 = ~n22918 ;
  assign n22919 = n22829 & n35110 ;
  assign n35111 = ~n22919 ;
  assign n22921 = n22818 & n35111 ;
  assign n35112 = ~n22921 ;
  assign n22922 = n22816 & n35112 ;
  assign n22923 = n22805 & n22922 ;
  assign n22108 = n22036 & n22107 ;
  assign n22924 = n22036 | n22107 ;
  assign n35113 = ~n22108 ;
  assign n22925 = n35113 & n22924 ;
  assign n22926 = n22805 | n22922 ;
  assign n35114 = ~n22923 ;
  assign n22927 = n35114 & n22926 ;
  assign n22928 = n22925 & n22927 ;
  assign n22929 = n22923 | n22928 ;
  assign n35115 = ~n22929 ;
  assign n22931 = n22798 & n35115 ;
  assign n35116 = ~n22931 ;
  assign n22932 = n22796 & n35116 ;
  assign n35117 = ~n22932 ;
  assign n22934 = n22785 & n35117 ;
  assign n35118 = ~n22934 ;
  assign n22935 = n22783 & n35118 ;
  assign n35119 = ~n22935 ;
  assign n22937 = n22772 & n35119 ;
  assign n35120 = ~n22937 ;
  assign n22938 = n22771 & n35120 ;
  assign n22759 = n22751 & n22758 ;
  assign n35121 = ~n22759 ;
  assign n22939 = n35121 & n22760 ;
  assign n35122 = ~n22938 ;
  assign n22940 = n35122 & n22939 ;
  assign n35123 = ~n22940 ;
  assign n22941 = n22760 & n35123 ;
  assign n22748 = n22740 & n22747 ;
  assign n35124 = ~n22748 ;
  assign n22942 = n35124 & n22749 ;
  assign n35125 = ~n22941 ;
  assign n22944 = n35125 & n22942 ;
  assign n35126 = ~n22944 ;
  assign n22945 = n22749 & n35126 ;
  assign n35127 = ~n22945 ;
  assign n22947 = n22738 & n35127 ;
  assign n35128 = ~n22947 ;
  assign n22948 = n22736 & n35128 ;
  assign n35129 = ~n22948 ;
  assign n22949 = n22725 & n35129 ;
  assign n35130 = ~n22949 ;
  assign n22950 = n22723 & n35130 ;
  assign n35131 = ~n22950 ;
  assign n22952 = n22713 & n35131 ;
  assign n35132 = ~n22952 ;
  assign n22953 = n22712 & n35132 ;
  assign n35133 = ~n22953 ;
  assign n22954 = n22701 & n35133 ;
  assign n35134 = ~n22954 ;
  assign n22955 = n22699 & n35134 ;
  assign n35135 = ~n22955 ;
  assign n22957 = n22689 & n35135 ;
  assign n35136 = ~n22957 ;
  assign n22958 = n22688 & n35136 ;
  assign n35137 = ~n22958 ;
  assign n22959 = n22677 & n35137 ;
  assign n35138 = ~n22959 ;
  assign n22960 = n22675 & n35138 ;
  assign n22962 = n22664 | n22960 ;
  assign n35139 = ~n22663 ;
  assign n22963 = n35139 & n22962 ;
  assign n35140 = ~n22612 ;
  assign n22639 = n35140 & n22638 ;
  assign n22964 = n22639 | n22640 ;
  assign n22965 = n22963 | n22964 ;
  assign n35141 = ~n22640 ;
  assign n22966 = n35141 & n22965 ;
  assign n22967 = n22610 & n22966 ;
  assign n22968 = n22610 | n22966 ;
  assign n35142 = ~n22967 ;
  assign n22969 = n35142 & n22968 ;
  assign n22970 = n22215 | n22237 ;
  assign n22971 = n34921 & n22970 ;
  assign n35143 = ~n22401 ;
  assign n22402 = n22237 & n35143 ;
  assign n22972 = n34914 & n22401 ;
  assign n22973 = n22402 | n22972 ;
  assign n22974 = n1271 | n2503 ;
  assign n22975 = n5486 | n22974 ;
  assign n22976 = n797 | n996 ;
  assign n22977 = n3678 | n22976 ;
  assign n22978 = n1422 | n1472 ;
  assign n22979 = n2364 | n12731 ;
  assign n22980 = n22978 | n22979 ;
  assign n22981 = n489 | n989 ;
  assign n22982 = n575 | n22981 ;
  assign n22983 = n22980 | n22982 ;
  assign n22984 = n22977 | n22983 ;
  assign n22985 = n22975 | n22984 ;
  assign n22986 = n3906 | n12952 ;
  assign n22987 = n319 | n354 ;
  assign n22988 = n550 | n857 ;
  assign n22989 = n22987 | n22988 ;
  assign n22990 = n1528 | n22989 ;
  assign n22991 = n2395 | n2999 ;
  assign n22992 = n22990 | n22991 ;
  assign n22993 = n22986 | n22992 ;
  assign n22994 = n2581 | n22993 ;
  assign n22995 = n22985 | n22994 ;
  assign n22996 = n11238 | n14315 ;
  assign n22997 = n22995 | n22996 ;
  assign n35144 = ~n22997 ;
  assign n22998 = n22973 & n35144 ;
  assign n35145 = ~n22973 ;
  assign n22999 = n35145 & n22997 ;
  assign n23000 = n22998 | n22999 ;
  assign n13118 = n889 & n32455 ;
  assign n13054 = n3329 & n32456 ;
  assign n13098 = n3311 & n13077 ;
  assign n23001 = n13054 | n13098 ;
  assign n23002 = n3343 & n13027 ;
  assign n23003 = n23001 | n23002 ;
  assign n23004 = n13118 | n23003 ;
  assign n23005 = n23000 | n23004 ;
  assign n23006 = n23000 & n23004 ;
  assign n35146 = ~n23006 ;
  assign n23007 = n23005 & n35146 ;
  assign n23008 = n22971 & n23007 ;
  assign n23009 = n22971 | n23007 ;
  assign n35147 = ~n23008 ;
  assign n23010 = n35147 & n23009 ;
  assign n14194 = n895 & n14183 ;
  assign n14144 = n2849 & n14124 ;
  assign n14168 = n2861 & n14147 ;
  assign n23011 = n14144 | n14168 ;
  assign n23012 = n894 & n14196 ;
  assign n23013 = n23011 | n23012 ;
  assign n23014 = n14194 | n23013 ;
  assign n35148 = ~n23014 ;
  assign n23015 = x29 & n35148 ;
  assign n23016 = n30024 & n23014 ;
  assign n23017 = n23015 | n23016 ;
  assign n23018 = n23010 | n23017 ;
  assign n23019 = n23010 & n23017 ;
  assign n35149 = ~n23019 ;
  assign n23020 = n23018 & n35149 ;
  assign n23021 = n22282 | n22284 ;
  assign n35150 = ~n23021 ;
  assign n23022 = n23020 & n35150 ;
  assign n35151 = ~n23020 ;
  assign n23023 = n35151 & n23021 ;
  assign n23024 = n23022 | n23023 ;
  assign n14580 = n3791 & n14570 ;
  assign n14531 = n3802 & n32706 ;
  assign n14547 = n209 & n14536 ;
  assign n23025 = n14531 | n14547 ;
  assign n23026 = n3818 & n32707 ;
  assign n23027 = n23025 | n23026 ;
  assign n23028 = n14580 | n23027 ;
  assign n35152 = ~n23028 ;
  assign n23029 = x26 & n35152 ;
  assign n23030 = n30019 & n23028 ;
  assign n23031 = n23029 | n23030 ;
  assign n23032 = n23024 | n23031 ;
  assign n23033 = n23024 & n23031 ;
  assign n35153 = ~n23033 ;
  assign n23034 = n23032 & n35153 ;
  assign n23035 = n22167 | n22316 ;
  assign n35154 = ~n22315 ;
  assign n23036 = n35154 & n23035 ;
  assign n23037 = n23034 & n23036 ;
  assign n23038 = n23034 | n23036 ;
  assign n35155 = ~n23037 ;
  assign n23039 = n35155 & n23038 ;
  assign n15194 = n4135 & n32875 ;
  assign n15073 = n4148 & n32856 ;
  assign n15102 = n4185 & n15081 ;
  assign n23040 = n15073 | n15102 ;
  assign n23041 = n4165 & n32876 ;
  assign n23042 = n23040 | n23041 ;
  assign n23043 = n15194 | n23042 ;
  assign n23044 = x23 | n23043 ;
  assign n23045 = x23 & n23043 ;
  assign n35156 = ~n23045 ;
  assign n23046 = n23044 & n35156 ;
  assign n23048 = n23039 | n23046 ;
  assign n35157 = ~n23039 ;
  assign n23047 = n35157 & n23046 ;
  assign n35158 = ~n23046 ;
  assign n23049 = n23039 & n35158 ;
  assign n23050 = n23047 | n23049 ;
  assign n35159 = ~n22354 ;
  assign n23051 = n35159 & n22356 ;
  assign n35160 = ~n23051 ;
  assign n23053 = n23050 & n35160 ;
  assign n35161 = ~n23053 ;
  assign n23054 = n23048 & n35161 ;
  assign n4725 = x20 & n4724 ;
  assign n15242 = x19 & n15221 ;
  assign n15237 = x20 & n32883 ;
  assign n23055 = n4724 | n15237 ;
  assign n23056 = n15242 | n23055 ;
  assign n35162 = ~n4725 ;
  assign n23057 = n35162 & n23056 ;
  assign n23058 = n23054 & n23057 ;
  assign n15294 = n3791 & n15288 ;
  assign n14510 = n3802 & n32707 ;
  assign n14523 = n209 & n32706 ;
  assign n23059 = n14510 | n14523 ;
  assign n23060 = n3818 & n15081 ;
  assign n23061 = n23059 | n23060 ;
  assign n23062 = n15294 | n23061 ;
  assign n35163 = ~n23062 ;
  assign n23063 = x26 & n35163 ;
  assign n23064 = n30019 & n23062 ;
  assign n23065 = n23063 | n23064 ;
  assign n14975 = n895 & n14965 ;
  assign n14119 = n2849 & n14101 ;
  assign n14127 = n2861 & n14124 ;
  assign n23066 = n14119 | n14127 ;
  assign n23067 = n894 & n14536 ;
  assign n23068 = n23066 | n23067 ;
  assign n23069 = n14975 | n23068 ;
  assign n35164 = ~n23069 ;
  assign n23070 = x29 & n35164 ;
  assign n23071 = n30024 & n23069 ;
  assign n23072 = n23070 | n23071 ;
  assign n35165 = ~n22971 ;
  assign n23073 = n35165 & n23007 ;
  assign n35166 = ~n23073 ;
  assign n23074 = n23005 & n35166 ;
  assign n23075 = n22237 | n22401 ;
  assign n23076 = n22973 & n22997 ;
  assign n35167 = ~n23076 ;
  assign n23077 = n23075 & n35167 ;
  assign n23078 = n1718 | n2122 ;
  assign n23079 = n5378 | n23078 ;
  assign n23080 = n630 | n989 ;
  assign n23081 = n1308 | n23080 ;
  assign n23082 = n5321 | n23081 ;
  assign n23083 = n23079 | n23082 ;
  assign n23084 = n249 | n764 ;
  assign n23085 = n1049 | n23084 ;
  assign n23086 = n2029 | n23085 ;
  assign n23087 = n2722 | n23086 ;
  assign n23088 = n130 | n221 ;
  assign n23089 = n684 | n23088 ;
  assign n23090 = n4073 | n23089 ;
  assign n23091 = n472 | n23090 ;
  assign n23092 = n2991 | n23091 ;
  assign n23093 = n23087 | n23092 ;
  assign n23094 = n23083 | n23093 ;
  assign n23095 = n1146 | n2140 ;
  assign n23096 = n2686 | n2767 ;
  assign n23097 = n23095 | n23096 ;
  assign n23098 = n682 | n750 ;
  assign n23099 = n811 | n23098 ;
  assign n23100 = n384 | n447 ;
  assign n23101 = n23099 | n23100 ;
  assign n23102 = n11127 | n23101 ;
  assign n23103 = n23097 | n23102 ;
  assign n23104 = n270 | n272 ;
  assign n23105 = n310 | n23104 ;
  assign n23106 = n553 | n13252 ;
  assign n23107 = n23105 | n23106 ;
  assign n23108 = n13721 | n23107 ;
  assign n23109 = n203 | n320 ;
  assign n23110 = n506 | n23109 ;
  assign n23111 = n337 | n428 ;
  assign n35168 = ~n23111 ;
  assign n23112 = n11669 & n35168 ;
  assign n35169 = ~n23110 ;
  assign n23113 = n35169 & n23112 ;
  assign n35170 = ~n23108 ;
  assign n23114 = n35170 & n23113 ;
  assign n35171 = ~n23103 ;
  assign n23115 = n35171 & n23114 ;
  assign n35172 = ~n22993 ;
  assign n23116 = n35172 & n23115 ;
  assign n35173 = ~n2599 ;
  assign n23117 = n35173 & n23116 ;
  assign n35174 = ~n23094 ;
  assign n23118 = n35174 & n23117 ;
  assign n23119 = n23077 & n23118 ;
  assign n23120 = n23077 | n23118 ;
  assign n35175 = ~n23119 ;
  assign n23121 = n35175 & n23120 ;
  assign n14665 = n889 & n14655 ;
  assign n13045 = n3329 & n13027 ;
  assign n13071 = n3311 & n32456 ;
  assign n23122 = n13045 | n13071 ;
  assign n23123 = n3343 & n14147 ;
  assign n23124 = n23122 | n23123 ;
  assign n23125 = n14665 | n23124 ;
  assign n35176 = ~n23125 ;
  assign n23126 = n23121 & n35176 ;
  assign n35177 = ~n23121 ;
  assign n23127 = n35177 & n23125 ;
  assign n23128 = n23126 | n23127 ;
  assign n35178 = ~n23128 ;
  assign n23129 = n23074 & n35178 ;
  assign n35179 = ~n23074 ;
  assign n23130 = n35179 & n23128 ;
  assign n23131 = n23129 | n23130 ;
  assign n23132 = n23072 | n23131 ;
  assign n23133 = n23072 & n23131 ;
  assign n35180 = ~n23133 ;
  assign n23134 = n23132 & n35180 ;
  assign n35181 = ~n23022 ;
  assign n23135 = n23018 & n35181 ;
  assign n23136 = n23134 & n23135 ;
  assign n23137 = n23134 | n23135 ;
  assign n35182 = ~n23136 ;
  assign n23138 = n35182 & n23137 ;
  assign n23139 = n23065 | n23138 ;
  assign n23140 = n23065 & n23138 ;
  assign n35183 = ~n23140 ;
  assign n23141 = n23139 & n35183 ;
  assign n35184 = ~n23036 ;
  assign n23142 = n23034 & n35184 ;
  assign n35185 = ~n23142 ;
  assign n23143 = n23032 & n35185 ;
  assign n23144 = n23141 & n23143 ;
  assign n23145 = n23141 | n23143 ;
  assign n35186 = ~n23144 ;
  assign n23146 = n35186 & n23145 ;
  assign n15266 = n4135 & n32889 ;
  assign n15074 = n4185 & n32856 ;
  assign n15176 = n4148 & n32876 ;
  assign n23147 = n15074 | n15176 ;
  assign n23148 = n4165 & n32890 ;
  assign n23149 = n23147 | n23148 ;
  assign n23150 = n15266 | n23149 ;
  assign n35187 = ~n23150 ;
  assign n23151 = x23 & n35187 ;
  assign n23152 = n30030 & n23150 ;
  assign n23153 = n23151 | n23152 ;
  assign n23154 = n23146 | n23153 ;
  assign n23155 = n23146 & n23153 ;
  assign n35188 = ~n23155 ;
  assign n23156 = n23154 & n35188 ;
  assign n23157 = n23054 | n23057 ;
  assign n35189 = ~n23058 ;
  assign n23158 = n35189 & n23157 ;
  assign n35190 = ~n23156 ;
  assign n23160 = n35190 & n23158 ;
  assign n23161 = n23058 | n23160 ;
  assign n35191 = ~n23077 ;
  assign n23162 = n35191 & n23118 ;
  assign n23163 = n23127 | n23162 ;
  assign n23164 = n512 | n538 ;
  assign n23165 = n630 | n23164 ;
  assign n23166 = n359 | n506 ;
  assign n23167 = n428 | n23166 ;
  assign n23168 = n23165 | n23167 ;
  assign n23169 = n291 | n11154 ;
  assign n23170 = n23168 | n23169 ;
  assign n23171 = n788 | n2410 ;
  assign n23172 = n4310 | n5806 ;
  assign n23173 = n23171 | n23172 ;
  assign n23174 = n1014 | n23173 ;
  assign n23175 = n332 | n1099 ;
  assign n23176 = n1126 | n23175 ;
  assign n23177 = n464 | n631 ;
  assign n23178 = n4010 | n23177 ;
  assign n23179 = n23176 | n23178 ;
  assign n23180 = n23174 | n23179 ;
  assign n23181 = n23170 | n23180 ;
  assign n23182 = n1852 | n23181 ;
  assign n23183 = n3294 & n32117 ;
  assign n35192 = ~n23182 ;
  assign n23184 = n35192 & n23183 ;
  assign n35193 = ~n23118 ;
  assign n23185 = n35193 & n23184 ;
  assign n35194 = ~n23184 ;
  assign n23186 = n23118 & n35194 ;
  assign n23187 = n23185 | n23186 ;
  assign n14294 = n889 & n14283 ;
  assign n13033 = n3311 & n13027 ;
  assign n14165 = n3329 & n14147 ;
  assign n23188 = n13033 | n14165 ;
  assign n23189 = n3343 & n14295 ;
  assign n23190 = n23188 | n23189 ;
  assign n23191 = n14294 | n23190 ;
  assign n35195 = ~n23191 ;
  assign n23192 = n23187 & n35195 ;
  assign n35196 = ~n23187 ;
  assign n23194 = n35196 & n23191 ;
  assign n23195 = n23192 | n23194 ;
  assign n35197 = ~n23195 ;
  assign n23196 = n23163 & n35197 ;
  assign n35198 = ~n23163 ;
  assign n23197 = n35198 & n23195 ;
  assign n23198 = n23196 | n23197 ;
  assign n35199 = ~n23130 ;
  assign n23199 = n35199 & n23132 ;
  assign n35200 = ~n23198 ;
  assign n23200 = n35200 & n23199 ;
  assign n35201 = ~n23199 ;
  assign n23201 = n23198 & n35201 ;
  assign n23202 = n23200 | n23201 ;
  assign n14690 = n895 & n32735 ;
  assign n14109 = n2861 & n14101 ;
  assign n14554 = n2849 & n14536 ;
  assign n23203 = n14109 | n14554 ;
  assign n23204 = n894 & n32706 ;
  assign n23205 = n23203 | n23204 ;
  assign n23206 = n14690 | n23205 ;
  assign n23207 = x29 | n23206 ;
  assign n23208 = x29 & n23206 ;
  assign n35202 = ~n23208 ;
  assign n23209 = n23207 & n35202 ;
  assign n23210 = n23202 & n23209 ;
  assign n23211 = n23202 | n23209 ;
  assign n35203 = ~n23210 ;
  assign n23212 = n35203 & n23211 ;
  assign n15119 = n3791 & n15111 ;
  assign n14500 = n209 & n32707 ;
  assign n15103 = n3802 & n15081 ;
  assign n23213 = n14500 | n15103 ;
  assign n23214 = n3818 & n32856 ;
  assign n23215 = n23213 | n23214 ;
  assign n23216 = n15119 | n23215 ;
  assign n35204 = ~n23216 ;
  assign n23217 = x26 & n35204 ;
  assign n23218 = n30019 & n23216 ;
  assign n23219 = n23217 | n23218 ;
  assign n35205 = ~n23219 ;
  assign n23220 = n23212 & n35205 ;
  assign n35206 = ~n23212 ;
  assign n23221 = n35206 & n23219 ;
  assign n23222 = n23220 | n23221 ;
  assign n15535 = n4135 & n15526 ;
  assign n15177 = n4185 & n32876 ;
  assign n15227 = n4165 & n15221 ;
  assign n23223 = n15177 | n15227 ;
  assign n23224 = n4148 & n32890 ;
  assign n23225 = n23223 | n23224 ;
  assign n23226 = n15535 | n23225 ;
  assign n23227 = x23 | n23226 ;
  assign n23228 = x23 & n23226 ;
  assign n35207 = ~n23228 ;
  assign n23229 = n23227 & n35207 ;
  assign n35208 = ~n23135 ;
  assign n23230 = n23134 & n35208 ;
  assign n35209 = ~n23230 ;
  assign n23231 = n23139 & n35209 ;
  assign n23232 = n23229 & n23231 ;
  assign n23233 = n23229 | n23231 ;
  assign n35210 = ~n23232 ;
  assign n23234 = n35210 & n23233 ;
  assign n35211 = ~n23222 ;
  assign n23235 = n35211 & n23234 ;
  assign n35212 = ~n23234 ;
  assign n23236 = n23222 & n35212 ;
  assign n23237 = n23235 | n23236 ;
  assign n4682 = x19 | n4680 ;
  assign n23238 = n4682 & n35162 ;
  assign n35213 = ~n23143 ;
  assign n23239 = n23141 & n35213 ;
  assign n35214 = ~n23239 ;
  assign n23240 = n23154 & n35214 ;
  assign n23241 = n23238 & n23240 ;
  assign n23242 = n23238 | n23240 ;
  assign n35215 = ~n23241 ;
  assign n23243 = n35215 & n23242 ;
  assign n23244 = n23237 & n23243 ;
  assign n23245 = n23237 | n23243 ;
  assign n35216 = ~n23244 ;
  assign n23246 = n35216 & n23245 ;
  assign n35217 = ~n23161 ;
  assign n23247 = n35217 & n23246 ;
  assign n35218 = ~n23246 ;
  assign n23248 = n23161 & n35218 ;
  assign n23249 = n23247 | n23248 ;
  assign n23159 = n23156 & n23158 ;
  assign n23250 = n23156 | n23158 ;
  assign n35219 = ~n23159 ;
  assign n23251 = n35219 & n23250 ;
  assign n15518 = n4683 & n15516 ;
  assign n15243 = n4706 & n15221 ;
  assign n23252 = n4748 | n15243 ;
  assign n23253 = n4726 & n32890 ;
  assign n23254 = n23252 | n23253 ;
  assign n23255 = n15518 | n23254 ;
  assign n35220 = ~n23255 ;
  assign n23256 = x20 & n35220 ;
  assign n23257 = n30374 & n23255 ;
  assign n23258 = n23256 | n23257 ;
  assign n35221 = ~n22358 ;
  assign n23259 = n35221 & n22397 ;
  assign n23260 = n22395 | n23259 ;
  assign n23261 = n23258 | n23260 ;
  assign n23052 = n23050 & n23051 ;
  assign n23262 = n23050 | n23051 ;
  assign n35222 = ~n23052 ;
  assign n23263 = n35222 & n23262 ;
  assign n23264 = n23258 & n23260 ;
  assign n35223 = ~n23264 ;
  assign n23265 = n23261 & n35223 ;
  assign n35224 = ~n23263 ;
  assign n23266 = n35224 & n23265 ;
  assign n35225 = ~n23266 ;
  assign n23267 = n23261 & n35225 ;
  assign n35226 = ~n23267 ;
  assign n23269 = n23251 & n35226 ;
  assign n35227 = ~n23251 ;
  assign n23268 = n35227 & n23267 ;
  assign n23270 = n23268 | n23269 ;
  assign n35228 = ~n23265 ;
  assign n23271 = n23263 & n35228 ;
  assign n23272 = n23266 | n23271 ;
  assign n23273 = n22437 & n34981 ;
  assign n23275 = n23272 | n23273 ;
  assign n35229 = ~n23272 ;
  assign n23274 = n35229 & n23273 ;
  assign n35230 = ~n23273 ;
  assign n23276 = n23272 & n35230 ;
  assign n23277 = n23274 | n23276 ;
  assign n35231 = ~n22469 ;
  assign n23278 = n22442 & n35231 ;
  assign n23279 = n22472 | n22506 ;
  assign n35232 = ~n23278 ;
  assign n23280 = n35232 & n23279 ;
  assign n35233 = ~n23280 ;
  assign n23283 = n23277 & n35233 ;
  assign n35234 = ~n23283 ;
  assign n23284 = n23275 & n35234 ;
  assign n23285 = n23270 | n23284 ;
  assign n35235 = ~n23269 ;
  assign n23286 = n35235 & n23285 ;
  assign n35236 = ~n23249 ;
  assign n23287 = n35236 & n23286 ;
  assign n35237 = ~n23286 ;
  assign n23289 = n23249 & n35237 ;
  assign n23290 = n23287 | n23289 ;
  assign n35238 = ~n23270 ;
  assign n23313 = n35238 & n23284 ;
  assign n35239 = ~n23284 ;
  assign n23315 = n23270 & n35239 ;
  assign n23316 = n23313 | n23315 ;
  assign n23281 = n23277 & n23280 ;
  assign n23338 = n23277 | n23280 ;
  assign n35240 = ~n23281 ;
  assign n23339 = n35240 & n23338 ;
  assign n23365 = n35020 & n22562 ;
  assign n23366 = n23339 | n23365 ;
  assign n23367 = n23316 | n23366 ;
  assign n23362 = n22509 & n35019 ;
  assign n35241 = ~n23362 ;
  assign n23364 = n23339 & n35241 ;
  assign n23368 = n23316 & n23364 ;
  assign n35242 = ~n23368 ;
  assign n23369 = n23367 & n35242 ;
  assign n23370 = n23290 | n23369 ;
  assign n23371 = n23290 & n23369 ;
  assign n35243 = ~n23371 ;
  assign n23372 = n23370 & n35243 ;
  assign n23373 = n7068 & n23372 ;
  assign n35244 = ~n23316 ;
  assign n23322 = n69 & n35244 ;
  assign n23352 = n7041 & n23339 ;
  assign n23386 = n23322 | n23352 ;
  assign n23288 = n23249 & n23286 ;
  assign n23384 = n23249 | n23286 ;
  assign n35245 = ~n23288 ;
  assign n23385 = n35245 & n23384 ;
  assign n35246 = ~n23385 ;
  assign n23387 = n7017 & n35246 ;
  assign n23388 = n23386 | n23387 ;
  assign n23389 = n23373 | n23388 ;
  assign n23390 = x8 | n23389 ;
  assign n23391 = x8 & n23389 ;
  assign n35247 = ~n23391 ;
  assign n23392 = n23390 & n35247 ;
  assign n23393 = n22969 & n23392 ;
  assign n23394 = n22969 | n23392 ;
  assign n35248 = ~n23393 ;
  assign n23395 = n35248 & n23394 ;
  assign n23396 = n22963 & n22964 ;
  assign n35249 = ~n23396 ;
  assign n23397 = n22965 & n35249 ;
  assign n23363 = n23339 & n23362 ;
  assign n35250 = ~n23339 ;
  assign n23398 = n35250 & n23365 ;
  assign n23399 = n23363 | n23398 ;
  assign n23400 = n35244 & n23399 ;
  assign n35251 = ~n23399 ;
  assign n23401 = n23316 & n35251 ;
  assign n23402 = n23400 | n23401 ;
  assign n35252 = ~n23402 ;
  assign n23403 = n7068 & n35252 ;
  assign n22522 = n7041 & n35020 ;
  assign n23350 = n69 & n23339 ;
  assign n23415 = n22522 | n23350 ;
  assign n23314 = n23270 & n23284 ;
  assign n35253 = ~n23314 ;
  assign n23414 = n23285 & n35253 ;
  assign n35254 = ~n23414 ;
  assign n23416 = n7017 & n35254 ;
  assign n23417 = n23415 | n23416 ;
  assign n23418 = n23403 | n23417 ;
  assign n23419 = x8 | n23418 ;
  assign n23420 = x8 & n23418 ;
  assign n35255 = ~n23420 ;
  assign n23421 = n23419 & n35255 ;
  assign n35256 = ~n23421 ;
  assign n23423 = n23397 & n35256 ;
  assign n23422 = n23397 & n23421 ;
  assign n23424 = n23397 | n23421 ;
  assign n35257 = ~n23422 ;
  assign n23425 = n35257 & n23424 ;
  assign n35258 = ~n22664 ;
  assign n22961 = n35258 & n22960 ;
  assign n35259 = ~n22960 ;
  assign n23426 = n22664 & n35259 ;
  assign n23427 = n22961 | n23426 ;
  assign n22577 = n22509 & n22559 ;
  assign n23428 = n22509 | n22562 ;
  assign n35260 = ~n22577 ;
  assign n23429 = n35260 & n23428 ;
  assign n35261 = ~n23429 ;
  assign n23430 = n23339 & n35261 ;
  assign n23431 = n35250 & n23429 ;
  assign n23432 = n23430 | n23431 ;
  assign n35262 = ~n23432 ;
  assign n23433 = n7068 & n35262 ;
  assign n22519 = n69 & n35020 ;
  assign n22587 = n7041 & n22533 ;
  assign n23445 = n22519 | n22587 ;
  assign n35263 = ~n23277 ;
  assign n23282 = n35263 & n23280 ;
  assign n23444 = n23282 | n23283 ;
  assign n23446 = n7017 & n23444 ;
  assign n23447 = n23445 | n23446 ;
  assign n23448 = n23433 | n23447 ;
  assign n23449 = x8 | n23448 ;
  assign n23450 = x8 & n23448 ;
  assign n35264 = ~n23450 ;
  assign n23451 = n23449 & n35264 ;
  assign n35265 = ~n23451 ;
  assign n23453 = n23427 & n35265 ;
  assign n35266 = ~n23427 ;
  assign n23452 = n35266 & n23451 ;
  assign n23454 = n23452 | n23453 ;
  assign n22568 = n7068 & n35022 ;
  assign n22543 = n7041 & n35018 ;
  assign n22586 = n69 & n22533 ;
  assign n23455 = n22543 | n22586 ;
  assign n23456 = n7017 & n35020 ;
  assign n23457 = n23455 | n23456 ;
  assign n23458 = n22568 | n23457 ;
  assign n23459 = x8 | n23458 ;
  assign n23460 = x8 & n23458 ;
  assign n35267 = ~n23460 ;
  assign n23461 = n23459 & n35267 ;
  assign n22956 = n22689 & n22955 ;
  assign n23462 = n22689 | n22955 ;
  assign n35268 = ~n22956 ;
  assign n23463 = n35268 & n23462 ;
  assign n22624 = n7068 & n35030 ;
  assign n21738 = n7041 & n21729 ;
  assign n22549 = n69 & n35018 ;
  assign n23464 = n21738 | n22549 ;
  assign n23465 = n7017 & n22533 ;
  assign n23466 = n23464 | n23465 ;
  assign n23467 = n22624 | n23466 ;
  assign n23468 = x8 | n23467 ;
  assign n23469 = x8 & n23467 ;
  assign n35269 = ~n23469 ;
  assign n23470 = n23468 & n35269 ;
  assign n23472 = n23463 | n23470 ;
  assign n35270 = ~n23463 ;
  assign n23471 = n35270 & n23470 ;
  assign n35271 = ~n23470 ;
  assign n23473 = n23463 & n35271 ;
  assign n23474 = n23471 | n23473 ;
  assign n22645 = n7068 & n35035 ;
  assign n21736 = n69 & n21729 ;
  assign n21815 = n7041 & n21753 ;
  assign n23475 = n21736 | n21815 ;
  assign n23476 = n7017 & n35018 ;
  assign n23477 = n23475 | n23476 ;
  assign n23478 = n22645 | n23477 ;
  assign n23479 = x8 | n23478 ;
  assign n23480 = x8 & n23478 ;
  assign n35272 = ~n23480 ;
  assign n23481 = n23479 & n35272 ;
  assign n22951 = n22713 & n22950 ;
  assign n23482 = n22713 | n22950 ;
  assign n35273 = ~n22951 ;
  assign n23483 = n35273 & n23482 ;
  assign n21794 = n7068 & n34802 ;
  assign n21760 = n7041 & n34803 ;
  assign n21817 = n69 & n21753 ;
  assign n23484 = n21760 | n21817 ;
  assign n23485 = n7017 & n21804 ;
  assign n23486 = n23484 | n23485 ;
  assign n23487 = n21794 | n23486 ;
  assign n23488 = x8 | n23487 ;
  assign n23489 = x8 & n23487 ;
  assign n35274 = ~n23489 ;
  assign n23490 = n23488 & n35274 ;
  assign n23492 = n23483 | n23490 ;
  assign n35275 = ~n22725 ;
  assign n23493 = n35275 & n22948 ;
  assign n23494 = n22949 | n23493 ;
  assign n21852 = n7068 & n21848 ;
  assign n19661 = n7041 & n34360 ;
  assign n21766 = n69 & n34803 ;
  assign n23495 = n19661 | n21766 ;
  assign n23496 = n7017 & n21753 ;
  assign n23497 = n23495 | n23496 ;
  assign n23498 = n21852 | n23497 ;
  assign n23499 = x8 | n23498 ;
  assign n23500 = x8 & n23498 ;
  assign n35276 = ~n23500 ;
  assign n23501 = n23499 & n35276 ;
  assign n23503 = n23494 | n23501 ;
  assign n23502 = n23494 & n23501 ;
  assign n35277 = ~n23502 ;
  assign n23504 = n35277 & n23503 ;
  assign n35278 = ~n22738 ;
  assign n22946 = n35278 & n22945 ;
  assign n23505 = n22946 | n22947 ;
  assign n21877 = n7068 & n34817 ;
  assign n19669 = n69 & n34360 ;
  assign n19696 = n7041 & n34349 ;
  assign n23506 = n19669 | n19696 ;
  assign n23507 = n7017 & n34803 ;
  assign n23508 = n23506 | n23507 ;
  assign n23509 = n21877 | n23508 ;
  assign n23510 = x8 | n23509 ;
  assign n23511 = x8 & n23509 ;
  assign n35279 = ~n23511 ;
  assign n23512 = n23510 & n35279 ;
  assign n23514 = n23505 | n23512 ;
  assign n35280 = ~n23505 ;
  assign n23513 = n35280 & n23512 ;
  assign n35281 = ~n23512 ;
  assign n23515 = n23505 & n35281 ;
  assign n23516 = n23513 | n23515 ;
  assign n20154 = n7068 & n34362 ;
  assign n19686 = n69 & n34349 ;
  assign n19711 = n7041 & n34363 ;
  assign n23517 = n19686 | n19711 ;
  assign n23518 = n7017 & n34365 ;
  assign n23519 = n23517 | n23518 ;
  assign n23520 = n20154 | n23519 ;
  assign n23521 = x8 | n23520 ;
  assign n23522 = x8 & n23520 ;
  assign n35282 = ~n23522 ;
  assign n23523 = n23521 & n35282 ;
  assign n22943 = n22941 & n22942 ;
  assign n23524 = n22941 | n22942 ;
  assign n35283 = ~n22943 ;
  assign n23525 = n35283 & n23524 ;
  assign n23526 = n23523 | n23525 ;
  assign n35284 = ~n22939 ;
  assign n23527 = n22938 & n35284 ;
  assign n23528 = n22940 | n23527 ;
  assign n21074 = n7068 & n34598 ;
  assign n19721 = n69 & n34363 ;
  assign n19735 = n7041 & n34520 ;
  assign n23529 = n19721 | n19735 ;
  assign n23530 = n7017 & n34349 ;
  assign n23531 = n23529 | n23530 ;
  assign n23532 = n21074 | n23531 ;
  assign n23533 = x8 | n23532 ;
  assign n23534 = x8 & n23532 ;
  assign n35285 = ~n23534 ;
  assign n23535 = n23533 & n35285 ;
  assign n23537 = n23528 & n23535 ;
  assign n35286 = ~n23528 ;
  assign n23536 = n35286 & n23535 ;
  assign n35287 = ~n23535 ;
  assign n23538 = n23528 & n35287 ;
  assign n23539 = n23536 | n23538 ;
  assign n35288 = ~n22772 ;
  assign n22936 = n35288 & n22935 ;
  assign n23540 = n22936 | n22937 ;
  assign n21098 = n7068 & n34603 ;
  assign n19744 = n69 & n34520 ;
  assign n19757 = n7041 & n19752 ;
  assign n23541 = n19744 | n19757 ;
  assign n23542 = n7017 & n34596 ;
  assign n23543 = n23541 | n23542 ;
  assign n23544 = n21098 | n23543 ;
  assign n23545 = x8 | n23544 ;
  assign n23546 = x8 & n23544 ;
  assign n35289 = ~n23546 ;
  assign n23547 = n23545 & n35289 ;
  assign n23549 = n23540 | n23547 ;
  assign n22933 = n22785 & n22932 ;
  assign n23550 = n22785 | n22932 ;
  assign n35290 = ~n22933 ;
  assign n23551 = n35290 & n23550 ;
  assign n20810 = n7068 & n20805 ;
  assign n19756 = n69 & n19752 ;
  assign n19777 = n7041 & n34519 ;
  assign n23552 = n19756 | n19777 ;
  assign n23553 = n7017 & n34520 ;
  assign n23554 = n23552 | n23553 ;
  assign n23555 = n20810 | n23554 ;
  assign n23556 = x8 | n23555 ;
  assign n23557 = x8 & n23555 ;
  assign n35291 = ~n23557 ;
  assign n23558 = n23556 & n35291 ;
  assign n23560 = n23551 | n23558 ;
  assign n35292 = ~n23551 ;
  assign n23559 = n35292 & n23558 ;
  assign n35293 = ~n23558 ;
  assign n23561 = n23551 & n35293 ;
  assign n23562 = n23559 | n23561 ;
  assign n20839 = n7068 & n20833 ;
  assign n19789 = n69 & n34519 ;
  assign n19805 = n7041 & n34355 ;
  assign n23563 = n19789 | n19805 ;
  assign n23564 = n7017 & n20845 ;
  assign n23565 = n23563 | n23564 ;
  assign n23566 = n20839 | n23565 ;
  assign n23567 = x8 | n23566 ;
  assign n23568 = x8 & n23566 ;
  assign n35294 = ~n23568 ;
  assign n23569 = n23567 & n35294 ;
  assign n23570 = n22925 | n22927 ;
  assign n35295 = ~n22928 ;
  assign n23571 = n35295 & n23570 ;
  assign n20869 = n7068 & n20863 ;
  assign n19803 = n69 & n34355 ;
  assign n19825 = n7041 & n19824 ;
  assign n23572 = n19803 | n19825 ;
  assign n23573 = n7017 & n34536 ;
  assign n23574 = n23572 | n23573 ;
  assign n23575 = n20869 | n23574 ;
  assign n23576 = x8 | n23575 ;
  assign n23577 = x8 & n23575 ;
  assign n35296 = ~n23577 ;
  assign n23578 = n23576 & n35296 ;
  assign n23580 = n23571 | n23578 ;
  assign n23579 = n23571 & n23578 ;
  assign n35297 = ~n23579 ;
  assign n23581 = n35297 & n23580 ;
  assign n22920 = n22818 & n22919 ;
  assign n23582 = n22818 | n22919 ;
  assign n35298 = ~n22920 ;
  assign n23583 = n35298 & n23582 ;
  assign n20781 = n7068 & n34511 ;
  assign n19839 = n69 & n19824 ;
  assign n20095 = n7041 & n34354 ;
  assign n23584 = n19839 | n20095 ;
  assign n23585 = n7017 & n34513 ;
  assign n23586 = n23584 | n23585 ;
  assign n23587 = n20781 | n23586 ;
  assign n23588 = x8 | n23587 ;
  assign n23589 = x8 & n23587 ;
  assign n35299 = ~n23589 ;
  assign n23590 = n23588 & n35299 ;
  assign n23592 = n23583 | n23590 ;
  assign n23591 = n23583 & n23590 ;
  assign n35300 = ~n23591 ;
  assign n23593 = n35300 & n23592 ;
  assign n22917 = n22830 | n22916 ;
  assign n23594 = n22830 & n22916 ;
  assign n35301 = ~n23594 ;
  assign n23595 = n22917 & n35301 ;
  assign n20521 = n7068 & n34442 ;
  assign n20083 = n7041 & n20067 ;
  assign n20108 = n69 & n34354 ;
  assign n23596 = n20083 | n20108 ;
  assign n23597 = n7017 & n20527 ;
  assign n23598 = n23596 | n23597 ;
  assign n23599 = n20521 | n23598 ;
  assign n23600 = x8 | n23599 ;
  assign n23601 = x8 & n23599 ;
  assign n35302 = ~n23601 ;
  assign n23602 = n23600 & n35302 ;
  assign n23604 = n23595 | n23602 ;
  assign n35303 = ~n23595 ;
  assign n23603 = n35303 & n23602 ;
  assign n35304 = ~n23602 ;
  assign n23605 = n23595 & n35304 ;
  assign n23606 = n23603 | n23605 ;
  assign n20551 = n7068 & n34450 ;
  assign n19862 = n7041 & n19846 ;
  assign n20082 = n69 & n20067 ;
  assign n23607 = n19862 | n20082 ;
  assign n23608 = n7017 & n34452 ;
  assign n23609 = n23607 | n23608 ;
  assign n23610 = n20551 | n23609 ;
  assign n23611 = x8 | n23610 ;
  assign n23612 = x8 & n23610 ;
  assign n35305 = ~n23612 ;
  assign n23613 = n23611 & n35305 ;
  assign n23614 = n22912 | n22914 ;
  assign n35306 = ~n22915 ;
  assign n23615 = n35306 & n23614 ;
  assign n23617 = n23613 | n23615 ;
  assign n23616 = n23613 & n23615 ;
  assign n35307 = ~n23616 ;
  assign n23618 = n35307 & n23617 ;
  assign n35308 = ~n22910 ;
  assign n23619 = n22909 & n35308 ;
  assign n23620 = n22911 | n23619 ;
  assign n20582 = n7068 & n20579 ;
  assign n19863 = n69 & n19846 ;
  assign n19887 = n7041 & n19870 ;
  assign n23621 = n19863 | n19887 ;
  assign n23622 = n7017 & n20067 ;
  assign n23623 = n23621 | n23622 ;
  assign n23624 = n20582 | n23623 ;
  assign n23625 = x8 | n23624 ;
  assign n23626 = x8 & n23624 ;
  assign n35309 = ~n23626 ;
  assign n23627 = n23625 & n35309 ;
  assign n23629 = n23620 | n23627 ;
  assign n35310 = ~n23620 ;
  assign n23628 = n35310 & n23627 ;
  assign n35311 = ~n23627 ;
  assign n23630 = n23620 & n35311 ;
  assign n23631 = n23628 | n23630 ;
  assign n35312 = ~n22898 ;
  assign n23632 = n22897 & n35312 ;
  assign n23633 = n22899 | n23632 ;
  assign n20493 = n7068 & n20486 ;
  assign n19881 = n69 & n19870 ;
  assign n19903 = n7041 & n19893 ;
  assign n23634 = n19881 | n19903 ;
  assign n23635 = n7017 & n19846 ;
  assign n23636 = n23634 | n23635 ;
  assign n23637 = n20493 | n23636 ;
  assign n23638 = x8 | n23637 ;
  assign n23639 = x8 & n23637 ;
  assign n35313 = ~n23639 ;
  assign n23640 = n23638 & n35313 ;
  assign n23642 = n23633 | n23640 ;
  assign n23641 = n23633 & n23640 ;
  assign n35314 = ~n23641 ;
  assign n23643 = n35314 & n23642 ;
  assign n35315 = ~n22879 ;
  assign n23644 = n35315 & n22886 ;
  assign n23645 = n22887 | n23644 ;
  assign n20319 = n7068 & n20311 ;
  assign n19909 = n69 & n19893 ;
  assign n19929 = n7041 & n19917 ;
  assign n23646 = n19909 | n19929 ;
  assign n23647 = n7017 & n19870 ;
  assign n23648 = n23646 | n23647 ;
  assign n23649 = n20319 | n23648 ;
  assign n23650 = x8 | n23649 ;
  assign n23651 = x8 & n23649 ;
  assign n35316 = ~n23651 ;
  assign n23652 = n23650 & n35316 ;
  assign n23654 = n23645 | n23652 ;
  assign n23653 = n23645 & n23652 ;
  assign n35317 = ~n23653 ;
  assign n23655 = n35317 & n23654 ;
  assign n35318 = ~n20040 ;
  assign n22863 = n35318 & n22862 ;
  assign n35319 = ~n22862 ;
  assign n23656 = n20040 & n35319 ;
  assign n23657 = n22863 | n23656 ;
  assign n35320 = ~n22871 ;
  assign n23658 = n35320 & n23657 ;
  assign n35321 = ~n23657 ;
  assign n23659 = n22871 & n35321 ;
  assign n23660 = n23658 | n23659 ;
  assign n22860 = n22853 & n22859 ;
  assign n35322 = ~n22860 ;
  assign n23661 = n35322 & n22861 ;
  assign n20039 = n67 & n34367 ;
  assign n23662 = x8 & n20039 ;
  assign n20178 = n7068 & n20170 ;
  assign n23663 = n7017 & n34350 ;
  assign n23664 = n69 & n34367 ;
  assign n23665 = n23663 | n23664 ;
  assign n23666 = n20178 | n23665 ;
  assign n23668 = n23662 | n23666 ;
  assign n23669 = x8 & n23668 ;
  assign n20014 = n7017 & n19991 ;
  assign n23670 = n69 & n34350 ;
  assign n23671 = n7041 & n34367 ;
  assign n23672 = n23670 | n23671 ;
  assign n23673 = n20014 | n23672 ;
  assign n23674 = n7068 & n20189 ;
  assign n23675 = n23673 | n23674 ;
  assign n23677 = n23669 | n23675 ;
  assign n35323 = ~n23677 ;
  assign n23678 = x8 & n35323 ;
  assign n23680 = n20041 | n23678 ;
  assign n20209 = n7068 & n20207 ;
  assign n19993 = n69 & n19991 ;
  assign n20034 = n7041 & n34350 ;
  assign n23681 = n19993 | n20034 ;
  assign n23682 = n7017 & n34372 ;
  assign n23683 = n23681 | n23682 ;
  assign n23684 = n20209 | n23683 ;
  assign n35324 = ~n23684 ;
  assign n23685 = x8 & n35324 ;
  assign n23686 = n30185 & n23684 ;
  assign n23687 = n23685 | n23686 ;
  assign n23688 = n23680 & n23687 ;
  assign n23689 = x11 & n20041 ;
  assign n23690 = n22851 | n23689 ;
  assign n23691 = n22851 & n23689 ;
  assign n35325 = ~n23691 ;
  assign n23692 = n23690 & n35325 ;
  assign n23694 = n23688 | n23692 ;
  assign n23693 = n23688 & n23692 ;
  assign n35326 = ~n23693 ;
  assign n23695 = n35326 & n23694 ;
  assign n20284 = n7068 & n34383 ;
  assign n19984 = n69 & n34372 ;
  assign n19992 = n7041 & n19991 ;
  assign n23696 = n19984 | n19992 ;
  assign n23697 = n7017 & n34381 ;
  assign n23698 = n23696 | n23697 ;
  assign n23699 = n20284 | n23698 ;
  assign n35327 = ~n23699 ;
  assign n23700 = x8 & n35327 ;
  assign n23701 = n30185 & n23699 ;
  assign n23702 = n23700 | n23701 ;
  assign n35328 = ~n23702 ;
  assign n23703 = n23695 & n35328 ;
  assign n35329 = ~n23703 ;
  assign n23704 = n23694 & n35329 ;
  assign n23706 = n23661 | n23704 ;
  assign n20421 = n7068 & n20412 ;
  assign n19949 = n69 & n34381 ;
  assign n19974 = n7041 & n34372 ;
  assign n23707 = n19949 | n19974 ;
  assign n23708 = n7017 & n19917 ;
  assign n23709 = n23707 | n23708 ;
  assign n23710 = n20421 | n23709 ;
  assign n35330 = ~n23710 ;
  assign n23711 = x8 & n35330 ;
  assign n23712 = n30185 & n23710 ;
  assign n23713 = n23711 | n23712 ;
  assign n23705 = n23661 & n23704 ;
  assign n35331 = ~n23705 ;
  assign n23714 = n35331 & n23706 ;
  assign n35332 = ~n23713 ;
  assign n23715 = n35332 & n23714 ;
  assign n35333 = ~n23715 ;
  assign n23716 = n23706 & n35333 ;
  assign n23718 = n23660 | n23716 ;
  assign n20351 = n7068 & n34399 ;
  assign n19936 = n69 & n19917 ;
  assign n19957 = n7041 & n34381 ;
  assign n23719 = n19936 | n19957 ;
  assign n23720 = n7017 & n19893 ;
  assign n23721 = n23719 | n23720 ;
  assign n23722 = n20351 | n23721 ;
  assign n23723 = x8 | n23722 ;
  assign n23724 = x8 & n23722 ;
  assign n35334 = ~n23724 ;
  assign n23725 = n23723 & n35334 ;
  assign n23717 = n23660 & n23716 ;
  assign n35335 = ~n23717 ;
  assign n23726 = n35335 & n23718 ;
  assign n35336 = ~n23725 ;
  assign n23727 = n35336 & n23726 ;
  assign n35337 = ~n23727 ;
  assign n23729 = n23718 & n35337 ;
  assign n35338 = ~n23729 ;
  assign n23731 = n23655 & n35338 ;
  assign n35339 = ~n23731 ;
  assign n23732 = n23654 & n35339 ;
  assign n35340 = ~n23732 ;
  assign n23734 = n23643 & n35340 ;
  assign n35341 = ~n23734 ;
  assign n23735 = n23642 & n35341 ;
  assign n35342 = ~n23735 ;
  assign n23737 = n23631 & n35342 ;
  assign n35343 = ~n23737 ;
  assign n23738 = n23629 & n35343 ;
  assign n35344 = ~n23738 ;
  assign n23740 = n23618 & n35344 ;
  assign n35345 = ~n23740 ;
  assign n23741 = n23617 & n35345 ;
  assign n35346 = ~n23741 ;
  assign n23742 = n23606 & n35346 ;
  assign n35347 = ~n23742 ;
  assign n23743 = n23604 & n35347 ;
  assign n35348 = ~n23743 ;
  assign n23745 = n23593 & n35348 ;
  assign n35349 = ~n23745 ;
  assign n23746 = n23592 & n35349 ;
  assign n35350 = ~n23746 ;
  assign n23747 = n23581 & n35350 ;
  assign n35351 = ~n23747 ;
  assign n23748 = n23580 & n35351 ;
  assign n23749 = n23569 & n23748 ;
  assign n22930 = n22798 | n22929 ;
  assign n23750 = n22798 & n22929 ;
  assign n35352 = ~n23750 ;
  assign n23751 = n22930 & n35352 ;
  assign n23752 = n23569 | n23748 ;
  assign n35353 = ~n23749 ;
  assign n23753 = n35353 & n23752 ;
  assign n23754 = n23751 & n23753 ;
  assign n23755 = n23749 | n23754 ;
  assign n35354 = ~n23755 ;
  assign n23757 = n23562 & n35354 ;
  assign n35355 = ~n23757 ;
  assign n23758 = n23560 & n35355 ;
  assign n35356 = ~n23540 ;
  assign n23548 = n35356 & n23547 ;
  assign n35357 = ~n23547 ;
  assign n23759 = n23540 & n35357 ;
  assign n23760 = n23548 | n23759 ;
  assign n35358 = ~n23758 ;
  assign n23761 = n35358 & n23760 ;
  assign n35359 = ~n23761 ;
  assign n23762 = n23549 & n35359 ;
  assign n23764 = n23539 & n23762 ;
  assign n23765 = n23537 | n23764 ;
  assign n23766 = n23523 & n23525 ;
  assign n23767 = n23765 | n23766 ;
  assign n23768 = n23526 & n23767 ;
  assign n35360 = ~n23768 ;
  assign n23769 = n23516 & n35360 ;
  assign n35361 = ~n23769 ;
  assign n23770 = n23514 & n35361 ;
  assign n35362 = ~n23770 ;
  assign n23772 = n23504 & n35362 ;
  assign n35363 = ~n23772 ;
  assign n23773 = n23503 & n35363 ;
  assign n23491 = n23483 & n23490 ;
  assign n35364 = ~n23491 ;
  assign n23774 = n35364 & n23492 ;
  assign n35365 = ~n23773 ;
  assign n23775 = n35365 & n23774 ;
  assign n35366 = ~n23775 ;
  assign n23776 = n23492 & n35366 ;
  assign n23777 = n23481 & n23776 ;
  assign n35367 = ~n22701 ;
  assign n23778 = n35367 & n22953 ;
  assign n23779 = n22954 | n23778 ;
  assign n23780 = n23481 | n23776 ;
  assign n35368 = ~n23777 ;
  assign n23781 = n35368 & n23780 ;
  assign n23782 = n23779 & n23781 ;
  assign n23783 = n23777 | n23782 ;
  assign n35369 = ~n23783 ;
  assign n23784 = n23474 & n35369 ;
  assign n35370 = ~n23784 ;
  assign n23785 = n23472 & n35370 ;
  assign n23787 = n23461 | n23785 ;
  assign n35371 = ~n22677 ;
  assign n23788 = n35371 & n22958 ;
  assign n23789 = n22959 | n23788 ;
  assign n23786 = n23461 & n23785 ;
  assign n35372 = ~n23786 ;
  assign n23790 = n35372 & n23787 ;
  assign n35373 = ~n23789 ;
  assign n23791 = n35373 & n23790 ;
  assign n35374 = ~n23791 ;
  assign n23792 = n23787 & n35374 ;
  assign n23794 = n23454 | n23792 ;
  assign n35375 = ~n23453 ;
  assign n23795 = n35375 & n23794 ;
  assign n23796 = n23425 | n23795 ;
  assign n35376 = ~n23423 ;
  assign n23797 = n35376 & n23796 ;
  assign n23798 = n23395 & n23797 ;
  assign n23799 = n23395 | n23797 ;
  assign n35377 = ~n23798 ;
  assign n23800 = n35377 & n23799 ;
  assign n23801 = n140 | n1047 ;
  assign n23802 = n2940 | n2955 ;
  assign n23803 = n23801 | n23802 ;
  assign n23804 = n5100 | n23803 ;
  assign n23805 = n1126 | n2231 ;
  assign n23806 = n11572 | n23805 ;
  assign n23807 = n23804 | n23806 ;
  assign n23808 = n771 | n3141 ;
  assign n23809 = n22203 | n23808 ;
  assign n23810 = n1196 | n23809 ;
  assign n23811 = n23807 | n23810 ;
  assign n23812 = n324 | n346 ;
  assign n23813 = n383 | n795 ;
  assign n23814 = n23812 | n23813 ;
  assign n23815 = n533 | n677 ;
  assign n23816 = n23814 | n23815 ;
  assign n23817 = n1641 | n3682 ;
  assign n23818 = n23816 | n23817 ;
  assign n23819 = n2659 | n2749 ;
  assign n23820 = n3075 | n23819 ;
  assign n23821 = n854 | n23820 ;
  assign n23822 = n23818 | n23821 ;
  assign n23823 = n3725 | n23822 ;
  assign n23824 = n2545 | n23823 ;
  assign n23825 = n23811 | n23824 ;
  assign n35378 = ~n23825 ;
  assign n23826 = n1603 & n35378 ;
  assign n23827 = n23238 & n23826 ;
  assign n23828 = n23238 | n23826 ;
  assign n35379 = ~n23827 ;
  assign n23829 = n35379 & n23828 ;
  assign n23830 = n23118 & n23829 ;
  assign n23831 = n23118 | n23829 ;
  assign n35380 = ~n23830 ;
  assign n23832 = n35380 & n23831 ;
  assign n14192 = n889 & n14183 ;
  assign n14142 = n3329 & n14124 ;
  assign n14169 = n3311 & n14147 ;
  assign n23833 = n14142 | n14169 ;
  assign n23834 = n3343 & n14196 ;
  assign n23835 = n23833 | n23834 ;
  assign n23836 = n14192 | n23835 ;
  assign n23837 = n23832 | n23836 ;
  assign n23838 = n23832 & n23836 ;
  assign n35381 = ~n23838 ;
  assign n23839 = n23837 & n35381 ;
  assign n23193 = n23186 | n23191 ;
  assign n35382 = ~n23185 ;
  assign n23840 = n35382 & n23193 ;
  assign n35383 = ~n23839 ;
  assign n23841 = n35383 & n23840 ;
  assign n35384 = ~n23840 ;
  assign n23842 = n23839 & n35384 ;
  assign n23843 = n23841 | n23842 ;
  assign n14576 = n895 & n14570 ;
  assign n14532 = n2849 & n32706 ;
  assign n14555 = n2861 & n14536 ;
  assign n23844 = n14532 | n14555 ;
  assign n23845 = n894 & n32707 ;
  assign n23846 = n23844 | n23845 ;
  assign n23847 = n14576 | n23846 ;
  assign n35385 = ~n23847 ;
  assign n23848 = x29 & n35385 ;
  assign n23849 = n30024 & n23847 ;
  assign n23850 = n23848 | n23849 ;
  assign n35386 = ~n23850 ;
  assign n23851 = n23843 & n35386 ;
  assign n35387 = ~n23843 ;
  assign n23852 = n35387 & n23850 ;
  assign n23853 = n23851 | n23852 ;
  assign n23854 = n23198 | n23199 ;
  assign n35388 = ~n23197 ;
  assign n23855 = n35388 & n23854 ;
  assign n35389 = ~n23853 ;
  assign n23856 = n35389 & n23855 ;
  assign n35390 = ~n23855 ;
  assign n23857 = n23853 & n35390 ;
  assign n23858 = n23856 | n23857 ;
  assign n15189 = n3791 & n32875 ;
  assign n15076 = n3802 & n32856 ;
  assign n15097 = n209 & n15081 ;
  assign n23859 = n15076 | n15097 ;
  assign n23860 = n3818 & n32876 ;
  assign n23861 = n23859 | n23860 ;
  assign n23862 = n15189 | n23861 ;
  assign n23863 = x26 | n23862 ;
  assign n23864 = x26 & n23862 ;
  assign n35391 = ~n23864 ;
  assign n23865 = n23863 & n35391 ;
  assign n35392 = ~n23865 ;
  assign n23867 = n23858 & n35392 ;
  assign n23866 = n23858 & n23865 ;
  assign n23868 = n23858 | n23865 ;
  assign n35393 = ~n23866 ;
  assign n23869 = n35393 & n23868 ;
  assign n35394 = ~n23209 ;
  assign n23870 = n23202 & n35394 ;
  assign n23871 = n23212 | n23219 ;
  assign n35395 = ~n23870 ;
  assign n23872 = n35395 & n23871 ;
  assign n23874 = n23869 | n23872 ;
  assign n35396 = ~n23867 ;
  assign n23875 = n35396 & n23874 ;
  assign n4184 = x23 & n4183 ;
  assign n15241 = x22 & n15221 ;
  assign n23876 = x23 & n32883 ;
  assign n23877 = n4183 | n23876 ;
  assign n23878 = n15241 | n23877 ;
  assign n35397 = ~n4184 ;
  assign n23879 = n35397 & n23878 ;
  assign n23880 = n23875 & n23879 ;
  assign n35398 = ~n23836 ;
  assign n23881 = n23832 & n35398 ;
  assign n23882 = n23839 | n23840 ;
  assign n35399 = ~n23881 ;
  assign n23883 = n35399 & n23882 ;
  assign n23884 = n35193 & n23829 ;
  assign n35400 = ~n23884 ;
  assign n23885 = n23828 & n35400 ;
  assign n23886 = n131 | n621 ;
  assign n23887 = n2573 | n23886 ;
  assign n23888 = n348 | n433 ;
  assign n23889 = n660 | n750 ;
  assign n23890 = n23888 | n23889 ;
  assign n23891 = n2169 | n23890 ;
  assign n23892 = n2430 | n3187 ;
  assign n23893 = n23891 | n23892 ;
  assign n23894 = n23887 | n23893 ;
  assign n23895 = n181 | n318 ;
  assign n23896 = n564 | n23895 ;
  assign n23897 = n698 | n808 ;
  assign n23898 = n11607 | n23897 ;
  assign n23899 = n23896 | n23898 ;
  assign n23900 = n2528 | n23899 ;
  assign n23901 = n23894 | n23900 ;
  assign n23902 = n1377 | n23901 ;
  assign n23903 = n14002 | n23902 ;
  assign n35401 = ~n23903 ;
  assign n23904 = n23885 & n35401 ;
  assign n35402 = ~n23885 ;
  assign n23905 = n35402 & n23903 ;
  assign n23906 = n23904 | n23905 ;
  assign n14976 = n889 & n14965 ;
  assign n14121 = n3329 & n14101 ;
  assign n14145 = n3311 & n14124 ;
  assign n23907 = n14121 | n14145 ;
  assign n23908 = n3343 & n14536 ;
  assign n23909 = n23907 | n23908 ;
  assign n23910 = n14976 | n23909 ;
  assign n23911 = n23906 | n23910 ;
  assign n23912 = n23906 & n23910 ;
  assign n35403 = ~n23912 ;
  assign n23913 = n23911 & n35403 ;
  assign n23914 = n23883 & n23913 ;
  assign n23915 = n23883 | n23913 ;
  assign n35404 = ~n23914 ;
  assign n23916 = n35404 & n23915 ;
  assign n15297 = n895 & n15288 ;
  assign n14497 = n2849 & n32707 ;
  assign n14528 = n2861 & n32706 ;
  assign n23917 = n14497 | n14528 ;
  assign n23918 = n894 & n15081 ;
  assign n23919 = n23917 | n23918 ;
  assign n23920 = n15297 | n23919 ;
  assign n35405 = ~n23920 ;
  assign n23921 = x29 & n35405 ;
  assign n23922 = n30024 & n23920 ;
  assign n23923 = n23921 | n23922 ;
  assign n35406 = ~n23923 ;
  assign n23924 = n23916 & n35406 ;
  assign n35407 = ~n23916 ;
  assign n23925 = n35407 & n23923 ;
  assign n23926 = n23924 | n23925 ;
  assign n23927 = n23853 | n23855 ;
  assign n35408 = ~n23851 ;
  assign n23928 = n35408 & n23927 ;
  assign n35409 = ~n23926 ;
  assign n23929 = n35409 & n23928 ;
  assign n35410 = ~n23928 ;
  assign n23930 = n23926 & n35410 ;
  assign n23931 = n23929 | n23930 ;
  assign n15271 = n3791 & n32889 ;
  assign n15066 = n209 & n32856 ;
  assign n15174 = n3802 & n32876 ;
  assign n23932 = n15066 | n15174 ;
  assign n23933 = n3818 & n32890 ;
  assign n23934 = n23932 | n23933 ;
  assign n23935 = n15271 | n23934 ;
  assign n35411 = ~n23935 ;
  assign n23936 = x26 & n35411 ;
  assign n23937 = n30019 & n23935 ;
  assign n23938 = n23936 | n23937 ;
  assign n35412 = ~n23938 ;
  assign n23939 = n23931 & n35412 ;
  assign n35413 = ~n23931 ;
  assign n23940 = n35413 & n23938 ;
  assign n23941 = n23939 | n23940 ;
  assign n23942 = n23875 | n23879 ;
  assign n35414 = ~n23880 ;
  assign n23943 = n35414 & n23942 ;
  assign n23945 = n23941 & n23943 ;
  assign n23946 = n23880 | n23945 ;
  assign n23947 = n869 | n2252 ;
  assign n23948 = n21355 | n23947 ;
  assign n23949 = n326 | n331 ;
  assign n23950 = n661 | n23949 ;
  assign n23951 = n11226 | n23950 ;
  assign n23952 = n23948 | n23951 ;
  assign n23953 = n238 | n4995 ;
  assign n23954 = n23952 | n23953 ;
  assign n23955 = n658 | n767 ;
  assign n23956 = n755 | n23955 ;
  assign n23957 = n2951 | n4804 ;
  assign n23958 = n23956 | n23957 ;
  assign n23959 = n1066 | n23958 ;
  assign n23960 = n3112 | n3453 ;
  assign n23961 = n5032 | n13889 ;
  assign n23962 = n23960 | n23961 ;
  assign n23963 = n23959 | n23962 ;
  assign n23964 = n23954 | n23963 ;
  assign n23965 = n11115 | n23964 ;
  assign n23966 = n23094 | n23965 ;
  assign n23967 = n23903 | n23966 ;
  assign n23968 = n23903 & n23966 ;
  assign n35415 = ~n23968 ;
  assign n23969 = n23967 & n35415 ;
  assign n23970 = n23885 | n23903 ;
  assign n23971 = n35403 & n23970 ;
  assign n35416 = ~n23969 ;
  assign n23972 = n35416 & n23971 ;
  assign n35417 = ~n23971 ;
  assign n23973 = n23969 & n35417 ;
  assign n23974 = n23972 | n23973 ;
  assign n14692 = n889 & n32735 ;
  assign n14122 = n3311 & n14101 ;
  assign n14556 = n3329 & n14536 ;
  assign n23975 = n14122 | n14556 ;
  assign n23976 = n3343 & n32706 ;
  assign n23977 = n23975 | n23976 ;
  assign n23978 = n14692 | n23977 ;
  assign n23979 = n23974 | n23978 ;
  assign n23980 = n23974 & n23978 ;
  assign n35418 = ~n23980 ;
  assign n23981 = n23979 & n35418 ;
  assign n15113 = n895 & n15111 ;
  assign n14501 = n2861 & n32707 ;
  assign n15104 = n2849 & n15081 ;
  assign n23982 = n14501 | n15104 ;
  assign n23983 = n894 & n32856 ;
  assign n23984 = n23982 | n23983 ;
  assign n23985 = n15113 | n23984 ;
  assign n35419 = ~n23985 ;
  assign n23986 = x29 & n35419 ;
  assign n23987 = n30024 & n23985 ;
  assign n23988 = n23986 | n23987 ;
  assign n35420 = ~n23988 ;
  assign n23989 = n23981 & n35420 ;
  assign n35421 = ~n23981 ;
  assign n23990 = n35421 & n23988 ;
  assign n23991 = n23989 | n23990 ;
  assign n15529 = n3791 & n15526 ;
  assign n15178 = n209 & n32876 ;
  assign n15245 = n3818 & n15221 ;
  assign n23992 = n15178 | n15245 ;
  assign n23993 = n3802 & n32890 ;
  assign n23994 = n23992 | n23993 ;
  assign n23995 = n15529 | n23994 ;
  assign n23996 = x26 | n23995 ;
  assign n23997 = x26 & n23995 ;
  assign n35422 = ~n23997 ;
  assign n23998 = n23996 & n35422 ;
  assign n35423 = ~n23924 ;
  assign n23999 = n23915 & n35423 ;
  assign n24000 = n23998 & n23999 ;
  assign n24001 = n23998 | n23999 ;
  assign n35424 = ~n24000 ;
  assign n24002 = n35424 & n24001 ;
  assign n24003 = n23991 & n24002 ;
  assign n24004 = n23991 | n24002 ;
  assign n35425 = ~n24003 ;
  assign n24005 = n35425 & n24004 ;
  assign n4131 = x22 | n4129 ;
  assign n24006 = n4131 & n35397 ;
  assign n24007 = n23926 | n23928 ;
  assign n35426 = ~n23939 ;
  assign n24008 = n35426 & n24007 ;
  assign n24009 = n24006 & n24008 ;
  assign n24010 = n24006 | n24008 ;
  assign n35427 = ~n24009 ;
  assign n24011 = n35427 & n24010 ;
  assign n35428 = ~n24005 ;
  assign n24012 = n35428 & n24011 ;
  assign n35429 = ~n24011 ;
  assign n24013 = n24005 & n35429 ;
  assign n24014 = n24012 | n24013 ;
  assign n24015 = n23946 | n24014 ;
  assign n24016 = n23946 & n24014 ;
  assign n35430 = ~n24016 ;
  assign n24017 = n24015 & n35430 ;
  assign n35431 = ~n23941 ;
  assign n23944 = n35431 & n23943 ;
  assign n35432 = ~n23943 ;
  assign n24018 = n23941 & n35432 ;
  assign n24019 = n23944 | n24018 ;
  assign n15520 = n4132 & n15516 ;
  assign n15244 = n4148 & n15221 ;
  assign n24020 = n4165 | n15244 ;
  assign n24021 = n4185 & n32890 ;
  assign n24022 = n24020 | n24021 ;
  assign n24023 = n15520 | n24022 ;
  assign n24024 = x23 | n24023 ;
  assign n24025 = x23 & n24023 ;
  assign n35433 = ~n24025 ;
  assign n24026 = n24024 & n35433 ;
  assign n24027 = n23232 | n23235 ;
  assign n24029 = n24026 & n24027 ;
  assign n35434 = ~n23869 ;
  assign n23873 = n35434 & n23872 ;
  assign n35435 = ~n23872 ;
  assign n24030 = n23869 & n35435 ;
  assign n24031 = n23873 | n24030 ;
  assign n35436 = ~n24027 ;
  assign n24028 = n24026 & n35436 ;
  assign n35437 = ~n24026 ;
  assign n24032 = n35437 & n24027 ;
  assign n24033 = n24028 | n24032 ;
  assign n35438 = ~n24031 ;
  assign n24034 = n35438 & n24033 ;
  assign n24036 = n24029 | n24034 ;
  assign n24038 = n24019 | n24036 ;
  assign n35439 = ~n24036 ;
  assign n24037 = n24019 & n35439 ;
  assign n35440 = ~n24019 ;
  assign n24039 = n35440 & n24036 ;
  assign n24040 = n24037 | n24039 ;
  assign n24035 = n24031 & n24033 ;
  assign n24041 = n24031 | n24033 ;
  assign n35441 = ~n24035 ;
  assign n24042 = n35441 & n24041 ;
  assign n24043 = n23242 & n35216 ;
  assign n35442 = ~n24043 ;
  assign n24045 = n24042 & n35442 ;
  assign n35443 = ~n24042 ;
  assign n24044 = n35443 & n24043 ;
  assign n24046 = n24044 | n24045 ;
  assign n35444 = ~n23247 ;
  assign n24047 = n35444 & n23384 ;
  assign n24050 = n24046 | n24047 ;
  assign n35445 = ~n24045 ;
  assign n24051 = n35445 & n24050 ;
  assign n35446 = ~n24051 ;
  assign n24052 = n24040 & n35446 ;
  assign n35447 = ~n24052 ;
  assign n24053 = n24038 & n35447 ;
  assign n24054 = n24017 & n24053 ;
  assign n24056 = n24017 | n24053 ;
  assign n35448 = ~n24054 ;
  assign n24057 = n35448 & n24056 ;
  assign n35449 = ~n24040 ;
  assign n24079 = n35449 & n24051 ;
  assign n24080 = n24052 | n24079 ;
  assign n35450 = ~n24046 ;
  assign n24048 = n35450 & n24047 ;
  assign n35451 = ~n24047 ;
  assign n24102 = n24046 & n35451 ;
  assign n24103 = n24048 | n24102 ;
  assign n35452 = ~n23364 ;
  assign n24126 = n23316 & n35452 ;
  assign n24128 = n23290 | n24126 ;
  assign n24129 = n24103 & n24128 ;
  assign n24130 = n24080 & n24129 ;
  assign n24131 = n35244 & n23366 ;
  assign n35453 = ~n24131 ;
  assign n24132 = n23290 & n35453 ;
  assign n24133 = n24103 | n24132 ;
  assign n24134 = n24080 | n24133 ;
  assign n35454 = ~n24130 ;
  assign n24135 = n35454 & n24134 ;
  assign n35455 = ~n24135 ;
  assign n24136 = n24057 & n35455 ;
  assign n35456 = ~n24057 ;
  assign n24137 = n35456 & n24135 ;
  assign n24138 = n24136 | n24137 ;
  assign n35457 = ~n24138 ;
  assign n24139 = n8157 & n35457 ;
  assign n24094 = n740 & n24080 ;
  assign n35458 = ~n24103 ;
  assign n24112 = n8195 & n35458 ;
  assign n24152 = n24094 | n24112 ;
  assign n35459 = ~n24017 ;
  assign n24055 = n35459 & n24053 ;
  assign n35460 = ~n24053 ;
  assign n24150 = n24017 & n35460 ;
  assign n24151 = n24055 | n24150 ;
  assign n24153 = n9052 & n24151 ;
  assign n24154 = n24152 | n24153 ;
  assign n24155 = n24139 | n24154 ;
  assign n24156 = x5 | n24155 ;
  assign n24157 = x5 & n24155 ;
  assign n35461 = ~n24157 ;
  assign n24158 = n24156 & n35461 ;
  assign n24159 = n23800 & n24158 ;
  assign n24160 = n23800 | n24158 ;
  assign n35462 = ~n24159 ;
  assign n24161 = n35462 & n24160 ;
  assign n24049 = n24046 & n24047 ;
  assign n35463 = ~n24049 ;
  assign n24162 = n35463 & n24050 ;
  assign n35464 = ~n24128 ;
  assign n24163 = n35464 & n24162 ;
  assign n35465 = ~n24162 ;
  assign n24164 = n24132 & n35465 ;
  assign n24165 = n24163 | n24164 ;
  assign n24166 = n24080 & n24165 ;
  assign n24167 = n24080 | n24165 ;
  assign n35466 = ~n24166 ;
  assign n24168 = n35466 & n24167 ;
  assign n24169 = n8157 & n24168 ;
  assign n35467 = ~n23290 ;
  assign n23304 = n8195 & n35467 ;
  assign n24116 = n740 & n35458 ;
  assign n24180 = n23304 | n24116 ;
  assign n24181 = n9052 & n24080 ;
  assign n24182 = n24180 | n24181 ;
  assign n24183 = n24169 | n24182 ;
  assign n35468 = ~n24183 ;
  assign n24184 = x5 & n35468 ;
  assign n24185 = n30053 & n24183 ;
  assign n24186 = n24184 | n24185 ;
  assign n35469 = ~n23454 ;
  assign n23793 = n35469 & n23792 ;
  assign n35470 = ~n23792 ;
  assign n24187 = n23454 & n35470 ;
  assign n24188 = n23793 | n24187 ;
  assign n24127 = n35467 & n24126 ;
  assign n24189 = n23290 & n24131 ;
  assign n24190 = n24127 | n24189 ;
  assign n24191 = n35458 & n24190 ;
  assign n35471 = ~n24190 ;
  assign n24192 = n24103 & n35471 ;
  assign n24193 = n24191 | n24192 ;
  assign n35472 = ~n24193 ;
  assign n24194 = n8157 & n35472 ;
  assign n23297 = n740 & n35467 ;
  assign n23321 = n8195 & n35244 ;
  assign n24205 = n23297 | n23321 ;
  assign n24206 = n9052 & n35465 ;
  assign n24207 = n24205 | n24206 ;
  assign n24208 = n24194 | n24207 ;
  assign n24209 = x5 | n24208 ;
  assign n24210 = x5 & n24208 ;
  assign n35473 = ~n24210 ;
  assign n24211 = n24209 & n35473 ;
  assign n35474 = ~n24211 ;
  assign n24213 = n24188 & n35474 ;
  assign n35475 = ~n24188 ;
  assign n24212 = n35475 & n24211 ;
  assign n24214 = n24212 | n24213 ;
  assign n35476 = ~n23790 ;
  assign n24215 = n23789 & n35476 ;
  assign n24216 = n23791 | n24215 ;
  assign n23374 = n8157 & n23372 ;
  assign n23327 = n740 & n35244 ;
  assign n23349 = n8195 & n23339 ;
  assign n24217 = n23327 | n23349 ;
  assign n24218 = n9052 & n35246 ;
  assign n24219 = n24217 | n24218 ;
  assign n24220 = n23374 | n24219 ;
  assign n24221 = x5 | n24220 ;
  assign n24222 = x5 & n24220 ;
  assign n35477 = ~n24222 ;
  assign n24223 = n24221 & n35477 ;
  assign n24225 = n24216 | n24223 ;
  assign n35478 = ~n24216 ;
  assign n24224 = n35478 & n24223 ;
  assign n35479 = ~n24223 ;
  assign n24226 = n24216 & n35479 ;
  assign n24227 = n24224 | n24226 ;
  assign n35480 = ~n23474 ;
  assign n24228 = n35480 & n23783 ;
  assign n24229 = n23784 | n24228 ;
  assign n23405 = n8157 & n35252 ;
  assign n22521 = n8195 & n35020 ;
  assign n23341 = n740 & n23339 ;
  assign n24230 = n22521 | n23341 ;
  assign n24231 = n9052 & n35254 ;
  assign n24232 = n24230 | n24231 ;
  assign n24233 = n23405 | n24232 ;
  assign n24234 = x5 | n24233 ;
  assign n24235 = x5 & n24233 ;
  assign n35481 = ~n24235 ;
  assign n24236 = n24234 & n35481 ;
  assign n24237 = n24229 & n24236 ;
  assign n24238 = n23779 | n23781 ;
  assign n35482 = ~n23782 ;
  assign n24239 = n35482 & n24238 ;
  assign n23436 = n8157 & n35262 ;
  assign n22518 = n740 & n35020 ;
  assign n22585 = n8195 & n22533 ;
  assign n24240 = n22518 | n22585 ;
  assign n24241 = n9052 & n23444 ;
  assign n24242 = n24240 | n24241 ;
  assign n24243 = n23436 | n24242 ;
  assign n24244 = x5 | n24243 ;
  assign n24245 = x5 & n24243 ;
  assign n35483 = ~n24245 ;
  assign n24246 = n24244 & n35483 ;
  assign n24248 = n24239 | n24246 ;
  assign n35484 = ~n23774 ;
  assign n24249 = n23773 & n35484 ;
  assign n24250 = n23775 | n24249 ;
  assign n22569 = n8157 & n35022 ;
  assign n22540 = n8195 & n35018 ;
  assign n22590 = n740 & n22533 ;
  assign n24251 = n22540 | n22590 ;
  assign n24252 = n9052 & n35020 ;
  assign n24253 = n24251 | n24252 ;
  assign n24254 = n22569 | n24253 ;
  assign n24255 = x5 | n24254 ;
  assign n24256 = x5 & n24254 ;
  assign n35485 = ~n24256 ;
  assign n24257 = n24255 & n35485 ;
  assign n24259 = n24250 | n24257 ;
  assign n24258 = n24250 & n24257 ;
  assign n35486 = ~n24258 ;
  assign n24260 = n35486 & n24259 ;
  assign n35487 = ~n23504 ;
  assign n23771 = n35487 & n23770 ;
  assign n24261 = n23771 | n23772 ;
  assign n22625 = n8157 & n35030 ;
  assign n21740 = n8195 & n21729 ;
  assign n22539 = n740 & n35018 ;
  assign n24262 = n21740 | n22539 ;
  assign n24263 = n9052 & n22533 ;
  assign n24264 = n24262 | n24263 ;
  assign n24265 = n22625 | n24264 ;
  assign n24266 = x5 | n24265 ;
  assign n24267 = x5 & n24265 ;
  assign n35488 = ~n24267 ;
  assign n24268 = n24266 & n35488 ;
  assign n24270 = n24261 | n24268 ;
  assign n35489 = ~n24261 ;
  assign n24269 = n35489 & n24268 ;
  assign n35490 = ~n24268 ;
  assign n24271 = n24261 & n35490 ;
  assign n24272 = n24269 | n24271 ;
  assign n22647 = n8157 & n35035 ;
  assign n21735 = n740 & n21729 ;
  assign n21812 = n8195 & n21753 ;
  assign n24273 = n21735 | n21812 ;
  assign n24274 = n9052 & n35018 ;
  assign n24275 = n24273 | n24274 ;
  assign n24276 = n22647 | n24275 ;
  assign n24277 = x5 | n24276 ;
  assign n24278 = x5 & n24276 ;
  assign n35491 = ~n24278 ;
  assign n24279 = n24277 & n35491 ;
  assign n35492 = ~n23766 ;
  assign n24280 = n23526 & n35492 ;
  assign n24281 = n23765 & n24280 ;
  assign n24282 = n23765 | n24280 ;
  assign n35493 = ~n24281 ;
  assign n24283 = n35493 & n24282 ;
  assign n21795 = n8157 & n34802 ;
  assign n21757 = n8195 & n34803 ;
  assign n21810 = n740 & n21753 ;
  assign n24284 = n21757 | n21810 ;
  assign n24285 = n9052 & n21804 ;
  assign n24286 = n24284 | n24285 ;
  assign n24287 = n21795 | n24286 ;
  assign n24288 = x5 | n24287 ;
  assign n24289 = x5 & n24287 ;
  assign n35494 = ~n24289 ;
  assign n24290 = n24288 & n35494 ;
  assign n24292 = n24283 | n24290 ;
  assign n21854 = n8157 & n21848 ;
  assign n19660 = n8195 & n34360 ;
  assign n21756 = n740 & n34803 ;
  assign n24293 = n19660 | n21756 ;
  assign n24294 = n9052 & n21753 ;
  assign n24295 = n24293 | n24294 ;
  assign n24296 = n21854 | n24295 ;
  assign n35495 = ~n24296 ;
  assign n24297 = x5 & n35495 ;
  assign n24298 = n30053 & n24296 ;
  assign n24299 = n24297 | n24298 ;
  assign n35496 = ~n23760 ;
  assign n24300 = n23758 & n35496 ;
  assign n24301 = n23761 | n24300 ;
  assign n21876 = n8157 & n34817 ;
  assign n19662 = n740 & n34360 ;
  assign n19685 = n8195 & n34349 ;
  assign n24302 = n19662 | n19685 ;
  assign n24303 = n9052 & n34803 ;
  assign n24304 = n24302 | n24303 ;
  assign n24305 = n21876 | n24304 ;
  assign n24306 = x5 | n24305 ;
  assign n24307 = x5 & n24305 ;
  assign n35497 = ~n24307 ;
  assign n24308 = n24306 & n35497 ;
  assign n24309 = n24301 & n24308 ;
  assign n24310 = n24301 | n24308 ;
  assign n20153 = n8157 & n34362 ;
  assign n19693 = n740 & n34349 ;
  assign n19712 = n8195 & n34363 ;
  assign n24311 = n19693 | n19712 ;
  assign n24312 = n9052 & n34365 ;
  assign n24313 = n24311 | n24312 ;
  assign n24314 = n20153 | n24313 ;
  assign n35498 = ~n24314 ;
  assign n24315 = x5 & n35498 ;
  assign n24316 = n30053 & n24314 ;
  assign n24317 = n24315 | n24316 ;
  assign n24318 = n23751 | n23753 ;
  assign n35499 = ~n23754 ;
  assign n24319 = n35499 & n24318 ;
  assign n21076 = n8157 & n34598 ;
  assign n19708 = n740 & n34363 ;
  assign n19730 = n8195 & n34520 ;
  assign n24320 = n19708 | n19730 ;
  assign n24321 = n9052 & n34349 ;
  assign n24322 = n24320 | n24321 ;
  assign n24323 = n21076 | n24322 ;
  assign n24324 = x5 | n24323 ;
  assign n24325 = x5 & n24323 ;
  assign n35500 = ~n24325 ;
  assign n24326 = n24324 & n35500 ;
  assign n24328 = n24319 | n24326 ;
  assign n24327 = n24319 & n24326 ;
  assign n35501 = ~n24327 ;
  assign n24329 = n35501 & n24328 ;
  assign n35502 = ~n23581 ;
  assign n24330 = n35502 & n23746 ;
  assign n24331 = n23747 | n24330 ;
  assign n21099 = n8157 & n34603 ;
  assign n19741 = n740 & n34520 ;
  assign n19753 = n8195 & n19752 ;
  assign n24332 = n19741 | n19753 ;
  assign n24333 = n9052 & n34596 ;
  assign n24334 = n24332 | n24333 ;
  assign n24335 = n21099 | n24334 ;
  assign n24336 = x5 | n24335 ;
  assign n24337 = x5 & n24335 ;
  assign n35503 = ~n24337 ;
  assign n24338 = n24336 & n35503 ;
  assign n24340 = n24331 | n24338 ;
  assign n35504 = ~n24331 ;
  assign n24339 = n35504 & n24338 ;
  assign n35505 = ~n24338 ;
  assign n24341 = n24331 & n35505 ;
  assign n24342 = n24339 | n24341 ;
  assign n35506 = ~n23593 ;
  assign n23744 = n35506 & n23743 ;
  assign n24343 = n23744 | n23745 ;
  assign n20812 = n8157 & n20805 ;
  assign n19758 = n740 & n19752 ;
  assign n19783 = n8195 & n34519 ;
  assign n24344 = n19758 | n19783 ;
  assign n24345 = n9052 & n34520 ;
  assign n24346 = n24344 | n24345 ;
  assign n24347 = n20812 | n24346 ;
  assign n24348 = x5 | n24347 ;
  assign n24349 = x5 & n24347 ;
  assign n35507 = ~n24349 ;
  assign n24350 = n24348 & n35507 ;
  assign n24351 = n24343 | n24350 ;
  assign n35508 = ~n23606 ;
  assign n24352 = n35508 & n23741 ;
  assign n24353 = n23742 | n24352 ;
  assign n20840 = n8157 & n20833 ;
  assign n19790 = n740 & n34519 ;
  assign n19801 = n8195 & n34355 ;
  assign n24354 = n19790 | n19801 ;
  assign n24355 = n9052 & n20845 ;
  assign n24356 = n24354 | n24355 ;
  assign n24357 = n20840 | n24356 ;
  assign n24358 = x5 | n24357 ;
  assign n24359 = x5 & n24357 ;
  assign n35509 = ~n24359 ;
  assign n24360 = n24358 & n35509 ;
  assign n24362 = n24353 & n24360 ;
  assign n35510 = ~n24353 ;
  assign n24361 = n35510 & n24360 ;
  assign n35511 = ~n24360 ;
  assign n24363 = n24353 & n35511 ;
  assign n24364 = n24361 | n24363 ;
  assign n35512 = ~n23618 ;
  assign n23739 = n35512 & n23738 ;
  assign n24365 = n23739 | n23740 ;
  assign n20870 = n8157 & n20863 ;
  assign n19811 = n740 & n34355 ;
  assign n19840 = n8195 & n19824 ;
  assign n24366 = n19811 | n19840 ;
  assign n24367 = n9052 & n34536 ;
  assign n24368 = n24366 | n24367 ;
  assign n24369 = n20870 | n24368 ;
  assign n24370 = x5 | n24369 ;
  assign n24371 = x5 & n24369 ;
  assign n35513 = ~n24371 ;
  assign n24372 = n24370 & n35513 ;
  assign n24373 = n24365 & n24372 ;
  assign n24374 = n24365 | n24372 ;
  assign n35514 = ~n24373 ;
  assign n24375 = n35514 & n24374 ;
  assign n35515 = ~n23631 ;
  assign n23736 = n35515 & n23735 ;
  assign n24376 = n23736 | n23737 ;
  assign n20782 = n8157 & n34511 ;
  assign n19827 = n740 & n19824 ;
  assign n20109 = n8195 & n34354 ;
  assign n24377 = n19827 | n20109 ;
  assign n24378 = n9052 & n34513 ;
  assign n24379 = n24377 | n24378 ;
  assign n24380 = n20782 | n24379 ;
  assign n24381 = x5 | n24380 ;
  assign n24382 = x5 & n24380 ;
  assign n35516 = ~n24382 ;
  assign n24383 = n24381 & n35516 ;
  assign n24384 = n24376 | n24383 ;
  assign n23733 = n23643 & n23732 ;
  assign n24385 = n23643 | n23732 ;
  assign n35517 = ~n23733 ;
  assign n24386 = n35517 & n24385 ;
  assign n20522 = n8157 & n34442 ;
  assign n20084 = n8195 & n20067 ;
  assign n20110 = n740 & n34354 ;
  assign n24387 = n20084 | n20110 ;
  assign n24388 = n9052 & n20527 ;
  assign n24389 = n24387 | n24388 ;
  assign n24390 = n20522 | n24389 ;
  assign n24391 = x5 | n24390 ;
  assign n24392 = x5 & n24390 ;
  assign n35518 = ~n24392 ;
  assign n24393 = n24391 & n35518 ;
  assign n24395 = n24386 | n24393 ;
  assign n35519 = ~n24386 ;
  assign n24394 = n35519 & n24393 ;
  assign n35520 = ~n24393 ;
  assign n24396 = n24386 & n35520 ;
  assign n24397 = n24394 | n24396 ;
  assign n23730 = n23655 & n23729 ;
  assign n24398 = n23655 | n23729 ;
  assign n35521 = ~n23730 ;
  assign n24399 = n35521 & n24398 ;
  assign n20552 = n8157 & n34450 ;
  assign n19858 = n8195 & n19846 ;
  assign n20085 = n740 & n20067 ;
  assign n24400 = n19858 | n20085 ;
  assign n24401 = n9052 & n34452 ;
  assign n24402 = n24400 | n24401 ;
  assign n24403 = n20552 | n24402 ;
  assign n24404 = x5 | n24403 ;
  assign n24405 = x5 & n24403 ;
  assign n35522 = ~n24405 ;
  assign n24406 = n24404 & n35522 ;
  assign n24408 = n24399 | n24406 ;
  assign n35523 = ~n24399 ;
  assign n24407 = n35523 & n24406 ;
  assign n35524 = ~n24406 ;
  assign n24409 = n24399 & n35524 ;
  assign n24410 = n24407 | n24409 ;
  assign n23728 = n23725 & n23726 ;
  assign n24411 = n23725 | n23726 ;
  assign n35525 = ~n23728 ;
  assign n24412 = n35525 & n24411 ;
  assign n20584 = n8157 & n20579 ;
  assign n19859 = n740 & n19846 ;
  assign n19889 = n8195 & n19870 ;
  assign n24413 = n19859 | n19889 ;
  assign n24414 = n9052 & n20067 ;
  assign n24415 = n24413 | n24414 ;
  assign n24416 = n20584 | n24415 ;
  assign n24417 = x5 | n24416 ;
  assign n24418 = x5 & n24416 ;
  assign n35526 = ~n24418 ;
  assign n24419 = n24417 & n35526 ;
  assign n24421 = n24412 | n24419 ;
  assign n24420 = n24412 & n24419 ;
  assign n35527 = ~n24420 ;
  assign n24422 = n35527 & n24421 ;
  assign n35528 = ~n23714 ;
  assign n24423 = n23713 & n35528 ;
  assign n24424 = n23715 | n24423 ;
  assign n20494 = n8157 & n20486 ;
  assign n19883 = n740 & n19870 ;
  assign n19908 = n8195 & n19893 ;
  assign n24425 = n19883 | n19908 ;
  assign n24426 = n9052 & n19846 ;
  assign n24427 = n24425 | n24426 ;
  assign n24428 = n20494 | n24427 ;
  assign n24429 = x5 | n24428 ;
  assign n24430 = x5 & n24428 ;
  assign n35529 = ~n24430 ;
  assign n24431 = n24429 & n35529 ;
  assign n24433 = n24424 | n24431 ;
  assign n24432 = n24424 & n24431 ;
  assign n35530 = ~n24432 ;
  assign n24434 = n35530 & n24433 ;
  assign n35531 = ~n23695 ;
  assign n24435 = n35531 & n23702 ;
  assign n24436 = n23703 | n24435 ;
  assign n20320 = n8157 & n20311 ;
  assign n19911 = n740 & n19893 ;
  assign n19938 = n8195 & n19917 ;
  assign n24437 = n19911 | n19938 ;
  assign n24438 = n9052 & n19870 ;
  assign n24439 = n24437 | n24438 ;
  assign n24440 = n20320 | n24439 ;
  assign n24441 = x5 | n24440 ;
  assign n24442 = x5 & n24440 ;
  assign n35532 = ~n24442 ;
  assign n24443 = n24441 & n35532 ;
  assign n24445 = n24436 | n24443 ;
  assign n24444 = n24436 & n24443 ;
  assign n35533 = ~n24444 ;
  assign n24446 = n35533 & n24445 ;
  assign n35534 = ~n20041 ;
  assign n23679 = n35534 & n23678 ;
  assign n35535 = ~n23678 ;
  assign n24447 = n20041 & n35535 ;
  assign n24448 = n23679 | n24447 ;
  assign n35536 = ~n23687 ;
  assign n24449 = n35536 & n24448 ;
  assign n35537 = ~n24448 ;
  assign n24450 = n23687 & n35537 ;
  assign n24451 = n24449 | n24450 ;
  assign n20346 = n8157 & n34399 ;
  assign n19939 = n740 & n19917 ;
  assign n19961 = n8195 & n34381 ;
  assign n24452 = n19939 | n19961 ;
  assign n24453 = n9052 & n19893 ;
  assign n24454 = n24452 | n24453 ;
  assign n24455 = n20346 | n24454 ;
  assign n24456 = x5 | n24455 ;
  assign n24457 = x5 & n24455 ;
  assign n35538 = ~n24457 ;
  assign n24458 = n24456 & n35538 ;
  assign n24460 = n24451 | n24458 ;
  assign n24459 = n24451 & n24458 ;
  assign n35539 = ~n24459 ;
  assign n24461 = n35539 & n24460 ;
  assign n20416 = n8157 & n20412 ;
  assign n19950 = n740 & n34381 ;
  assign n19988 = n8195 & n34372 ;
  assign n24462 = n19950 | n19988 ;
  assign n24463 = n9052 & n19917 ;
  assign n24464 = n24462 | n24463 ;
  assign n24465 = n20416 | n24464 ;
  assign n24466 = x5 | n24465 ;
  assign n24467 = x5 & n24465 ;
  assign n35540 = ~n24467 ;
  assign n24468 = n24466 & n35540 ;
  assign n35541 = ~n23669 ;
  assign n23676 = n35541 & n23675 ;
  assign n35542 = ~n23675 ;
  assign n24469 = n23669 & n35542 ;
  assign n24470 = n23676 | n24469 ;
  assign n24472 = n24468 | n24470 ;
  assign n24471 = n24468 & n24470 ;
  assign n35543 = ~n24471 ;
  assign n24473 = n35543 & n24472 ;
  assign n20043 = n9969 & n34367 ;
  assign n20179 = n8157 & n20170 ;
  assign n24474 = n9052 & n34350 ;
  assign n24475 = n740 & n34367 ;
  assign n24476 = n24474 | n24475 ;
  assign n24477 = n20179 | n24476 ;
  assign n24478 = n20043 | n24477 ;
  assign n24480 = x5 & n24478 ;
  assign n20003 = n9052 & n19991 ;
  assign n24481 = n740 & n34350 ;
  assign n24482 = n8195 & n34367 ;
  assign n24483 = n24481 | n24482 ;
  assign n24484 = n20003 | n24483 ;
  assign n24485 = n8157 & n20189 ;
  assign n24486 = n24484 | n24485 ;
  assign n24488 = n24480 | n24486 ;
  assign n35544 = ~n24488 ;
  assign n24489 = x5 & n35544 ;
  assign n24491 = n20039 | n24489 ;
  assign n20217 = n8157 & n20207 ;
  assign n20019 = n740 & n19991 ;
  assign n20035 = n8195 & n34350 ;
  assign n24492 = n20019 | n20035 ;
  assign n24493 = n9052 & n34372 ;
  assign n24494 = n24492 | n24493 ;
  assign n24495 = n20217 | n24494 ;
  assign n35545 = ~n24495 ;
  assign n24496 = x5 & n35545 ;
  assign n24497 = n30053 & n24495 ;
  assign n24498 = n24496 | n24497 ;
  assign n24499 = n24491 & n24498 ;
  assign n35546 = ~n23666 ;
  assign n23667 = n23662 & n35546 ;
  assign n35547 = ~n23662 ;
  assign n24500 = n35547 & n23666 ;
  assign n24501 = n23667 | n24500 ;
  assign n24502 = n24499 & n24501 ;
  assign n20281 = n8157 & n34383 ;
  assign n19970 = n740 & n34372 ;
  assign n20010 = n8195 & n19991 ;
  assign n24503 = n19970 | n20010 ;
  assign n24504 = n9052 & n34381 ;
  assign n24505 = n24503 | n24504 ;
  assign n24506 = n20281 | n24505 ;
  assign n35548 = ~n24506 ;
  assign n24507 = x5 & n35548 ;
  assign n24508 = n30053 & n24506 ;
  assign n24509 = n24507 | n24508 ;
  assign n24510 = n24499 | n24501 ;
  assign n35549 = ~n24502 ;
  assign n24511 = n35549 & n24510 ;
  assign n24513 = n24509 & n24511 ;
  assign n24514 = n24502 | n24513 ;
  assign n35550 = ~n24514 ;
  assign n24516 = n24473 & n35550 ;
  assign n35551 = ~n24516 ;
  assign n24517 = n24472 & n35551 ;
  assign n35552 = ~n24517 ;
  assign n24519 = n24461 & n35552 ;
  assign n35553 = ~n24519 ;
  assign n24520 = n24460 & n35553 ;
  assign n35554 = ~n24520 ;
  assign n24522 = n24446 & n35554 ;
  assign n35555 = ~n24522 ;
  assign n24523 = n24445 & n35555 ;
  assign n35556 = ~n24523 ;
  assign n24525 = n24434 & n35556 ;
  assign n35557 = ~n24525 ;
  assign n24526 = n24433 & n35557 ;
  assign n35558 = ~n24526 ;
  assign n24528 = n24422 & n35558 ;
  assign n35559 = ~n24528 ;
  assign n24529 = n24421 & n35559 ;
  assign n35560 = ~n24529 ;
  assign n24530 = n24410 & n35560 ;
  assign n35561 = ~n24530 ;
  assign n24531 = n24408 & n35561 ;
  assign n35562 = ~n24531 ;
  assign n24533 = n24397 & n35562 ;
  assign n35563 = ~n24533 ;
  assign n24534 = n24395 & n35563 ;
  assign n24535 = n24376 & n24383 ;
  assign n35564 = ~n24535 ;
  assign n24536 = n24384 & n35564 ;
  assign n35565 = ~n24534 ;
  assign n24537 = n35565 & n24536 ;
  assign n35566 = ~n24537 ;
  assign n24538 = n24384 & n35566 ;
  assign n24539 = n24375 & n24538 ;
  assign n24540 = n24373 | n24539 ;
  assign n24542 = n24364 & n24540 ;
  assign n24543 = n24362 | n24542 ;
  assign n24544 = n24343 & n24350 ;
  assign n24545 = n24543 | n24544 ;
  assign n24546 = n24351 & n24545 ;
  assign n35567 = ~n24546 ;
  assign n24547 = n24342 & n35567 ;
  assign n35568 = ~n24547 ;
  assign n24548 = n24340 & n35568 ;
  assign n35569 = ~n24548 ;
  assign n24550 = n24329 & n35569 ;
  assign n35570 = ~n24550 ;
  assign n24551 = n24328 & n35570 ;
  assign n24553 = n24317 & n24551 ;
  assign n23756 = n23562 | n23755 ;
  assign n24554 = n23562 & n23755 ;
  assign n35571 = ~n24554 ;
  assign n24555 = n23756 & n35571 ;
  assign n24552 = n24317 | n24551 ;
  assign n35572 = ~n24553 ;
  assign n24556 = n24552 & n35572 ;
  assign n24558 = n24555 & n24556 ;
  assign n24559 = n24553 | n24558 ;
  assign n24560 = n24310 & n24559 ;
  assign n24561 = n24309 | n24560 ;
  assign n24562 = n24299 | n24561 ;
  assign n23763 = n23539 | n23762 ;
  assign n35573 = ~n23764 ;
  assign n24563 = n23763 & n35573 ;
  assign n24564 = n24299 & n24561 ;
  assign n35574 = ~n24564 ;
  assign n24565 = n24562 & n35574 ;
  assign n35575 = ~n24563 ;
  assign n24567 = n35575 & n24565 ;
  assign n35576 = ~n24567 ;
  assign n24568 = n24562 & n35576 ;
  assign n24291 = n24283 & n24290 ;
  assign n35577 = ~n24291 ;
  assign n24569 = n35577 & n24292 ;
  assign n35578 = ~n24568 ;
  assign n24570 = n35578 & n24569 ;
  assign n35579 = ~n24570 ;
  assign n24571 = n24292 & n35579 ;
  assign n24572 = n24279 & n24571 ;
  assign n35580 = ~n23516 ;
  assign n24573 = n35580 & n23768 ;
  assign n24574 = n23769 | n24573 ;
  assign n24575 = n24279 | n24571 ;
  assign n35581 = ~n24572 ;
  assign n24576 = n35581 & n24575 ;
  assign n24577 = n24574 & n24576 ;
  assign n24578 = n24572 | n24577 ;
  assign n35582 = ~n24578 ;
  assign n24579 = n24272 & n35582 ;
  assign n35583 = ~n24579 ;
  assign n24580 = n24270 & n35583 ;
  assign n35584 = ~n24580 ;
  assign n24582 = n24260 & n35584 ;
  assign n35585 = ~n24582 ;
  assign n24583 = n24259 & n35585 ;
  assign n24247 = n24239 & n24246 ;
  assign n35586 = ~n24247 ;
  assign n24584 = n35586 & n24248 ;
  assign n35587 = ~n24583 ;
  assign n24585 = n35587 & n24584 ;
  assign n35588 = ~n24585 ;
  assign n24586 = n24248 & n35588 ;
  assign n24587 = n24229 | n24236 ;
  assign n35589 = ~n24237 ;
  assign n24588 = n35589 & n24587 ;
  assign n24589 = n24586 & n24588 ;
  assign n24590 = n24237 | n24589 ;
  assign n35590 = ~n24590 ;
  assign n24591 = n24227 & n35590 ;
  assign n35591 = ~n24591 ;
  assign n24592 = n24225 & n35591 ;
  assign n24594 = n24214 | n24592 ;
  assign n35592 = ~n24213 ;
  assign n24595 = n35592 & n24594 ;
  assign n24597 = n24186 & n24595 ;
  assign n24598 = n23425 & n23795 ;
  assign n35593 = ~n24598 ;
  assign n24599 = n23796 & n35593 ;
  assign n24596 = n24186 | n24595 ;
  assign n35594 = ~n24597 ;
  assign n24600 = n24596 & n35594 ;
  assign n35595 = ~n24599 ;
  assign n24601 = n35595 & n24600 ;
  assign n24602 = n24597 | n24601 ;
  assign n24603 = n24161 | n24602 ;
  assign n24604 = n24161 & n24602 ;
  assign n35596 = ~n24604 ;
  assign n24605 = n24603 & n35596 ;
  assign n15195 = n895 & n32875 ;
  assign n15075 = n2849 & n32856 ;
  assign n15085 = n2861 & n15081 ;
  assign n24606 = n15075 | n15085 ;
  assign n24607 = n894 & n32876 ;
  assign n24608 = n24606 | n24607 ;
  assign n24609 = n15195 | n24608 ;
  assign n24610 = x29 | n24609 ;
  assign n24611 = x29 & n24609 ;
  assign n35597 = ~n24611 ;
  assign n24612 = n24610 & n35597 ;
  assign n24613 = n35401 & n23966 ;
  assign n24614 = n23972 | n24613 ;
  assign n24615 = n190 | n489 ;
  assign n24616 = n534 | n24615 ;
  assign n24617 = n689 | n823 ;
  assign n24618 = n24616 | n24617 ;
  assign n24619 = n13351 | n24618 ;
  assign n24620 = n874 | n1147 ;
  assign n24621 = n12831 | n24620 ;
  assign n24622 = n4966 | n24621 ;
  assign n24623 = n5365 | n24622 ;
  assign n24624 = n24619 | n24623 ;
  assign n24625 = n578 | n11196 ;
  assign n24626 = n24624 | n24625 ;
  assign n24627 = n13614 | n24626 ;
  assign n24628 = n22191 | n24627 ;
  assign n35598 = ~n24628 ;
  assign n24629 = n24006 & n35598 ;
  assign n35599 = ~n24006 ;
  assign n24630 = n35599 & n24628 ;
  assign n24631 = n24629 | n24630 ;
  assign n24632 = n23966 | n24631 ;
  assign n24633 = n23966 & n24631 ;
  assign n35600 = ~n24633 ;
  assign n24634 = n24632 & n35600 ;
  assign n14577 = n889 & n14570 ;
  assign n14533 = n3329 & n32706 ;
  assign n14557 = n3311 & n14536 ;
  assign n24635 = n14533 | n14557 ;
  assign n24636 = n3343 & n32707 ;
  assign n24637 = n24635 | n24636 ;
  assign n24638 = n14577 | n24637 ;
  assign n35601 = ~n24638 ;
  assign n24639 = n24634 & n35601 ;
  assign n35602 = ~n24634 ;
  assign n24640 = n35602 & n24638 ;
  assign n24641 = n24639 | n24640 ;
  assign n35603 = ~n24641 ;
  assign n24642 = n24614 & n35603 ;
  assign n35604 = ~n24614 ;
  assign n24643 = n35604 & n24641 ;
  assign n24644 = n24642 | n24643 ;
  assign n35605 = ~n23989 ;
  assign n24645 = n23979 & n35605 ;
  assign n24646 = n24644 & n24645 ;
  assign n24647 = n24644 | n24645 ;
  assign n35606 = ~n24646 ;
  assign n24648 = n35606 & n24647 ;
  assign n24649 = n24612 & n24648 ;
  assign n24651 = n24612 | n24648 ;
  assign n35607 = ~n24649 ;
  assign n24652 = n35607 & n24651 ;
  assign n24653 = n260 & n15516 ;
  assign n15256 = n209 & n32890 ;
  assign n24654 = n3818 | n15256 ;
  assign n24655 = n3802 & n15221 ;
  assign n24656 = n24654 | n24655 ;
  assign n24657 = n24653 | n24656 ;
  assign n24658 = x26 | n24657 ;
  assign n24659 = x26 & n24657 ;
  assign n35608 = ~n24659 ;
  assign n24660 = n24658 & n35608 ;
  assign n24661 = n24000 | n24003 ;
  assign n35609 = ~n24661 ;
  assign n24662 = n24660 & n35609 ;
  assign n35610 = ~n24660 ;
  assign n24663 = n35610 & n24661 ;
  assign n24664 = n24662 | n24663 ;
  assign n35611 = ~n24652 ;
  assign n24665 = n35611 & n24664 ;
  assign n35612 = ~n24664 ;
  assign n24667 = n24652 & n35612 ;
  assign n24668 = n24665 | n24667 ;
  assign n35613 = ~n24012 ;
  assign n24669 = n24010 & n35613 ;
  assign n24670 = n24668 & n24669 ;
  assign n24671 = n24668 | n24669 ;
  assign n35614 = ~n24670 ;
  assign n24672 = n35614 & n24671 ;
  assign n35615 = ~n24150 ;
  assign n24673 = n24015 & n35615 ;
  assign n35616 = ~n24673 ;
  assign n24674 = n24672 & n35616 ;
  assign n35617 = ~n24672 ;
  assign n24675 = n35617 & n24673 ;
  assign n24676 = n24674 | n24675 ;
  assign n24690 = n9552 & n24676 ;
  assign n24699 = n461 | n495 ;
  assign n24700 = n897 | n24699 ;
  assign n24701 = n5861 | n24700 ;
  assign n24702 = n4854 | n5591 ;
  assign n24703 = n24701 | n24702 ;
  assign n24704 = n1135 | n1311 ;
  assign n24705 = n1468 | n24704 ;
  assign n24706 = n905 | n972 ;
  assign n24707 = n2208 | n24706 ;
  assign n24708 = n24705 | n24707 ;
  assign n24709 = n5014 | n24708 ;
  assign n24710 = n24703 | n24709 ;
  assign n35618 = ~n24710 ;
  assign n24711 = n5080 & n35618 ;
  assign n24712 = n32836 & n24711 ;
  assign n35619 = ~n24631 ;
  assign n24713 = n23966 & n35619 ;
  assign n24714 = n24630 | n24713 ;
  assign n35620 = ~n24714 ;
  assign n24715 = n24712 & n35620 ;
  assign n35621 = ~n24712 ;
  assign n24716 = n35621 & n24714 ;
  assign n24717 = n24715 | n24716 ;
  assign n15299 = n889 & n15288 ;
  assign n14511 = n3329 & n32707 ;
  assign n14534 = n3311 & n32706 ;
  assign n24718 = n14511 | n14534 ;
  assign n24719 = n3343 & n15081 ;
  assign n24720 = n24718 | n24719 ;
  assign n24721 = n15299 | n24720 ;
  assign n35622 = ~n24721 ;
  assign n24722 = n24717 & n35622 ;
  assign n35623 = ~n24717 ;
  assign n24723 = n35623 & n24721 ;
  assign n24724 = n24722 | n24723 ;
  assign n24725 = n24639 | n24642 ;
  assign n35624 = ~n24725 ;
  assign n24726 = n24724 & n35624 ;
  assign n35625 = ~n24724 ;
  assign n24727 = n35625 & n24725 ;
  assign n24728 = n24726 | n24727 ;
  assign n15268 = n895 & n32889 ;
  assign n15077 = n2861 & n32856 ;
  assign n15179 = n2849 & n32876 ;
  assign n24729 = n15077 | n15179 ;
  assign n24730 = n894 & n32890 ;
  assign n24731 = n24729 | n24730 ;
  assign n24732 = n15268 | n24731 ;
  assign n35626 = ~n24732 ;
  assign n24733 = x29 & n35626 ;
  assign n24734 = n30024 & n24732 ;
  assign n24735 = n24733 | n24734 ;
  assign n24736 = n24728 | n24735 ;
  assign n24737 = n24728 & n24735 ;
  assign n35627 = ~n24737 ;
  assign n24738 = n24736 & n35627 ;
  assign n24739 = n191 & n23876 ;
  assign n24740 = n30019 & n114 ;
  assign n24741 = n122 | n24740 ;
  assign n24742 = n115 | n24741 ;
  assign n24744 = n128 & n15221 ;
  assign n35628 = ~n24744 ;
  assign n24745 = n24742 & n35628 ;
  assign n35629 = ~n24739 ;
  assign n24746 = n35629 & n24745 ;
  assign n24747 = n24738 & n24746 ;
  assign n24748 = n24738 | n24746 ;
  assign n35630 = ~n24747 ;
  assign n24749 = n35630 & n24748 ;
  assign n35631 = ~n24612 ;
  assign n24650 = n35631 & n24648 ;
  assign n35632 = ~n24650 ;
  assign n24750 = n24647 & n35632 ;
  assign n35633 = ~n24749 ;
  assign n24751 = n35633 & n24750 ;
  assign n35634 = ~n24750 ;
  assign n24752 = n24749 & n35634 ;
  assign n24753 = n24751 | n24752 ;
  assign n24666 = n24652 & n24664 ;
  assign n24754 = n24660 & n24661 ;
  assign n24755 = n24666 | n24754 ;
  assign n35635 = ~n24755 ;
  assign n24756 = n24753 & n35635 ;
  assign n35636 = ~n24753 ;
  assign n24757 = n35636 & n24755 ;
  assign n24758 = n24756 | n24757 ;
  assign n35637 = ~n24674 ;
  assign n24759 = n24671 & n35637 ;
  assign n24761 = n24758 | n24759 ;
  assign n35638 = ~n24756 ;
  assign n24762 = n35638 & n24761 ;
  assign n24763 = n487 | n845 ;
  assign n24764 = n1596 | n24763 ;
  assign n24765 = n4630 | n13571 ;
  assign n24766 = n24764 | n24765 ;
  assign n24767 = n3737 | n3963 ;
  assign n24768 = n24766 | n24767 ;
  assign n24769 = n1633 | n24768 ;
  assign n24770 = n5865 | n24769 ;
  assign n24771 = n4993 | n24770 ;
  assign n24772 = n24711 | n24771 ;
  assign n24773 = n24712 & n24771 ;
  assign n35639 = ~n24773 ;
  assign n24774 = n24772 & n35639 ;
  assign n15117 = n889 & n15111 ;
  assign n14493 = n3311 & n32707 ;
  assign n15095 = n3329 & n15081 ;
  assign n24775 = n14493 | n15095 ;
  assign n24776 = n3343 & n32856 ;
  assign n24777 = n24775 | n24776 ;
  assign n24778 = n15117 | n24777 ;
  assign n35640 = ~n24778 ;
  assign n24779 = n24774 & n35640 ;
  assign n35641 = ~n24774 ;
  assign n24781 = n35641 & n24778 ;
  assign n24782 = n24779 | n24781 ;
  assign n24783 = n24712 & n24714 ;
  assign n24784 = n24717 & n24721 ;
  assign n24785 = n24783 | n24784 ;
  assign n35642 = ~n24785 ;
  assign n24786 = n24782 & n35642 ;
  assign n35643 = ~n24782 ;
  assign n24787 = n35643 & n24785 ;
  assign n24788 = n24786 | n24787 ;
  assign n35644 = ~n24727 ;
  assign n24789 = n35644 & n24736 ;
  assign n24790 = n24788 & n24789 ;
  assign n24791 = n24788 | n24789 ;
  assign n35645 = ~n24790 ;
  assign n24792 = n35645 & n24791 ;
  assign n15532 = n895 & n15526 ;
  assign n15166 = n2861 & n32876 ;
  assign n15246 = n894 & n15221 ;
  assign n24793 = n15166 | n15246 ;
  assign n24794 = n2849 & n32890 ;
  assign n24795 = n24793 | n24794 ;
  assign n24796 = n15532 | n24795 ;
  assign n35646 = ~n24796 ;
  assign n24797 = x29 & n35646 ;
  assign n24798 = n30024 & n24796 ;
  assign n24799 = n24797 | n24798 ;
  assign n24800 = n24741 | n24799 ;
  assign n24801 = n24741 & n24799 ;
  assign n35647 = ~n24801 ;
  assign n24802 = n24800 & n35647 ;
  assign n35648 = ~n24792 ;
  assign n24803 = n35648 & n24802 ;
  assign n35649 = ~n24802 ;
  assign n24805 = n24792 & n35649 ;
  assign n24806 = n24803 | n24805 ;
  assign n35650 = ~n24746 ;
  assign n24807 = n24738 & n35650 ;
  assign n24808 = n24749 | n24750 ;
  assign n35651 = ~n24807 ;
  assign n24809 = n35651 & n24808 ;
  assign n24810 = n24806 & n24809 ;
  assign n24811 = n24806 | n24809 ;
  assign n35652 = ~n24810 ;
  assign n24812 = n35652 & n24811 ;
  assign n24813 = n24762 & n24812 ;
  assign n24814 = n24762 | n24812 ;
  assign n35653 = ~n24813 ;
  assign n24815 = n35653 & n24814 ;
  assign n35654 = ~n24758 ;
  assign n24760 = n35654 & n24759 ;
  assign n35655 = ~n24759 ;
  assign n24837 = n24758 & n35655 ;
  assign n24838 = n24760 | n24837 ;
  assign n35656 = ~n24080 ;
  assign n24865 = n35656 & n24133 ;
  assign n35657 = ~n24865 ;
  assign n24866 = n24057 & n35657 ;
  assign n24867 = n24676 | n24866 ;
  assign n24868 = n24838 | n24867 ;
  assign n35658 = ~n24129 ;
  assign n24860 = n24080 & n35658 ;
  assign n24862 = n24057 | n24860 ;
  assign n24864 = n24676 & n24862 ;
  assign n24869 = n24838 & n24864 ;
  assign n35659 = ~n24869 ;
  assign n24870 = n24868 & n35659 ;
  assign n35660 = ~n24870 ;
  assign n24871 = n24815 & n35660 ;
  assign n35661 = ~n24815 ;
  assign n24872 = n35661 & n24870 ;
  assign n24873 = n24871 | n24872 ;
  assign n35662 = ~n24873 ;
  assign n24874 = n9562 & n35662 ;
  assign n24885 = n10105 & n24815 ;
  assign n35663 = ~n24838 ;
  assign n24886 = n10126 & n35663 ;
  assign n24887 = n24885 | n24886 ;
  assign n24888 = n24874 | n24887 ;
  assign n35664 = ~n24888 ;
  assign n24889 = x2 & n35664 ;
  assign n24890 = n30049 & n24888 ;
  assign n24891 = n24889 | n24890 ;
  assign n35665 = ~n24690 ;
  assign n24892 = n35665 & n24891 ;
  assign n24894 = n24605 | n24892 ;
  assign n24893 = n24605 & n24892 ;
  assign n35666 = ~n24600 ;
  assign n25312 = n24599 & n35666 ;
  assign n25313 = n24601 | n25312 ;
  assign n35667 = ~n24862 ;
  assign n24863 = n24676 & n35667 ;
  assign n35668 = ~n24676 ;
  assign n25314 = n35668 & n24866 ;
  assign n25315 = n24863 | n25314 ;
  assign n25316 = n35663 & n25315 ;
  assign n35669 = ~n25315 ;
  assign n25317 = n24838 & n35669 ;
  assign n25318 = n25316 | n25317 ;
  assign n35670 = ~n25318 ;
  assign n25319 = n9562 & n35670 ;
  assign n24072 = n9552 & n24057 ;
  assign n24685 = n10126 & n24676 ;
  assign n25330 = n24072 | n24685 ;
  assign n25331 = n10105 & n35663 ;
  assign n25332 = n25330 | n25331 ;
  assign n25333 = n25319 | n25332 ;
  assign n35671 = ~n25333 ;
  assign n25334 = x2 & n35671 ;
  assign n25335 = n30049 & n25333 ;
  assign n25336 = n25334 | n25335 ;
  assign n35672 = ~n25336 ;
  assign n25337 = n25313 & n35672 ;
  assign n35673 = ~n24227 ;
  assign n24895 = n35673 & n24590 ;
  assign n24896 = n24591 | n24895 ;
  assign n24118 = n9552 & n35458 ;
  assign n24140 = n9562 & n35457 ;
  assign n24897 = n10105 & n24151 ;
  assign n24898 = n10126 & n24080 ;
  assign n24899 = n24897 | n24898 ;
  assign n24900 = n24140 | n24899 ;
  assign n35674 = ~n24900 ;
  assign n24901 = x2 & n35674 ;
  assign n24902 = n30049 & n24900 ;
  assign n24903 = n24901 | n24902 ;
  assign n35675 = ~n24118 ;
  assign n24904 = n35675 & n24903 ;
  assign n24906 = n24896 | n24904 ;
  assign n24905 = n24896 & n24904 ;
  assign n24907 = n24586 | n24588 ;
  assign n35676 = ~n24589 ;
  assign n24908 = n35676 & n24907 ;
  assign n24170 = n9562 & n24168 ;
  assign n23295 = n9552 & n35467 ;
  assign n24121 = n10126 & n35458 ;
  assign n24909 = n23295 | n24121 ;
  assign n24910 = n10105 & n24080 ;
  assign n24911 = n24909 | n24910 ;
  assign n24912 = n24170 | n24911 ;
  assign n35677 = ~n24912 ;
  assign n24913 = x2 & n35677 ;
  assign n24914 = n30049 & n24912 ;
  assign n24915 = n24913 | n24914 ;
  assign n24916 = n24908 | n24915 ;
  assign n24917 = n24908 & n24915 ;
  assign n35678 = ~n24584 ;
  assign n24918 = n24583 & n35678 ;
  assign n24919 = n24585 | n24918 ;
  assign n24195 = n9562 & n35472 ;
  assign n23301 = n10126 & n35467 ;
  assign n23328 = n9552 & n35244 ;
  assign n24920 = n23301 | n23328 ;
  assign n24921 = n10105 & n35465 ;
  assign n24922 = n24920 | n24921 ;
  assign n24923 = n24195 | n24922 ;
  assign n35679 = ~n24923 ;
  assign n24924 = x2 & n35679 ;
  assign n24925 = n30049 & n24923 ;
  assign n24926 = n24924 | n24925 ;
  assign n24927 = n24919 | n24926 ;
  assign n24928 = n24919 & n24926 ;
  assign n35680 = ~n24260 ;
  assign n24581 = n35680 & n24580 ;
  assign n24929 = n24581 | n24582 ;
  assign n23354 = n9552 & n23339 ;
  assign n23375 = n9562 & n23372 ;
  assign n24930 = n10105 & n35246 ;
  assign n24931 = n10126 & n35254 ;
  assign n24932 = n24930 | n24931 ;
  assign n24933 = n23375 | n24932 ;
  assign n35681 = ~n24933 ;
  assign n24934 = x2 & n35681 ;
  assign n24935 = n30049 & n24933 ;
  assign n24936 = n24934 | n24935 ;
  assign n35682 = ~n23354 ;
  assign n24937 = n35682 & n24936 ;
  assign n25275 = n24929 | n24937 ;
  assign n24938 = n24574 | n24576 ;
  assign n35683 = ~n24577 ;
  assign n24939 = n35683 & n24938 ;
  assign n35684 = ~n24569 ;
  assign n24940 = n24568 & n35684 ;
  assign n24941 = n24570 | n24940 ;
  assign n24566 = n24563 & n24565 ;
  assign n24942 = n24563 | n24565 ;
  assign n35685 = ~n24566 ;
  assign n24943 = n35685 & n24942 ;
  assign n22548 = n10126 & n35018 ;
  assign n22584 = n10105 & n22533 ;
  assign n24944 = n22548 | n22584 ;
  assign n24945 = n9562 & n35030 ;
  assign n24946 = n24944 | n24945 ;
  assign n24947 = n30049 & n24946 ;
  assign n21737 = n31643 & n21729 ;
  assign n35686 = ~n21737 ;
  assign n24948 = x2 & n35686 ;
  assign n35687 = ~n24946 ;
  assign n24949 = n35687 & n24948 ;
  assign n24950 = n24947 | n24949 ;
  assign n24951 = n24943 & n24950 ;
  assign n24952 = n24943 | n24950 ;
  assign n35688 = ~n24309 ;
  assign n24953 = n35688 & n24310 ;
  assign n35689 = ~n24953 ;
  assign n24954 = n24559 & n35689 ;
  assign n35690 = ~n24559 ;
  assign n24955 = n35690 & n24953 ;
  assign n24956 = n24954 | n24955 ;
  assign n22648 = n9562 & n35035 ;
  assign n21732 = n10126 & n21729 ;
  assign n21816 = n9552 & n21753 ;
  assign n24957 = n21732 | n21816 ;
  assign n24958 = n10105 & n35018 ;
  assign n24959 = n24957 | n24958 ;
  assign n24960 = n22648 | n24959 ;
  assign n35691 = ~n24960 ;
  assign n24961 = x2 & n35691 ;
  assign n24963 = n30049 & n24960 ;
  assign n24964 = n24961 | n24963 ;
  assign n24965 = n24956 & n24964 ;
  assign n24962 = x2 | n24960 ;
  assign n24966 = x2 & n24960 ;
  assign n35692 = ~n24966 ;
  assign n24967 = n24962 & n35692 ;
  assign n24968 = n24956 | n24967 ;
  assign n24557 = n24555 | n24556 ;
  assign n35693 = ~n24558 ;
  assign n24969 = n24557 & n35693 ;
  assign n35694 = ~n24329 ;
  assign n24549 = n35694 & n24548 ;
  assign n24970 = n24549 | n24550 ;
  assign n35695 = ~n24342 ;
  assign n24971 = n35695 & n24546 ;
  assign n24972 = n24547 | n24971 ;
  assign n21873 = n9562 & n34817 ;
  assign n19668 = n10126 & n34360 ;
  assign n19683 = n9552 & n34349 ;
  assign n24973 = n19668 | n19683 ;
  assign n24974 = n10105 & n34803 ;
  assign n24975 = n24973 | n24974 ;
  assign n24976 = n21873 | n24975 ;
  assign n24977 = x2 | n24976 ;
  assign n24979 = x2 & n24976 ;
  assign n35696 = ~n24979 ;
  assign n24980 = n24977 & n35696 ;
  assign n24981 = n24972 | n24980 ;
  assign n35697 = ~n24976 ;
  assign n24978 = x2 & n35697 ;
  assign n24982 = n30049 & n24976 ;
  assign n24983 = n24978 | n24982 ;
  assign n24984 = n24972 & n24983 ;
  assign n35698 = ~n24544 ;
  assign n24985 = n24351 & n35698 ;
  assign n24986 = n24543 & n24985 ;
  assign n24987 = n24543 | n24985 ;
  assign n35699 = ~n24986 ;
  assign n24988 = n35699 & n24987 ;
  assign n20148 = n9562 & n34362 ;
  assign n24989 = n10105 & n34365 ;
  assign n24990 = n10126 & n34349 ;
  assign n24991 = n24989 | n24990 ;
  assign n24992 = n20148 | n24991 ;
  assign n24993 = n30049 & n24992 ;
  assign n19706 = n733 | n19705 ;
  assign n24994 = x2 & n19706 ;
  assign n35700 = ~n24992 ;
  assign n24995 = n35700 & n24994 ;
  assign n24996 = n24993 | n24995 ;
  assign n24997 = n24988 | n24996 ;
  assign n24998 = n24988 & n24996 ;
  assign n21077 = n9562 & n34598 ;
  assign n19719 = n10126 & n34363 ;
  assign n19742 = n9552 & n34520 ;
  assign n24999 = n19719 | n19742 ;
  assign n25000 = n10105 & n34349 ;
  assign n25001 = n24999 | n25000 ;
  assign n25002 = n21077 | n25001 ;
  assign n25003 = x2 | n25002 ;
  assign n25004 = x2 & n25002 ;
  assign n35701 = ~n25004 ;
  assign n25005 = n25003 & n35701 ;
  assign n24541 = n24364 | n24540 ;
  assign n35702 = ~n24542 ;
  assign n25006 = n24541 & n35702 ;
  assign n25007 = n25005 | n25006 ;
  assign n25008 = n25005 & n25006 ;
  assign n25009 = n24375 | n24538 ;
  assign n35703 = ~n24539 ;
  assign n25010 = n35703 & n25009 ;
  assign n19761 = n9552 & n19752 ;
  assign n21101 = n9562 & n34603 ;
  assign n25011 = n10105 & n34596 ;
  assign n25012 = n10126 & n34520 ;
  assign n25013 = n25011 | n25012 ;
  assign n25014 = n21101 | n25013 ;
  assign n35704 = ~n25014 ;
  assign n25015 = x2 & n35704 ;
  assign n25016 = n30049 & n25014 ;
  assign n25017 = n25015 | n25016 ;
  assign n35705 = ~n19761 ;
  assign n25018 = n35705 & n25017 ;
  assign n25019 = n25010 | n25018 ;
  assign n25020 = n25010 & n25018 ;
  assign n35706 = ~n24536 ;
  assign n25021 = n24534 & n35706 ;
  assign n25022 = n24537 | n25021 ;
  assign n19785 = n9552 & n34519 ;
  assign n20813 = n9562 & n20805 ;
  assign n25023 = n10105 & n34520 ;
  assign n25024 = n10126 & n20845 ;
  assign n25025 = n25023 | n25024 ;
  assign n25026 = n20813 | n25025 ;
  assign n35707 = ~n25026 ;
  assign n25027 = x2 & n35707 ;
  assign n25028 = n30049 & n25026 ;
  assign n25029 = n25027 | n25028 ;
  assign n35708 = ~n19785 ;
  assign n25030 = n35708 & n25029 ;
  assign n25031 = n25022 | n25030 ;
  assign n35709 = ~n24397 ;
  assign n24532 = n35709 & n24531 ;
  assign n25032 = n24532 | n24533 ;
  assign n20841 = n9562 & n20833 ;
  assign n19792 = n10126 & n34519 ;
  assign n19815 = n9552 & n34355 ;
  assign n25033 = n19792 | n19815 ;
  assign n25034 = n10105 & n20845 ;
  assign n25035 = n25033 | n25034 ;
  assign n25036 = n20841 | n25035 ;
  assign n25037 = x2 | n25036 ;
  assign n25038 = x2 & n25036 ;
  assign n35710 = ~n25038 ;
  assign n25039 = n25037 & n35710 ;
  assign n25040 = n25032 & n25039 ;
  assign n25192 = n25032 | n25039 ;
  assign n35711 = ~n24410 ;
  assign n25041 = n35711 & n24529 ;
  assign n25042 = n24530 | n25041 ;
  assign n20866 = n9562 & n20863 ;
  assign n19817 = n10126 & n34355 ;
  assign n19831 = n9552 & n19824 ;
  assign n25043 = n19817 | n19831 ;
  assign n25044 = n10105 & n34536 ;
  assign n25045 = n25043 | n25044 ;
  assign n25046 = n20866 | n25045 ;
  assign n35712 = ~n25046 ;
  assign n25047 = x2 & n35712 ;
  assign n25048 = n30049 & n25046 ;
  assign n25049 = n25047 | n25048 ;
  assign n25051 = n25042 & n25049 ;
  assign n25050 = n25042 | n25049 ;
  assign n24527 = n24422 & n24526 ;
  assign n25052 = n24422 | n24526 ;
  assign n35713 = ~n24527 ;
  assign n25053 = n35713 & n25052 ;
  assign n20107 = n9552 & n34354 ;
  assign n20783 = n9562 & n34511 ;
  assign n25054 = n10105 & n34513 ;
  assign n25055 = n10126 & n20527 ;
  assign n25056 = n25054 | n25055 ;
  assign n25057 = n20783 | n25056 ;
  assign n35714 = ~n25057 ;
  assign n25058 = x2 & n35714 ;
  assign n25059 = n30049 & n25057 ;
  assign n25060 = n25058 | n25059 ;
  assign n35715 = ~n20107 ;
  assign n25061 = n35715 & n25060 ;
  assign n25062 = n25053 & n25061 ;
  assign n25187 = n25053 | n25061 ;
  assign n24524 = n24434 & n24523 ;
  assign n25063 = n24434 | n24523 ;
  assign n35716 = ~n24524 ;
  assign n25064 = n35716 & n25063 ;
  assign n20523 = n9562 & n34442 ;
  assign n20086 = n9552 & n20067 ;
  assign n20106 = n10126 & n34354 ;
  assign n25065 = n20086 | n20106 ;
  assign n25066 = n10105 & n20527 ;
  assign n25067 = n25065 | n25066 ;
  assign n25068 = n20523 | n25067 ;
  assign n35717 = ~n25068 ;
  assign n25069 = x2 & n35717 ;
  assign n25070 = n30049 & n25068 ;
  assign n25071 = n25069 | n25070 ;
  assign n25073 = n25064 & n25071 ;
  assign n25072 = n25064 | n25071 ;
  assign n24521 = n24446 & n24520 ;
  assign n25074 = n24446 | n24520 ;
  assign n35718 = ~n24521 ;
  assign n25075 = n35718 & n25074 ;
  assign n20553 = n9562 & n34450 ;
  assign n19864 = n9552 & n19846 ;
  assign n20087 = n10126 & n20067 ;
  assign n25076 = n19864 | n20087 ;
  assign n25077 = n10105 & n34452 ;
  assign n25078 = n25076 | n25077 ;
  assign n25079 = n20553 | n25078 ;
  assign n35719 = ~n25079 ;
  assign n25080 = x2 & n35719 ;
  assign n25081 = n30049 & n25079 ;
  assign n25082 = n25080 | n25081 ;
  assign n25084 = n25075 & n25082 ;
  assign n25083 = n25075 | n25082 ;
  assign n24518 = n24461 & n24517 ;
  assign n25085 = n24461 | n24517 ;
  assign n35720 = ~n24518 ;
  assign n25086 = n35720 & n25085 ;
  assign n20589 = n9562 & n20579 ;
  assign n19860 = n10126 & n19846 ;
  assign n19885 = n9552 & n19870 ;
  assign n25087 = n19860 | n19885 ;
  assign n25088 = n10105 & n20067 ;
  assign n25089 = n25087 | n25088 ;
  assign n25090 = n20589 | n25089 ;
  assign n35721 = ~n25090 ;
  assign n25091 = x2 & n35721 ;
  assign n25092 = n30049 & n25090 ;
  assign n25093 = n25091 | n25092 ;
  assign n25095 = n25086 & n25093 ;
  assign n25094 = n25086 | n25093 ;
  assign n19913 = n9552 & n19893 ;
  assign n20496 = n9562 & n20486 ;
  assign n25096 = n10105 & n19846 ;
  assign n25097 = n10126 & n19870 ;
  assign n25098 = n25096 | n25097 ;
  assign n25099 = n20496 | n25098 ;
  assign n35722 = ~n25099 ;
  assign n25100 = x2 & n35722 ;
  assign n25101 = n30049 & n25099 ;
  assign n25102 = n25100 | n25101 ;
  assign n35723 = ~n19913 ;
  assign n25103 = n35723 & n25102 ;
  assign n35724 = ~n24509 ;
  assign n24512 = n35724 & n24511 ;
  assign n35725 = ~n24511 ;
  assign n25104 = n24509 & n35725 ;
  assign n25105 = n24512 | n25104 ;
  assign n19930 = n9552 & n19917 ;
  assign n20314 = n9562 & n20311 ;
  assign n25106 = n10105 & n19870 ;
  assign n25107 = n10126 & n19893 ;
  assign n25108 = n25106 | n25107 ;
  assign n25109 = n20314 | n25108 ;
  assign n35726 = ~n25109 ;
  assign n25110 = x2 & n35726 ;
  assign n25111 = n30049 & n25109 ;
  assign n25112 = n25110 | n25111 ;
  assign n35727 = ~n19930 ;
  assign n25113 = n35727 & n25112 ;
  assign n25115 = n25105 & n25113 ;
  assign n25114 = n25105 | n25113 ;
  assign n35728 = ~n20039 ;
  assign n24490 = n35728 & n24489 ;
  assign n35729 = ~n24489 ;
  assign n25116 = n20039 & n35729 ;
  assign n25117 = n24490 | n25116 ;
  assign n35730 = ~n24498 ;
  assign n25118 = n35730 & n25117 ;
  assign n35731 = ~n25117 ;
  assign n25119 = n24498 & n35731 ;
  assign n25120 = n25118 | n25119 ;
  assign n24487 = n24480 & n24486 ;
  assign n35732 = ~n24487 ;
  assign n25121 = n35732 & n24488 ;
  assign n19940 = n10105 & n19917 ;
  assign n19962 = n10126 & n34381 ;
  assign n25122 = n19940 | n19962 ;
  assign n25123 = n9562 & n20412 ;
  assign n25124 = n25122 | n25123 ;
  assign n25125 = x2 & n25124 ;
  assign n19989 = n733 | n19968 ;
  assign n25126 = x2 & n19989 ;
  assign n25127 = n25124 | n25126 ;
  assign n35733 = ~n25125 ;
  assign n25128 = n35733 & n25127 ;
  assign n25130 = n25121 & n25128 ;
  assign n25129 = n25121 | n25128 ;
  assign n35734 = ~n24477 ;
  assign n24479 = n20043 & n35734 ;
  assign n35735 = ~n20043 ;
  assign n25131 = n35735 & n24477 ;
  assign n25132 = n24479 | n25131 ;
  assign n19981 = n10105 & n34372 ;
  assign n20020 = n10126 & n19991 ;
  assign n25133 = n19981 | n20020 ;
  assign n25134 = n9562 & n20207 ;
  assign n25135 = n25133 | n25134 ;
  assign n25136 = x2 & n25135 ;
  assign n20036 = n733 | n20022 ;
  assign n25137 = x2 & n20036 ;
  assign n25143 = n25135 | n25137 ;
  assign n25138 = n738 & n34367 ;
  assign n20017 = x0 & n19991 ;
  assign n25139 = x2 & n20038 ;
  assign n25140 = n19346 & n34350 ;
  assign n35736 = ~n25140 ;
  assign n25141 = n25139 & n35736 ;
  assign n35737 = ~n20017 ;
  assign n25142 = n35737 & n25141 ;
  assign n25144 = n25138 | n25142 ;
  assign n25145 = n25143 & n25144 ;
  assign n35738 = ~n25136 ;
  assign n25146 = n35738 & n25145 ;
  assign n25147 = n25132 & n25146 ;
  assign n20280 = n9562 & n34383 ;
  assign n25148 = n10105 & n34381 ;
  assign n25149 = n10126 & n34372 ;
  assign n25150 = n25148 | n25149 ;
  assign n25151 = n20280 | n25150 ;
  assign n25153 = x2 | n25151 ;
  assign n25152 = x2 & n25151 ;
  assign n25154 = n9552 & n19991 ;
  assign n25155 = n25132 | n25146 ;
  assign n35739 = ~n25154 ;
  assign n25156 = n35739 & n25155 ;
  assign n35740 = ~n25152 ;
  assign n25157 = n35740 & n25156 ;
  assign n25158 = n25153 & n25157 ;
  assign n25159 = n25147 | n25158 ;
  assign n25160 = n25129 & n25159 ;
  assign n25161 = n25130 | n25160 ;
  assign n25163 = n25120 & n25161 ;
  assign n25162 = n25120 | n25161 ;
  assign n19914 = n10105 & n19893 ;
  assign n19937 = n10126 & n19917 ;
  assign n25164 = n19914 | n19937 ;
  assign n25165 = n9562 & n34399 ;
  assign n25166 = n25164 | n25165 ;
  assign n25167 = x2 & n25166 ;
  assign n25168 = n9552 & n34381 ;
  assign n25169 = x2 | n25166 ;
  assign n35741 = ~n25168 ;
  assign n25170 = n35741 & n25169 ;
  assign n35742 = ~n25167 ;
  assign n25171 = n35742 & n25170 ;
  assign n25172 = n25162 & n25171 ;
  assign n25173 = n25163 | n25172 ;
  assign n25174 = n25114 & n25173 ;
  assign n25175 = n25115 | n25174 ;
  assign n25176 = n25103 & n25175 ;
  assign n24515 = n24473 | n24514 ;
  assign n25177 = n24473 & n24514 ;
  assign n35743 = ~n25177 ;
  assign n25178 = n24515 & n35743 ;
  assign n25179 = n25176 | n25178 ;
  assign n25180 = n25103 | n25175 ;
  assign n25181 = n25179 & n25180 ;
  assign n25182 = n25094 & n25181 ;
  assign n25183 = n25095 | n25182 ;
  assign n25184 = n25083 & n25183 ;
  assign n25185 = n25084 | n25184 ;
  assign n25186 = n25072 & n25185 ;
  assign n25188 = n25073 | n25186 ;
  assign n25189 = n25187 & n25188 ;
  assign n25190 = n25062 | n25189 ;
  assign n25191 = n25050 & n25190 ;
  assign n25193 = n25051 | n25191 ;
  assign n25194 = n25192 & n25193 ;
  assign n25195 = n25040 | n25194 ;
  assign n25196 = n25031 & n25195 ;
  assign n25197 = n25022 & n25030 ;
  assign n25198 = n25196 | n25197 ;
  assign n25199 = n25020 | n25198 ;
  assign n25200 = n25019 & n25199 ;
  assign n25201 = n25008 | n25200 ;
  assign n25202 = n25007 & n25201 ;
  assign n25203 = n24998 | n25202 ;
  assign n25204 = n24997 & n25203 ;
  assign n25205 = n24984 | n25204 ;
  assign n25206 = n24981 & n25205 ;
  assign n25208 = n24970 & n25206 ;
  assign n25207 = n24970 | n25206 ;
  assign n21762 = n10126 & n34803 ;
  assign n21807 = n10105 & n21753 ;
  assign n25209 = n21762 | n21807 ;
  assign n25210 = n9562 & n21848 ;
  assign n25211 = n25209 | n25210 ;
  assign n25212 = x2 & n25211 ;
  assign n25213 = n9552 & n34365 ;
  assign n25214 = x2 | n25211 ;
  assign n35744 = ~n25213 ;
  assign n25215 = n35744 & n25214 ;
  assign n35745 = ~n25212 ;
  assign n25216 = n35745 & n25215 ;
  assign n25217 = n25207 & n25216 ;
  assign n25218 = n25208 | n25217 ;
  assign n25219 = n24969 | n25218 ;
  assign n21796 = n9562 & n34802 ;
  assign n25220 = n10105 & n21804 ;
  assign n25221 = n10126 & n21753 ;
  assign n25222 = n25220 | n25221 ;
  assign n25223 = n21796 | n25222 ;
  assign n25224 = x2 | n25223 ;
  assign n25225 = x2 & n25223 ;
  assign n35746 = ~n25225 ;
  assign n25226 = n25224 & n35746 ;
  assign n25227 = n9552 & n34803 ;
  assign n35747 = ~n25227 ;
  assign n25228 = n25226 & n35747 ;
  assign n25229 = n25219 & n25228 ;
  assign n25230 = n24969 & n25218 ;
  assign n25231 = n25229 | n25230 ;
  assign n25232 = n24968 & n25231 ;
  assign n25233 = n24965 | n25232 ;
  assign n25234 = n24952 & n25233 ;
  assign n25235 = n24951 | n25234 ;
  assign n25237 = n24941 & n25235 ;
  assign n25236 = n24941 | n25235 ;
  assign n22517 = n10105 & n35020 ;
  assign n22589 = n10126 & n22533 ;
  assign n25238 = n22517 | n22589 ;
  assign n25239 = n9562 & n35022 ;
  assign n25240 = n25238 | n25239 ;
  assign n25241 = x2 & n25240 ;
  assign n25242 = n9552 & n35018 ;
  assign n25243 = x2 | n25240 ;
  assign n35748 = ~n25242 ;
  assign n25244 = n35748 & n25243 ;
  assign n35749 = ~n25241 ;
  assign n25245 = n35749 & n25244 ;
  assign n25246 = n25236 & n25245 ;
  assign n25247 = n25237 | n25246 ;
  assign n25248 = n24939 | n25247 ;
  assign n23438 = n9562 & n35262 ;
  assign n25249 = n10126 & n35020 ;
  assign n25250 = n10105 & n23444 ;
  assign n25251 = n25249 | n25250 ;
  assign n25252 = n23438 | n25251 ;
  assign n25253 = x2 | n25252 ;
  assign n25254 = x2 & n25252 ;
  assign n35750 = ~n25254 ;
  assign n25255 = n25253 & n35750 ;
  assign n25256 = n9552 & n22533 ;
  assign n35751 = ~n25256 ;
  assign n25257 = n25255 & n35751 ;
  assign n25258 = n25248 & n25257 ;
  assign n25259 = n24939 & n25247 ;
  assign n25260 = n25258 | n25259 ;
  assign n35752 = ~n24272 ;
  assign n25261 = n35752 & n24578 ;
  assign n25262 = n24579 | n25261 ;
  assign n25263 = n25260 | n25262 ;
  assign n23407 = n9562 & n35252 ;
  assign n22516 = n9552 & n35020 ;
  assign n23348 = n10126 & n23339 ;
  assign n25264 = n22516 | n23348 ;
  assign n25265 = n10105 & n35254 ;
  assign n25266 = n25264 | n25265 ;
  assign n25267 = n23407 | n25266 ;
  assign n35753 = ~n25267 ;
  assign n25268 = x2 & n35753 ;
  assign n25269 = n30049 & n25267 ;
  assign n25270 = n25268 | n25269 ;
  assign n25271 = n25263 & n25270 ;
  assign n25272 = n24929 & n24937 ;
  assign n25273 = n25260 & n25262 ;
  assign n25274 = n25272 | n25273 ;
  assign n25276 = n25271 | n25274 ;
  assign n25277 = n25275 & n25276 ;
  assign n25278 = n24928 | n25277 ;
  assign n25279 = n24927 & n25278 ;
  assign n25280 = n24917 | n25279 ;
  assign n25281 = n24916 & n25280 ;
  assign n25282 = n24905 | n25281 ;
  assign n25283 = n24906 & n25282 ;
  assign n24091 = n9552 & n24080 ;
  assign n35754 = ~n24151 ;
  assign n24861 = n35754 & n24860 ;
  assign n25284 = n24151 & n24865 ;
  assign n25285 = n24861 | n25284 ;
  assign n25286 = n24676 & n25285 ;
  assign n25287 = n24676 | n25285 ;
  assign n35755 = ~n25286 ;
  assign n25288 = n35755 & n25287 ;
  assign n25289 = n9562 & n25288 ;
  assign n25300 = n10126 & n24151 ;
  assign n25301 = n10105 & n24676 ;
  assign n25302 = n25300 | n25301 ;
  assign n25303 = n25289 | n25302 ;
  assign n35756 = ~n25303 ;
  assign n25304 = x2 & n35756 ;
  assign n25305 = n30049 & n25303 ;
  assign n25306 = n25304 | n25305 ;
  assign n35757 = ~n24091 ;
  assign n25307 = n35757 & n25306 ;
  assign n25309 = n25283 | n25307 ;
  assign n25308 = n25283 & n25307 ;
  assign n24593 = n24214 & n24592 ;
  assign n35758 = ~n24593 ;
  assign n25310 = n35758 & n24594 ;
  assign n35759 = ~n25308 ;
  assign n25311 = n35759 & n25310 ;
  assign n35760 = ~n25311 ;
  assign n25338 = n25309 & n35760 ;
  assign n35761 = ~n25313 ;
  assign n25339 = n35761 & n25336 ;
  assign n25340 = n25338 | n25339 ;
  assign n35762 = ~n25337 ;
  assign n25341 = n35762 & n25340 ;
  assign n25342 = n24893 | n25341 ;
  assign n25343 = n24894 & n25342 ;
  assign n24850 = n9552 & n35663 ;
  assign n24780 = n24773 | n24778 ;
  assign n25346 = n24772 & n24780 ;
  assign n35763 = ~n24741 ;
  assign n24743 = n24712 & n35763 ;
  assign n25347 = n35621 & n24741 ;
  assign n25348 = n24743 | n25347 ;
  assign n25349 = n5791 | n5908 ;
  assign n25350 = n679 | n25349 ;
  assign n25351 = n249 | n2477 ;
  assign n25352 = n5859 | n25351 ;
  assign n35764 = ~n25352 ;
  assign n25353 = n5828 & n35764 ;
  assign n35765 = ~n25350 ;
  assign n25354 = n35765 & n25353 ;
  assign n25355 = n25348 & n25354 ;
  assign n25356 = n25348 | n25354 ;
  assign n35766 = ~n25355 ;
  assign n25357 = n35766 & n25356 ;
  assign n15190 = n889 & n32875 ;
  assign n25358 = n3328 & n32856 ;
  assign n25359 = n3343 & n32876 ;
  assign n25360 = n25358 | n25359 ;
  assign n25361 = n15190 | n25360 ;
  assign n35767 = ~n25361 ;
  assign n25362 = n25357 & n35767 ;
  assign n35768 = ~n25357 ;
  assign n25363 = n35768 & n25361 ;
  assign n25364 = n25362 | n25363 ;
  assign n35769 = ~n25364 ;
  assign n25365 = n25346 & n35769 ;
  assign n35770 = ~n25346 ;
  assign n25366 = n35770 & n25364 ;
  assign n25367 = n25365 | n25366 ;
  assign n15521 = n895 & n15516 ;
  assign n25368 = n894 | n2849 ;
  assign n25369 = n2861 & n32890 ;
  assign n25370 = n25368 | n25369 ;
  assign n25371 = n15521 | n25370 ;
  assign n25372 = x29 | n25371 ;
  assign n25373 = x29 & n25371 ;
  assign n35771 = ~n25373 ;
  assign n25374 = n25372 & n35771 ;
  assign n25375 = n25367 & n25374 ;
  assign n25376 = n25367 | n25374 ;
  assign n35772 = ~n25375 ;
  assign n25377 = n35772 & n25376 ;
  assign n25378 = n24782 | n24785 ;
  assign n35773 = ~n24789 ;
  assign n25379 = n24788 & n35773 ;
  assign n35774 = ~n25379 ;
  assign n25380 = n25378 & n35774 ;
  assign n35775 = ~n25377 ;
  assign n25381 = n35775 & n25380 ;
  assign n35776 = ~n25380 ;
  assign n25382 = n25377 & n35776 ;
  assign n25383 = n25381 | n25382 ;
  assign n24804 = n24792 & n24802 ;
  assign n25384 = n24801 | n24804 ;
  assign n35777 = ~n25384 ;
  assign n25385 = n25383 & n35777 ;
  assign n35778 = ~n25383 ;
  assign n25386 = n35778 & n25384 ;
  assign n25387 = n25385 | n25386 ;
  assign n25388 = n24762 | n24810 ;
  assign n25389 = n24811 & n25388 ;
  assign n25390 = n25387 | n25389 ;
  assign n25392 = n25387 & n25389 ;
  assign n35779 = ~n25392 ;
  assign n25393 = n25390 & n35779 ;
  assign n35780 = ~n24864 ;
  assign n25344 = n24838 & n35780 ;
  assign n35781 = ~n25344 ;
  assign n25345 = n24815 & n35781 ;
  assign n25415 = n35663 & n24867 ;
  assign n25416 = n24815 | n25415 ;
  assign n35782 = ~n25345 ;
  assign n25417 = n35782 & n25416 ;
  assign n35783 = ~n25417 ;
  assign n25418 = n25393 & n35783 ;
  assign n35784 = ~n25393 ;
  assign n25419 = n35784 & n25416 ;
  assign n25420 = n35782 & n25419 ;
  assign n25421 = n25418 | n25420 ;
  assign n35785 = ~n25421 ;
  assign n25422 = n9562 & n35785 ;
  assign n25433 = n10126 & n24815 ;
  assign n25434 = n10105 & n35784 ;
  assign n25435 = n25433 | n25434 ;
  assign n25436 = n25422 | n25435 ;
  assign n35786 = ~n25436 ;
  assign n25437 = x2 & n35786 ;
  assign n25438 = n30049 & n25436 ;
  assign n25439 = n25437 | n25438 ;
  assign n35787 = ~n24850 ;
  assign n25440 = n35787 & n25439 ;
  assign n25442 = n25343 | n25440 ;
  assign n20871 = n4135 & n20863 ;
  assign n19804 = n4148 & n34355 ;
  assign n19841 = n4185 & n19824 ;
  assign n25443 = n19804 | n19841 ;
  assign n25444 = n4165 & n34536 ;
  assign n25445 = n25443 | n25444 ;
  assign n25446 = n20871 | n25445 ;
  assign n25447 = x23 | n25446 ;
  assign n25448 = x23 & n25446 ;
  assign n35788 = ~n25448 ;
  assign n25449 = n25447 & n35788 ;
  assign n25450 = n20739 & n20743 ;
  assign n25451 = n20738 | n25450 ;
  assign n25452 = n294 | n1831 ;
  assign n25453 = n3460 | n25452 ;
  assign n25454 = n1528 | n1688 ;
  assign n25455 = n4302 | n25454 ;
  assign n25456 = n248 | n380 ;
  assign n25457 = n477 | n25456 ;
  assign n25458 = n150 | n900 ;
  assign n25459 = n25457 | n25458 ;
  assign n25460 = n25455 | n25459 ;
  assign n25461 = n25453 | n25460 ;
  assign n25462 = n23108 | n25461 ;
  assign n25463 = n23083 | n23954 ;
  assign n25464 = n25462 | n25463 ;
  assign n35789 = ~n25464 ;
  assign n25465 = n13489 & n35789 ;
  assign n35790 = ~n25451 ;
  assign n25466 = n35790 & n25465 ;
  assign n35791 = ~n25465 ;
  assign n25467 = n25451 & n35791 ;
  assign n25468 = n25466 | n25467 ;
  assign n20290 = n889 & n34383 ;
  assign n19972 = n3329 & n34372 ;
  assign n20021 = n3311 & n19991 ;
  assign n25469 = n19972 | n20021 ;
  assign n25470 = n3343 & n34381 ;
  assign n25471 = n25469 | n25470 ;
  assign n25472 = n20290 | n25471 ;
  assign n25473 = n25468 | n25472 ;
  assign n25474 = n25468 & n25472 ;
  assign n35792 = ~n25474 ;
  assign n25475 = n25473 & n35792 ;
  assign n20321 = n895 & n20311 ;
  assign n19915 = n2849 & n19893 ;
  assign n19932 = n2861 & n19917 ;
  assign n25476 = n19915 | n19932 ;
  assign n25477 = n894 & n19870 ;
  assign n25478 = n25476 | n25477 ;
  assign n25479 = n20321 | n25478 ;
  assign n25480 = x29 | n25479 ;
  assign n25481 = x29 & n25479 ;
  assign n35793 = ~n25481 ;
  assign n25482 = n25480 & n35793 ;
  assign n35794 = ~n25475 ;
  assign n25483 = n35794 & n25482 ;
  assign n35795 = ~n25482 ;
  assign n25484 = n25475 & n35795 ;
  assign n25485 = n25483 | n25484 ;
  assign n25486 = n20754 | n20759 ;
  assign n25487 = n25485 | n25486 ;
  assign n25488 = n25485 & n25486 ;
  assign n35796 = ~n25488 ;
  assign n25489 = n25487 & n35796 ;
  assign n20549 = n3791 & n34450 ;
  assign n19866 = n209 & n19846 ;
  assign n20088 = n3802 & n20067 ;
  assign n25490 = n19866 | n20088 ;
  assign n25491 = n3818 & n34452 ;
  assign n25492 = n25490 | n25491 ;
  assign n25493 = n20549 | n25492 ;
  assign n25494 = x26 | n25493 ;
  assign n25495 = x26 & n25493 ;
  assign n35797 = ~n25495 ;
  assign n25496 = n25494 & n35797 ;
  assign n35798 = ~n25489 ;
  assign n25497 = n35798 & n25496 ;
  assign n35799 = ~n25496 ;
  assign n25498 = n25489 & n35799 ;
  assign n25499 = n25497 | n25498 ;
  assign n35800 = ~n20766 ;
  assign n25500 = n20764 & n35800 ;
  assign n35801 = ~n25500 ;
  assign n25501 = n20763 & n35801 ;
  assign n25502 = n25499 & n25501 ;
  assign n25503 = n25499 | n25501 ;
  assign n35802 = ~n25502 ;
  assign n25504 = n35802 & n25503 ;
  assign n25505 = n25449 & n25504 ;
  assign n25506 = n25449 | n25504 ;
  assign n35803 = ~n25505 ;
  assign n25507 = n35803 & n25506 ;
  assign n35804 = ~n20710 ;
  assign n25508 = n35804 & n20797 ;
  assign n35805 = ~n25508 ;
  assign n25509 = n20796 & n35805 ;
  assign n35806 = ~n25507 ;
  assign n25510 = n35806 & n25509 ;
  assign n35807 = ~n25509 ;
  assign n25511 = n25507 & n35807 ;
  assign n25512 = n25510 | n25511 ;
  assign n21102 = n4686 & n34603 ;
  assign n19745 = n4706 & n34520 ;
  assign n19754 = n4726 & n19752 ;
  assign n25513 = n19745 | n19754 ;
  assign n25514 = n4748 & n34596 ;
  assign n25515 = n25513 | n25514 ;
  assign n25516 = n21102 | n25515 ;
  assign n25517 = x20 | n25516 ;
  assign n25518 = x20 & n25516 ;
  assign n35808 = ~n25518 ;
  assign n25519 = n25517 & n35808 ;
  assign n35809 = ~n25512 ;
  assign n25520 = n35809 & n25519 ;
  assign n35810 = ~n25519 ;
  assign n25521 = n25512 & n35810 ;
  assign n25522 = n25520 | n25521 ;
  assign n25523 = n20800 | n20823 ;
  assign n35811 = ~n21061 ;
  assign n25524 = n35811 & n25523 ;
  assign n35812 = ~n25522 ;
  assign n25525 = n35812 & n25524 ;
  assign n35813 = ~n25524 ;
  assign n25526 = n25522 & n35813 ;
  assign n25527 = n25525 | n25526 ;
  assign n21874 = n37300 & n34817 ;
  assign n19671 = n5144 & n34360 ;
  assign n19697 = n5166 & n34349 ;
  assign n25528 = n19671 | n19697 ;
  assign n25529 = n5191 & n34803 ;
  assign n25530 = n25528 | n25529 ;
  assign n25531 = n21874 | n25530 ;
  assign n25532 = x17 | n25531 ;
  assign n25533 = x17 & n25531 ;
  assign n35814 = ~n25533 ;
  assign n25534 = n25532 & n35814 ;
  assign n35815 = ~n21341 ;
  assign n25535 = n21338 & n35815 ;
  assign n25536 = n25534 & n25535 ;
  assign n25537 = n25534 | n25535 ;
  assign n35816 = ~n25536 ;
  assign n25538 = n35816 & n25537 ;
  assign n25539 = n25527 & n25538 ;
  assign n25540 = n25527 | n25538 ;
  assign n35817 = ~n25539 ;
  assign n25541 = n35817 & n25540 ;
  assign n22649 = n5937 & n35035 ;
  assign n21730 = n5970 & n21729 ;
  assign n21805 = n5994 & n21753 ;
  assign n25542 = n21730 | n21805 ;
  assign n25543 = n6018 & n35018 ;
  assign n25544 = n25542 | n25543 ;
  assign n25545 = n22649 | n25544 ;
  assign n25546 = x14 | n25545 ;
  assign n25547 = x14 & n25545 ;
  assign n35818 = ~n25547 ;
  assign n25548 = n25546 & n35818 ;
  assign n25549 = n25541 & n25548 ;
  assign n25550 = n25541 | n25548 ;
  assign n35819 = ~n25549 ;
  assign n25551 = n35819 & n25550 ;
  assign n35820 = ~n22152 ;
  assign n25552 = n21836 & n35820 ;
  assign n25553 = n25551 | n25552 ;
  assign n25554 = n25551 & n25552 ;
  assign n35821 = ~n25554 ;
  assign n25555 = n25553 & n35821 ;
  assign n23440 = n6272 & n35262 ;
  assign n22514 = n6190 & n35020 ;
  assign n22582 = n6244 & n22533 ;
  assign n25556 = n22514 | n22582 ;
  assign n25557 = n6217 & n23444 ;
  assign n25558 = n25556 | n25557 ;
  assign n25559 = n23440 | n25558 ;
  assign n25560 = x11 | n25559 ;
  assign n25561 = x11 & n25559 ;
  assign n35822 = ~n25561 ;
  assign n25562 = n25560 & n35822 ;
  assign n35823 = ~n25555 ;
  assign n25563 = n35823 & n25562 ;
  assign n35824 = ~n25562 ;
  assign n25564 = n25555 & n35824 ;
  assign n25565 = n25563 | n25564 ;
  assign n35825 = ~n22966 ;
  assign n25566 = n22610 & n35825 ;
  assign n35826 = ~n25566 ;
  assign n25567 = n22609 & n35826 ;
  assign n25568 = n25565 & n25567 ;
  assign n25569 = n25565 | n25567 ;
  assign n35827 = ~n25568 ;
  assign n25570 = n35827 & n25569 ;
  assign n24196 = n7068 & n35472 ;
  assign n23294 = n69 & n35467 ;
  assign n23326 = n7041 & n35244 ;
  assign n25571 = n23294 | n23326 ;
  assign n25572 = n7017 & n35465 ;
  assign n25573 = n25571 | n25572 ;
  assign n25574 = n24196 | n25573 ;
  assign n25575 = x8 | n25574 ;
  assign n25576 = x8 & n25574 ;
  assign n35828 = ~n25576 ;
  assign n25577 = n25575 & n35828 ;
  assign n25578 = n25570 & n25577 ;
  assign n25579 = n25570 | n25577 ;
  assign n35829 = ~n25578 ;
  assign n25580 = n35829 & n25579 ;
  assign n35830 = ~n23797 ;
  assign n25581 = n23395 & n35830 ;
  assign n35831 = ~n25581 ;
  assign n25582 = n23394 & n35831 ;
  assign n25583 = n25580 | n25582 ;
  assign n25584 = n25580 & n25582 ;
  assign n35832 = ~n25584 ;
  assign n25585 = n25583 & n35832 ;
  assign n25290 = n8157 & n25288 ;
  assign n24071 = n740 & n24057 ;
  assign n24086 = n8195 & n24080 ;
  assign n25586 = n24071 | n24086 ;
  assign n25587 = n9052 & n24676 ;
  assign n25588 = n25586 | n25587 ;
  assign n25589 = n25290 | n25588 ;
  assign n25590 = x5 | n25589 ;
  assign n25591 = x5 & n25589 ;
  assign n35833 = ~n25591 ;
  assign n25592 = n25590 & n35833 ;
  assign n25593 = n25585 & n25592 ;
  assign n25594 = n25585 | n25592 ;
  assign n35834 = ~n25593 ;
  assign n25595 = n35834 & n25594 ;
  assign n35835 = ~n24602 ;
  assign n25596 = n24161 & n35835 ;
  assign n35836 = ~n25596 ;
  assign n25597 = n24160 & n35836 ;
  assign n35837 = ~n25595 ;
  assign n25598 = n35837 & n25597 ;
  assign n35838 = ~n25597 ;
  assign n25599 = n25595 & n35838 ;
  assign n25600 = n25598 | n25599 ;
  assign n25441 = n25343 & n25440 ;
  assign n35839 = ~n25441 ;
  assign n25601 = n35839 & n25442 ;
  assign n25602 = n25600 & n25601 ;
  assign n35840 = ~n25602 ;
  assign n25603 = n25442 & n35840 ;
  assign n25604 = n956 | n971 ;
  assign n25605 = n1200 | n1565 ;
  assign n25606 = n25604 | n25605 ;
  assign n25607 = n1799 | n25606 ;
  assign n25608 = n11241 | n25607 ;
  assign n25609 = n528 | n868 ;
  assign n25610 = n697 | n25609 ;
  assign n25611 = n1141 | n25610 ;
  assign n25612 = n12766 | n25611 ;
  assign n35841 = ~n25612 ;
  assign n25613 = n22219 & n35841 ;
  assign n35842 = ~n25608 ;
  assign n25614 = n35842 & n25613 ;
  assign n35843 = ~n11133 ;
  assign n25615 = n35843 & n25614 ;
  assign n35844 = ~n22193 ;
  assign n25616 = n35844 & n25615 ;
  assign n20422 = n889 & n20412 ;
  assign n19958 = n3329 & n34381 ;
  assign n19990 = n3311 & n34372 ;
  assign n25617 = n19958 | n19990 ;
  assign n25618 = n3343 & n19917 ;
  assign n25619 = n25617 | n25618 ;
  assign n25620 = n20422 | n25619 ;
  assign n35845 = ~n25620 ;
  assign n25621 = n25616 & n35845 ;
  assign n35846 = ~n25616 ;
  assign n25622 = n35846 & n25620 ;
  assign n25623 = n25621 | n25622 ;
  assign n35847 = ~n25468 ;
  assign n25624 = n35847 & n25472 ;
  assign n25625 = n25467 | n25624 ;
  assign n25626 = n25623 | n25625 ;
  assign n25627 = n25623 & n25625 ;
  assign n35848 = ~n25627 ;
  assign n25628 = n25626 & n35848 ;
  assign n35849 = ~n25485 ;
  assign n25629 = n35849 & n25486 ;
  assign n25630 = n25483 | n25629 ;
  assign n35850 = ~n25630 ;
  assign n25631 = n25628 & n35850 ;
  assign n35851 = ~n25628 ;
  assign n25632 = n35851 & n25630 ;
  assign n25633 = n25631 | n25632 ;
  assign n20495 = n895 & n20486 ;
  assign n19882 = n2849 & n19870 ;
  assign n19895 = n2861 & n19893 ;
  assign n25634 = n19882 | n19895 ;
  assign n25635 = n894 & n19846 ;
  assign n25636 = n25634 | n25635 ;
  assign n25637 = n20495 | n25636 ;
  assign n35852 = ~n25637 ;
  assign n25638 = x29 & n35852 ;
  assign n25639 = n30024 & n25637 ;
  assign n25640 = n25638 | n25639 ;
  assign n25641 = n25633 | n25640 ;
  assign n25642 = n25633 & n25640 ;
  assign n35853 = ~n25642 ;
  assign n25643 = n25641 & n35853 ;
  assign n20524 = n3791 & n34442 ;
  assign n20069 = n209 & n20067 ;
  assign n20111 = n3802 & n34354 ;
  assign n25644 = n20069 | n20111 ;
  assign n25645 = n3818 & n20527 ;
  assign n25646 = n25644 | n25645 ;
  assign n25647 = n20524 | n25646 ;
  assign n25648 = x26 | n25647 ;
  assign n25649 = x26 & n25647 ;
  assign n35854 = ~n25649 ;
  assign n25650 = n25648 & n35854 ;
  assign n25651 = n25643 & n25650 ;
  assign n25652 = n25643 | n25650 ;
  assign n35855 = ~n25651 ;
  assign n25653 = n35855 & n25652 ;
  assign n35856 = ~n25498 ;
  assign n25654 = n35856 & n25503 ;
  assign n35857 = ~n25653 ;
  assign n25655 = n35857 & n25654 ;
  assign n35858 = ~n25654 ;
  assign n25656 = n25653 & n35858 ;
  assign n25657 = n25655 | n25656 ;
  assign n20842 = n4135 & n20833 ;
  assign n19791 = n4148 & n34519 ;
  assign n19818 = n4185 & n34355 ;
  assign n25658 = n19791 | n19818 ;
  assign n25659 = n4165 & n20845 ;
  assign n25660 = n25658 | n25659 ;
  assign n25661 = n20842 | n25660 ;
  assign n25662 = x23 | n25661 ;
  assign n25663 = x23 & n25661 ;
  assign n35859 = ~n25663 ;
  assign n25664 = n25662 & n35859 ;
  assign n35860 = ~n25657 ;
  assign n25665 = n35860 & n25664 ;
  assign n35861 = ~n25664 ;
  assign n25666 = n25657 & n35861 ;
  assign n25667 = n25665 | n25666 ;
  assign n35862 = ~n25504 ;
  assign n25668 = n25449 & n35862 ;
  assign n25669 = n25510 | n25668 ;
  assign n25670 = n25667 | n25669 ;
  assign n25671 = n25667 & n25669 ;
  assign n35863 = ~n25671 ;
  assign n25672 = n25670 & n35863 ;
  assign n21078 = n4686 & n34598 ;
  assign n19724 = n4706 & n34363 ;
  assign n19746 = n4726 & n34520 ;
  assign n25673 = n19724 | n19746 ;
  assign n25674 = n4748 & n34349 ;
  assign n25675 = n25673 | n25674 ;
  assign n25676 = n21078 | n25675 ;
  assign n25677 = x20 | n25676 ;
  assign n25678 = x20 & n25676 ;
  assign n35864 = ~n25678 ;
  assign n25679 = n25677 & n35864 ;
  assign n25680 = n25672 & n25679 ;
  assign n25681 = n25672 | n25679 ;
  assign n35865 = ~n25680 ;
  assign n25682 = n35865 & n25681 ;
  assign n25683 = n25522 | n25524 ;
  assign n35866 = ~n25521 ;
  assign n25684 = n35866 & n25683 ;
  assign n35867 = ~n25682 ;
  assign n25685 = n35867 & n25684 ;
  assign n35868 = ~n25684 ;
  assign n25686 = n25682 & n35868 ;
  assign n25687 = n25685 | n25686 ;
  assign n21855 = n37300 & n21848 ;
  assign n19672 = n5166 & n34360 ;
  assign n21759 = n5144 & n34803 ;
  assign n25688 = n19672 | n21759 ;
  assign n25689 = n5191 & n21753 ;
  assign n25690 = n25688 | n25689 ;
  assign n25691 = n21855 | n25690 ;
  assign n25692 = x17 | n25691 ;
  assign n25693 = x17 & n25691 ;
  assign n35869 = ~n25693 ;
  assign n25694 = n25692 & n35869 ;
  assign n25695 = n25537 & n35817 ;
  assign n25696 = n25694 & n25695 ;
  assign n25697 = n25694 | n25695 ;
  assign n35870 = ~n25696 ;
  assign n25698 = n35870 & n25697 ;
  assign n35871 = ~n25687 ;
  assign n25699 = n35871 & n25698 ;
  assign n35872 = ~n25698 ;
  assign n25700 = n25687 & n35872 ;
  assign n25701 = n25699 | n25700 ;
  assign n22626 = n5937 & n35030 ;
  assign n21733 = n5994 & n21729 ;
  assign n22551 = n5970 & n35018 ;
  assign n25702 = n21733 | n22551 ;
  assign n25703 = n6018 & n22533 ;
  assign n25704 = n25702 | n25703 ;
  assign n25705 = n22626 | n25704 ;
  assign n25706 = x14 | n25705 ;
  assign n25707 = x14 & n25705 ;
  assign n35873 = ~n25707 ;
  assign n25708 = n25706 & n35873 ;
  assign n35874 = ~n25548 ;
  assign n25709 = n25541 & n35874 ;
  assign n35875 = ~n25709 ;
  assign n25710 = n25553 & n35875 ;
  assign n25711 = n25708 & n25710 ;
  assign n25712 = n25708 | n25710 ;
  assign n35876 = ~n25711 ;
  assign n25713 = n35876 & n25712 ;
  assign n25714 = n25701 & n25713 ;
  assign n25715 = n25701 | n25713 ;
  assign n35877 = ~n25714 ;
  assign n25716 = n35877 & n25715 ;
  assign n23404 = n6272 & n35252 ;
  assign n22515 = n6244 & n35020 ;
  assign n23346 = n6190 & n23339 ;
  assign n25717 = n22515 | n23346 ;
  assign n25718 = n6217 & n35254 ;
  assign n25719 = n25717 | n25718 ;
  assign n25720 = n23404 | n25719 ;
  assign n25721 = x11 | n25720 ;
  assign n25722 = x11 & n25720 ;
  assign n35878 = ~n25722 ;
  assign n25723 = n25721 & n35878 ;
  assign n25724 = n25716 & n25723 ;
  assign n25725 = n25716 | n25723 ;
  assign n35879 = ~n25724 ;
  assign n25726 = n35879 & n25725 ;
  assign n35880 = ~n25564 ;
  assign n25727 = n35880 & n25569 ;
  assign n25728 = n25726 | n25727 ;
  assign n25729 = n25726 & n25727 ;
  assign n35881 = ~n25729 ;
  assign n25730 = n25728 & n35881 ;
  assign n24171 = n7068 & n24168 ;
  assign n23292 = n7041 & n35467 ;
  assign n24114 = n69 & n35458 ;
  assign n25731 = n23292 | n24114 ;
  assign n25732 = n7017 & n24080 ;
  assign n25733 = n25731 | n25732 ;
  assign n25734 = n24171 | n25733 ;
  assign n25735 = x8 | n25734 ;
  assign n25736 = x8 & n25734 ;
  assign n35882 = ~n25736 ;
  assign n25737 = n25735 & n35882 ;
  assign n35883 = ~n25730 ;
  assign n25738 = n35883 & n25737 ;
  assign n35884 = ~n25737 ;
  assign n25739 = n25730 & n35884 ;
  assign n25740 = n25738 | n25739 ;
  assign n35885 = ~n25577 ;
  assign n25741 = n25570 & n35885 ;
  assign n35886 = ~n25741 ;
  assign n25742 = n25583 & n35886 ;
  assign n35887 = ~n25740 ;
  assign n25743 = n35887 & n25742 ;
  assign n35888 = ~n25742 ;
  assign n25744 = n25740 & n35888 ;
  assign n25745 = n25743 | n25744 ;
  assign n25320 = n8157 & n35670 ;
  assign n24067 = n8195 & n24057 ;
  assign n24683 = n740 & n24676 ;
  assign n25746 = n24067 | n24683 ;
  assign n25747 = n9052 & n35663 ;
  assign n25748 = n25746 | n25747 ;
  assign n25749 = n25320 | n25748 ;
  assign n25750 = x5 | n25749 ;
  assign n25751 = x5 & n25749 ;
  assign n35889 = ~n25751 ;
  assign n25752 = n25750 & n35889 ;
  assign n35890 = ~n25745 ;
  assign n25753 = n35890 & n25752 ;
  assign n35891 = ~n25752 ;
  assign n25754 = n25745 & n35891 ;
  assign n25755 = n25753 | n25754 ;
  assign n35892 = ~n25585 ;
  assign n25756 = n35892 & n25592 ;
  assign n25757 = n25598 | n25756 ;
  assign n35893 = ~n25757 ;
  assign n25758 = n25755 & n35893 ;
  assign n35894 = ~n25755 ;
  assign n25759 = n35894 & n25757 ;
  assign n25760 = n25758 | n25759 ;
  assign n24827 = n9552 & n24815 ;
  assign n25761 = n24712 & n24741 ;
  assign n25762 = n25355 | n25761 ;
  assign n25763 = n5787 | n5847 ;
  assign n25764 = n25350 | n25763 ;
  assign n25765 = n25762 | n25764 ;
  assign n25767 = n25762 & n25764 ;
  assign n35895 = ~n25767 ;
  assign n25768 = n25765 & n35895 ;
  assign n15275 = n889 & n32889 ;
  assign n15086 = n3311 & n15081 ;
  assign n15175 = n3329 & n32876 ;
  assign n25769 = n15086 | n15175 ;
  assign n25770 = n3343 & n32890 ;
  assign n25771 = n25769 | n25770 ;
  assign n25772 = n15275 | n25771 ;
  assign n35896 = ~n25772 ;
  assign n25773 = n25768 & n35896 ;
  assign n35897 = ~n25768 ;
  assign n25774 = n35897 & n25772 ;
  assign n25775 = n25773 | n25774 ;
  assign n25776 = x26 | n98 ;
  assign n25777 = n30024 & n25776 ;
  assign n25778 = n14311 | n25777 ;
  assign n35898 = ~n25778 ;
  assign n25779 = n25775 & n35898 ;
  assign n35899 = ~n25775 ;
  assign n25780 = n35899 & n25778 ;
  assign n25781 = n25779 | n25780 ;
  assign n25782 = n25346 | n25364 ;
  assign n35900 = ~n25362 ;
  assign n25783 = n35900 & n25782 ;
  assign n25784 = n25781 & n25783 ;
  assign n25785 = n25781 | n25783 ;
  assign n35901 = ~n25784 ;
  assign n25786 = n35901 & n25785 ;
  assign n35902 = ~n25374 ;
  assign n25787 = n25367 & n35902 ;
  assign n25788 = n25377 | n25380 ;
  assign n35903 = ~n25787 ;
  assign n25789 = n35903 & n25788 ;
  assign n25790 = n25786 & n25789 ;
  assign n25791 = n25786 | n25789 ;
  assign n35904 = ~n25790 ;
  assign n25792 = n35904 & n25791 ;
  assign n25391 = n25386 | n25389 ;
  assign n35905 = ~n25385 ;
  assign n25793 = n35905 & n25391 ;
  assign n25794 = n25792 & n25793 ;
  assign n25795 = n25792 | n25793 ;
  assign n35906 = ~n25794 ;
  assign n25796 = n35906 & n25795 ;
  assign n25810 = n35784 & n25796 ;
  assign n35907 = ~n25796 ;
  assign n25818 = n25393 & n35907 ;
  assign n25819 = n25810 | n25818 ;
  assign n25820 = n25345 | n25419 ;
  assign n35908 = ~n25820 ;
  assign n25821 = n25819 & n35908 ;
  assign n35909 = ~n25819 ;
  assign n25823 = n35909 & n25820 ;
  assign n25824 = n25821 | n25823 ;
  assign n35910 = ~n25824 ;
  assign n25825 = n9562 & n35910 ;
  assign n25836 = n10126 & n35784 ;
  assign n25837 = n10105 & n25796 ;
  assign n25838 = n25836 | n25837 ;
  assign n25839 = n25825 | n25838 ;
  assign n35911 = ~n25839 ;
  assign n25840 = x2 & n35911 ;
  assign n25841 = n30049 & n25839 ;
  assign n25842 = n25840 | n25841 ;
  assign n35912 = ~n24827 ;
  assign n25843 = n35912 & n25842 ;
  assign n35913 = ~n25760 ;
  assign n25844 = n35913 & n25843 ;
  assign n35914 = ~n25843 ;
  assign n25845 = n25760 & n35914 ;
  assign n25846 = n25844 | n25845 ;
  assign n25847 = n25603 & n25846 ;
  assign n25848 = n25603 | n25846 ;
  assign n35915 = ~n25847 ;
  assign n25849 = n35915 & n25848 ;
  assign n25850 = n25600 | n25601 ;
  assign n25851 = n35840 & n25850 ;
  assign n25852 = n25849 & n25851 ;
  assign n25853 = n25849 | n25851 ;
  assign n35916 = ~n25852 ;
  assign n33 = n35916 & n25853 ;
  assign n22571 = n5937 & n35022 ;
  assign n22545 = n5994 & n35018 ;
  assign n22581 = n5970 & n22533 ;
  assign n25854 = n22545 | n22581 ;
  assign n25855 = n6018 & n35020 ;
  assign n25856 = n25854 | n25855 ;
  assign n25857 = n22571 | n25856 ;
  assign n25858 = x14 | n25857 ;
  assign n25859 = x14 & n25857 ;
  assign n35917 = ~n25859 ;
  assign n25860 = n25858 & n35917 ;
  assign n35918 = ~n25666 ;
  assign n25861 = n35918 & n25670 ;
  assign n35919 = ~n25621 ;
  assign n25862 = n35919 & n25626 ;
  assign n20352 = n889 & n34399 ;
  assign n19934 = n3329 & n19917 ;
  assign n19963 = n3311 & n34381 ;
  assign n25863 = n19934 | n19963 ;
  assign n25864 = n3343 & n19893 ;
  assign n25865 = n25863 | n25864 ;
  assign n25866 = n20352 | n25865 ;
  assign n35920 = ~n25866 ;
  assign n25867 = n25862 & n35920 ;
  assign n35921 = ~n25862 ;
  assign n25868 = n35921 & n25866 ;
  assign n25869 = n25867 | n25868 ;
  assign n25870 = n1952 | n4608 ;
  assign n25871 = n157 | n1389 ;
  assign n25872 = n234 | n1472 ;
  assign n25873 = n25871 | n25872 ;
  assign n25874 = n25870 | n25873 ;
  assign n25875 = n558 | n25874 ;
  assign n25876 = n2359 | n25875 ;
  assign n25877 = n309 | n811 ;
  assign n25878 = n795 | n865 ;
  assign n25879 = n25877 | n25878 ;
  assign n25880 = n1538 | n25879 ;
  assign n35922 = ~n2394 ;
  assign n25881 = n35922 & n11669 ;
  assign n35923 = ~n25880 ;
  assign n25882 = n35923 & n25881 ;
  assign n35924 = ~n5422 ;
  assign n25883 = n35924 & n25882 ;
  assign n35925 = ~n5526 ;
  assign n25884 = n35925 & n25883 ;
  assign n35926 = ~n3045 ;
  assign n25885 = n35926 & n25884 ;
  assign n35927 = ~n25876 ;
  assign n25886 = n35927 & n25885 ;
  assign n25887 = n25869 & n25886 ;
  assign n25888 = n25869 | n25886 ;
  assign n35928 = ~n25887 ;
  assign n25889 = n35928 & n25888 ;
  assign n20590 = n895 & n20579 ;
  assign n19867 = n2849 & n19846 ;
  assign n19878 = n2861 & n19870 ;
  assign n25890 = n19867 | n19878 ;
  assign n25891 = n894 & n20067 ;
  assign n25892 = n25890 | n25891 ;
  assign n25893 = n20590 | n25892 ;
  assign n25894 = x29 | n25893 ;
  assign n25895 = x29 & n25893 ;
  assign n35929 = ~n25895 ;
  assign n25896 = n25894 & n35929 ;
  assign n35930 = ~n25889 ;
  assign n25897 = n35930 & n25896 ;
  assign n35931 = ~n25896 ;
  assign n25898 = n25889 & n35931 ;
  assign n25899 = n25897 | n25898 ;
  assign n35932 = ~n25631 ;
  assign n25900 = n35932 & n25641 ;
  assign n35933 = ~n25899 ;
  assign n25901 = n35933 & n25900 ;
  assign n35934 = ~n25900 ;
  assign n25902 = n25899 & n35934 ;
  assign n25903 = n25901 | n25902 ;
  assign n20785 = n3791 & n34511 ;
  assign n19842 = n3802 & n19824 ;
  assign n20112 = n209 & n34354 ;
  assign n25904 = n19842 | n20112 ;
  assign n25905 = n3818 & n34513 ;
  assign n25906 = n25904 | n25905 ;
  assign n25907 = n20785 | n25906 ;
  assign n25908 = x26 | n25907 ;
  assign n25909 = x26 & n25907 ;
  assign n35935 = ~n25909 ;
  assign n25910 = n25908 & n35935 ;
  assign n35936 = ~n25903 ;
  assign n25911 = n35936 & n25910 ;
  assign n35937 = ~n25910 ;
  assign n25912 = n25903 & n35937 ;
  assign n25913 = n25911 | n25912 ;
  assign n35938 = ~n25643 ;
  assign n25914 = n35938 & n25650 ;
  assign n25915 = n25655 | n25914 ;
  assign n25916 = n25913 | n25915 ;
  assign n25917 = n25913 & n25915 ;
  assign n35939 = ~n25917 ;
  assign n25918 = n25916 & n35939 ;
  assign n20814 = n4135 & n20805 ;
  assign n19768 = n4148 & n19752 ;
  assign n19793 = n4185 & n34519 ;
  assign n25919 = n19768 | n19793 ;
  assign n25920 = n4165 & n34520 ;
  assign n25921 = n25919 | n25920 ;
  assign n25922 = n20814 | n25921 ;
  assign n25923 = x23 | n25922 ;
  assign n25924 = x23 & n25922 ;
  assign n35940 = ~n25924 ;
  assign n25925 = n25923 & n35940 ;
  assign n35941 = ~n25918 ;
  assign n25926 = n35941 & n25925 ;
  assign n35942 = ~n25925 ;
  assign n25927 = n25918 & n35942 ;
  assign n25928 = n25926 | n25927 ;
  assign n35943 = ~n25928 ;
  assign n25929 = n25861 & n35943 ;
  assign n35944 = ~n25861 ;
  assign n25930 = n35944 & n25928 ;
  assign n25931 = n25929 | n25930 ;
  assign n20157 = n4686 & n34362 ;
  assign n19684 = n4706 & n34349 ;
  assign n19715 = n4726 & n34363 ;
  assign n25932 = n19684 | n19715 ;
  assign n25933 = n4748 & n34365 ;
  assign n25934 = n25932 | n25933 ;
  assign n25935 = n20157 | n25934 ;
  assign n25936 = x20 | n25935 ;
  assign n25937 = x20 & n25935 ;
  assign n35945 = ~n25937 ;
  assign n25938 = n25936 & n35945 ;
  assign n25939 = n25931 & n25938 ;
  assign n25940 = n25931 | n25938 ;
  assign n35946 = ~n25939 ;
  assign n25941 = n35946 & n25940 ;
  assign n35947 = ~n25672 ;
  assign n25942 = n35947 & n25679 ;
  assign n25943 = n25685 | n25942 ;
  assign n25944 = n25941 | n25943 ;
  assign n25945 = n25941 & n25943 ;
  assign n35948 = ~n25945 ;
  assign n25946 = n25944 & n35948 ;
  assign n21797 = n37300 & n34802 ;
  assign n21768 = n5166 & n34803 ;
  assign n21811 = n5144 & n21753 ;
  assign n25947 = n21768 | n21811 ;
  assign n25948 = n5191 & n21804 ;
  assign n25949 = n25947 | n25948 ;
  assign n25950 = n21797 | n25949 ;
  assign n25951 = x17 | n25950 ;
  assign n25952 = x17 & n25950 ;
  assign n35949 = ~n25952 ;
  assign n25953 = n25951 & n35949 ;
  assign n35950 = ~n25946 ;
  assign n25954 = n35950 & n25953 ;
  assign n35951 = ~n25953 ;
  assign n25955 = n25946 & n35951 ;
  assign n25956 = n25954 | n25955 ;
  assign n25957 = n25687 & n25698 ;
  assign n35952 = ~n25957 ;
  assign n25958 = n25697 & n35952 ;
  assign n25959 = n25956 & n25958 ;
  assign n25960 = n25956 | n25958 ;
  assign n35953 = ~n25959 ;
  assign n25961 = n35953 & n25960 ;
  assign n35954 = ~n25961 ;
  assign n25962 = n25860 & n35954 ;
  assign n35955 = ~n25860 ;
  assign n25963 = n35955 & n25961 ;
  assign n25964 = n25962 | n25963 ;
  assign n25965 = n25712 & n35877 ;
  assign n35956 = ~n25964 ;
  assign n25966 = n35956 & n25965 ;
  assign n35957 = ~n25965 ;
  assign n25967 = n25964 & n35957 ;
  assign n25968 = n25966 | n25967 ;
  assign n23376 = n6272 & n23372 ;
  assign n23330 = n6190 & n35244 ;
  assign n23340 = n6244 & n23339 ;
  assign n25969 = n23330 | n23340 ;
  assign n25970 = n6217 & n35246 ;
  assign n25971 = n25969 | n25970 ;
  assign n25972 = n23376 | n25971 ;
  assign n25973 = x11 | n25972 ;
  assign n25974 = x11 & n25972 ;
  assign n35958 = ~n25974 ;
  assign n25975 = n25973 & n35958 ;
  assign n35959 = ~n25968 ;
  assign n25976 = n35959 & n25975 ;
  assign n35960 = ~n25975 ;
  assign n25977 = n25968 & n35960 ;
  assign n25978 = n25976 | n25977 ;
  assign n35961 = ~n25723 ;
  assign n25979 = n25716 & n35961 ;
  assign n35962 = ~n25979 ;
  assign n25980 = n25728 & n35962 ;
  assign n35963 = ~n25978 ;
  assign n25981 = n35963 & n25980 ;
  assign n35964 = ~n25980 ;
  assign n25982 = n25978 & n35964 ;
  assign n25983 = n25981 | n25982 ;
  assign n24142 = n7068 & n35457 ;
  assign n24085 = n69 & n24080 ;
  assign n24111 = n7041 & n35458 ;
  assign n25984 = n24085 | n24111 ;
  assign n25985 = n7017 & n24151 ;
  assign n25986 = n25984 | n25985 ;
  assign n25987 = n24142 | n25986 ;
  assign n25988 = x8 | n25987 ;
  assign n25989 = x8 & n25987 ;
  assign n35965 = ~n25989 ;
  assign n25990 = n25988 & n35965 ;
  assign n35966 = ~n25983 ;
  assign n25991 = n35966 & n25990 ;
  assign n35967 = ~n25990 ;
  assign n25992 = n25983 & n35967 ;
  assign n25993 = n25991 | n25992 ;
  assign n25994 = n25738 | n25743 ;
  assign n35968 = ~n25994 ;
  assign n25995 = n25993 & n35968 ;
  assign n35969 = ~n25993 ;
  assign n25996 = n35969 & n25994 ;
  assign n25997 = n25995 | n25996 ;
  assign n24876 = n8157 & n35662 ;
  assign n24682 = n8195 & n24676 ;
  assign n24845 = n740 & n35663 ;
  assign n25998 = n24682 | n24845 ;
  assign n25999 = n9052 & n24815 ;
  assign n26000 = n25998 | n25999 ;
  assign n26001 = n24876 | n26000 ;
  assign n26002 = x5 | n26001 ;
  assign n26003 = x5 & n26001 ;
  assign n35970 = ~n26003 ;
  assign n26004 = n26002 & n35970 ;
  assign n35971 = ~n25997 ;
  assign n26005 = n35971 & n26004 ;
  assign n35972 = ~n26004 ;
  assign n26006 = n25997 & n35972 ;
  assign n26007 = n26005 | n26006 ;
  assign n26008 = n25753 | n25759 ;
  assign n35973 = ~n26007 ;
  assign n26009 = n35973 & n26008 ;
  assign n35974 = ~n26008 ;
  assign n26010 = n26007 & n35974 ;
  assign n26011 = n26009 | n26010 ;
  assign n35975 = ~n25845 ;
  assign n26012 = n35975 & n25848 ;
  assign n25408 = n9552 & n35784 ;
  assign n35976 = ~n25793 ;
  assign n26013 = n25792 & n35976 ;
  assign n35977 = ~n26013 ;
  assign n26014 = n25791 & n35977 ;
  assign n26015 = n25775 | n25778 ;
  assign n35978 = ~n25783 ;
  assign n26016 = n25781 & n35978 ;
  assign n35979 = ~n26016 ;
  assign n26017 = n26015 & n35979 ;
  assign n35980 = ~n15526 ;
  assign n15536 = n6561 & n35980 ;
  assign n26018 = n3311 & n15158 ;
  assign n35981 = ~n26018 ;
  assign n26019 = n77 & n35981 ;
  assign n35982 = ~n15536 ;
  assign n26020 = n35982 & n26019 ;
  assign n26021 = n35898 & n26020 ;
  assign n35983 = ~n26020 ;
  assign n26022 = n25778 & n35983 ;
  assign n26023 = n26021 | n26022 ;
  assign n5899 = n5792 | n5898 ;
  assign n25766 = n5899 | n25764 ;
  assign n26024 = n5899 & n25764 ;
  assign n35984 = ~n26024 ;
  assign n26025 = n25766 & n35984 ;
  assign n26026 = n25768 & n25772 ;
  assign n35985 = ~n26026 ;
  assign n26027 = n25765 & n35985 ;
  assign n35986 = ~n26025 ;
  assign n26028 = n35986 & n26027 ;
  assign n35987 = ~n26027 ;
  assign n26029 = n26025 & n35987 ;
  assign n26030 = n26028 | n26029 ;
  assign n26031 = n26023 & n26030 ;
  assign n26032 = n26023 | n26030 ;
  assign n35988 = ~n26031 ;
  assign n26033 = n35988 & n26032 ;
  assign n35989 = ~n26033 ;
  assign n26034 = n26017 & n35989 ;
  assign n35990 = ~n26017 ;
  assign n26035 = n35990 & n26033 ;
  assign n26036 = n26034 | n26035 ;
  assign n26037 = n26014 & n26036 ;
  assign n26038 = n26014 | n26036 ;
  assign n35991 = ~n26037 ;
  assign n26039 = n35991 & n26038 ;
  assign n26059 = n25419 | n25796 ;
  assign n25822 = n25393 & n35908 ;
  assign n35992 = ~n25822 ;
  assign n26061 = n25796 & n35992 ;
  assign n35993 = ~n26061 ;
  assign n26062 = n26059 & n35993 ;
  assign n26063 = n26039 & n26062 ;
  assign n26064 = n26039 | n26062 ;
  assign n35994 = ~n26063 ;
  assign n26065 = n35994 & n26064 ;
  assign n26066 = n9562 & n26065 ;
  assign n26077 = n10126 & n25796 ;
  assign n26078 = n10105 & n26039 ;
  assign n26079 = n26077 | n26078 ;
  assign n26080 = n26066 | n26079 ;
  assign n35995 = ~n26080 ;
  assign n26081 = x2 & n35995 ;
  assign n26082 = n30049 & n26080 ;
  assign n26083 = n26081 | n26082 ;
  assign n35996 = ~n25408 ;
  assign n26084 = n35996 & n26083 ;
  assign n35997 = ~n26012 ;
  assign n26085 = n35997 & n26084 ;
  assign n35998 = ~n26084 ;
  assign n26086 = n26012 & n35998 ;
  assign n26087 = n26085 | n26086 ;
  assign n26088 = n26011 & n26087 ;
  assign n26089 = n26011 | n26087 ;
  assign n35999 = ~n26088 ;
  assign n26090 = n35999 & n26089 ;
  assign n26091 = n25853 & n26090 ;
  assign n26092 = n25853 | n26090 ;
  assign n36000 = ~n26091 ;
  assign n34 = n36000 & n26092 ;
  assign n23441 = n5937 & n35262 ;
  assign n22510 = n5970 & n35020 ;
  assign n22580 = n5994 & n22533 ;
  assign n26093 = n22510 | n22580 ;
  assign n26094 = n6018 & n23444 ;
  assign n26095 = n26093 | n26094 ;
  assign n26096 = n23441 | n26095 ;
  assign n26097 = x14 | n26096 ;
  assign n26098 = x14 & n26096 ;
  assign n36001 = ~n26098 ;
  assign n26099 = n26097 & n36001 ;
  assign n26100 = n25862 & n25866 ;
  assign n36002 = ~n25886 ;
  assign n26101 = n25869 & n36002 ;
  assign n26102 = n26100 | n26101 ;
  assign n26103 = n1361 | n2305 ;
  assign n26104 = n13659 | n26103 ;
  assign n26105 = n823 | n2111 ;
  assign n26106 = n4249 | n26105 ;
  assign n26107 = n162 | n360 ;
  assign n26108 = n542 | n26107 ;
  assign n26109 = n152 | n26108 ;
  assign n26110 = n26106 | n26109 ;
  assign n26111 = n26104 | n26110 ;
  assign n26112 = n607 | n26111 ;
  assign n26113 = n810 | n2601 ;
  assign n26114 = n5596 | n26113 ;
  assign n26115 = n3431 | n26114 ;
  assign n26116 = n26112 | n26115 ;
  assign n26117 = n1521 | n12746 ;
  assign n26118 = n26116 | n26117 ;
  assign n26119 = n26102 | n26118 ;
  assign n26120 = n26102 & n26118 ;
  assign n36003 = ~n26120 ;
  assign n26121 = n26119 & n36003 ;
  assign n20322 = n889 & n20311 ;
  assign n19910 = n3329 & n19893 ;
  assign n19924 = n3311 & n19917 ;
  assign n26122 = n19910 | n19924 ;
  assign n26123 = n3343 & n19870 ;
  assign n26124 = n26122 | n26123 ;
  assign n26125 = n20322 | n26124 ;
  assign n36004 = ~n26125 ;
  assign n26126 = n26121 & n36004 ;
  assign n36005 = ~n26121 ;
  assign n26127 = n36005 & n26125 ;
  assign n26128 = n26126 | n26127 ;
  assign n20554 = n895 & n34450 ;
  assign n19868 = n2861 & n19846 ;
  assign n20089 = n2849 & n20067 ;
  assign n26129 = n19868 | n20089 ;
  assign n26130 = n894 & n34452 ;
  assign n26131 = n26129 | n26130 ;
  assign n26132 = n20554 | n26131 ;
  assign n26133 = x29 | n26132 ;
  assign n26134 = x29 & n26132 ;
  assign n36006 = ~n26134 ;
  assign n26135 = n26133 & n36006 ;
  assign n26136 = n26128 & n26135 ;
  assign n26137 = n26128 | n26135 ;
  assign n36007 = ~n26136 ;
  assign n26138 = n36007 & n26137 ;
  assign n26139 = n25897 | n25901 ;
  assign n36008 = ~n26139 ;
  assign n26140 = n26138 & n36008 ;
  assign n36009 = ~n26138 ;
  assign n26141 = n36009 & n26139 ;
  assign n26142 = n26140 | n26141 ;
  assign n20872 = n3791 & n20863 ;
  assign n19816 = n3802 & n34355 ;
  assign n19833 = n209 & n19824 ;
  assign n26143 = n19816 | n19833 ;
  assign n26144 = n3818 & n34536 ;
  assign n26145 = n26143 | n26144 ;
  assign n26146 = n20872 | n26145 ;
  assign n26147 = x26 | n26146 ;
  assign n26148 = x26 & n26146 ;
  assign n36010 = ~n26148 ;
  assign n26149 = n26147 & n36010 ;
  assign n36011 = ~n26142 ;
  assign n26150 = n36011 & n26149 ;
  assign n36012 = ~n26149 ;
  assign n26151 = n26142 & n36012 ;
  assign n26152 = n26150 | n26151 ;
  assign n36013 = ~n25913 ;
  assign n26153 = n36013 & n25915 ;
  assign n26154 = n25911 | n26153 ;
  assign n36014 = ~n26154 ;
  assign n26155 = n26152 & n36014 ;
  assign n36015 = ~n26152 ;
  assign n26156 = n36015 & n26154 ;
  assign n26157 = n26155 | n26156 ;
  assign n21103 = n4135 & n34603 ;
  assign n19739 = n4148 & n34520 ;
  assign n19759 = n4185 & n19752 ;
  assign n26158 = n19739 | n19759 ;
  assign n26159 = n4165 & n34596 ;
  assign n26160 = n26158 | n26159 ;
  assign n26161 = n21103 | n26160 ;
  assign n26162 = x23 | n26161 ;
  assign n26163 = x23 & n26161 ;
  assign n36016 = ~n26163 ;
  assign n26164 = n26162 & n36016 ;
  assign n36017 = ~n26157 ;
  assign n26165 = n36017 & n26164 ;
  assign n36018 = ~n26164 ;
  assign n26166 = n26157 & n36018 ;
  assign n26167 = n26165 | n26166 ;
  assign n26168 = n25861 | n25928 ;
  assign n36019 = ~n25927 ;
  assign n26169 = n36019 & n26168 ;
  assign n26170 = n26167 & n26169 ;
  assign n26171 = n26167 | n26169 ;
  assign n36020 = ~n26170 ;
  assign n26172 = n36020 & n26171 ;
  assign n21878 = n4686 & n34817 ;
  assign n19674 = n4706 & n34360 ;
  assign n19688 = n4726 & n34349 ;
  assign n26173 = n19674 | n19688 ;
  assign n26174 = n4748 & n34803 ;
  assign n26175 = n26173 | n26174 ;
  assign n26176 = n21878 | n26175 ;
  assign n26177 = x20 | n26176 ;
  assign n26178 = x20 & n26176 ;
  assign n36021 = ~n26178 ;
  assign n26179 = n26177 & n36021 ;
  assign n36022 = ~n26172 ;
  assign n26180 = n36022 & n26179 ;
  assign n36023 = ~n26179 ;
  assign n26181 = n26172 & n36023 ;
  assign n26182 = n26180 | n26181 ;
  assign n36024 = ~n25938 ;
  assign n26183 = n25931 & n36024 ;
  assign n36025 = ~n26183 ;
  assign n26184 = n25944 & n36025 ;
  assign n26185 = n26182 & n26184 ;
  assign n26186 = n26182 | n26184 ;
  assign n36026 = ~n26185 ;
  assign n26187 = n36026 & n26186 ;
  assign n22650 = n37300 & n35035 ;
  assign n21742 = n5144 & n21729 ;
  assign n21814 = n5166 & n21753 ;
  assign n26188 = n21742 | n21814 ;
  assign n26189 = n5191 & n35018 ;
  assign n26190 = n26188 | n26189 ;
  assign n26191 = n22650 | n26190 ;
  assign n26192 = x17 | n26191 ;
  assign n26193 = x17 & n26191 ;
  assign n36027 = ~n26193 ;
  assign n26194 = n26192 & n36027 ;
  assign n36028 = ~n26187 ;
  assign n26195 = n36028 & n26194 ;
  assign n36029 = ~n26194 ;
  assign n26196 = n26187 & n36029 ;
  assign n26197 = n26195 | n26196 ;
  assign n26198 = n25954 | n25958 ;
  assign n36030 = ~n25955 ;
  assign n26199 = n36030 & n26198 ;
  assign n36031 = ~n26199 ;
  assign n26200 = n26197 & n36031 ;
  assign n36032 = ~n26197 ;
  assign n26201 = n36032 & n26199 ;
  assign n26202 = n26200 | n26201 ;
  assign n36033 = ~n26202 ;
  assign n26203 = n26099 & n36033 ;
  assign n36034 = ~n26099 ;
  assign n26204 = n36034 & n26202 ;
  assign n26205 = n26203 | n26204 ;
  assign n26206 = n25964 | n25965 ;
  assign n36035 = ~n25963 ;
  assign n26207 = n36035 & n26206 ;
  assign n36036 = ~n26207 ;
  assign n26208 = n26205 & n36036 ;
  assign n36037 = ~n26205 ;
  assign n26209 = n36037 & n26207 ;
  assign n26210 = n26208 | n26209 ;
  assign n24197 = n6272 & n35472 ;
  assign n23300 = n6190 & n35467 ;
  assign n23319 = n6244 & n35244 ;
  assign n26211 = n23300 | n23319 ;
  assign n26212 = n6217 & n35465 ;
  assign n26213 = n26211 | n26212 ;
  assign n26214 = n24197 | n26213 ;
  assign n26215 = x11 | n26214 ;
  assign n26216 = x11 & n26214 ;
  assign n36038 = ~n26216 ;
  assign n26217 = n26215 & n36038 ;
  assign n36039 = ~n26210 ;
  assign n26218 = n36039 & n26217 ;
  assign n36040 = ~n26217 ;
  assign n26219 = n26210 & n36040 ;
  assign n26220 = n26218 | n26219 ;
  assign n26221 = n25978 | n25980 ;
  assign n36041 = ~n25977 ;
  assign n26222 = n36041 & n26221 ;
  assign n36042 = ~n26222 ;
  assign n26223 = n26220 & n36042 ;
  assign n36043 = ~n26220 ;
  assign n26224 = n36043 & n26222 ;
  assign n26225 = n26223 | n26224 ;
  assign n25291 = n7068 & n25288 ;
  assign n24065 = n69 & n24057 ;
  assign n24084 = n7041 & n24080 ;
  assign n26226 = n24065 | n24084 ;
  assign n26227 = n7017 & n24676 ;
  assign n26228 = n26226 | n26227 ;
  assign n26229 = n25291 | n26228 ;
  assign n26230 = x8 | n26229 ;
  assign n26231 = x8 & n26229 ;
  assign n36044 = ~n26231 ;
  assign n26232 = n26230 & n36044 ;
  assign n26233 = n26225 & n26232 ;
  assign n26234 = n26225 | n26232 ;
  assign n36045 = ~n26233 ;
  assign n26235 = n36045 & n26234 ;
  assign n26236 = n25993 | n25994 ;
  assign n36046 = ~n25992 ;
  assign n26237 = n36046 & n26236 ;
  assign n36047 = ~n26237 ;
  assign n26238 = n26235 & n36047 ;
  assign n36048 = ~n26235 ;
  assign n26239 = n36048 & n26237 ;
  assign n26240 = n26238 | n26239 ;
  assign n25423 = n8157 & n35785 ;
  assign n24825 = n740 & n24815 ;
  assign n24849 = n8195 & n35663 ;
  assign n26241 = n24825 | n24849 ;
  assign n26242 = n9052 & n35784 ;
  assign n26243 = n26241 | n26242 ;
  assign n26244 = n25423 | n26243 ;
  assign n36049 = ~n26244 ;
  assign n26245 = x5 & n36049 ;
  assign n26246 = n30053 & n26244 ;
  assign n26247 = n26245 | n26246 ;
  assign n26248 = n26005 | n26009 ;
  assign n26249 = n26247 | n26248 ;
  assign n26250 = n26247 & n26248 ;
  assign n36050 = ~n26250 ;
  assign n26251 = n26249 & n36050 ;
  assign n26252 = n26240 & n26251 ;
  assign n26253 = n26240 | n26251 ;
  assign n36051 = ~n26252 ;
  assign n26254 = n36051 & n26253 ;
  assign n25808 = n9552 & n25796 ;
  assign n36052 = ~n5899 ;
  assign n26255 = n36052 & n25764 ;
  assign n26256 = n26025 | n26027 ;
  assign n36053 = ~n26255 ;
  assign n26257 = n36053 & n26256 ;
  assign n26258 = n25778 | n26020 ;
  assign n36054 = ~n26030 ;
  assign n26259 = n26023 & n36054 ;
  assign n36055 = ~n26259 ;
  assign n26260 = n26258 & n36055 ;
  assign n26261 = n26257 & n26260 ;
  assign n26262 = n26257 | n26260 ;
  assign n36056 = ~n26261 ;
  assign n26263 = n36056 & n26262 ;
  assign n26264 = n26017 | n26033 ;
  assign n36057 = ~n26014 ;
  assign n26265 = n36057 & n26036 ;
  assign n36058 = ~n26265 ;
  assign n26266 = n26264 & n36058 ;
  assign n5900 = n5793 & n32864 ;
  assign n26267 = x31 | n5793 ;
  assign n36059 = ~n5900 ;
  assign n26268 = n36059 & n26267 ;
  assign n26269 = n25778 | n26268 ;
  assign n26270 = x31 & n26268 ;
  assign n26271 = n25778 & n26270 ;
  assign n36060 = ~n26271 ;
  assign n26272 = n26269 & n36060 ;
  assign n26273 = n26266 | n26272 ;
  assign n26274 = n26266 & n26272 ;
  assign n36061 = ~n26274 ;
  assign n26275 = n26273 & n36061 ;
  assign n36062 = ~n26263 ;
  assign n26276 = n36062 & n26275 ;
  assign n36063 = ~n26275 ;
  assign n26277 = n26263 & n36063 ;
  assign n26278 = n26276 | n26277 ;
  assign n36064 = ~n26059 ;
  assign n26060 = n26039 & n36064 ;
  assign n36065 = ~n26039 ;
  assign n26280 = n36065 & n26061 ;
  assign n26281 = n26060 | n26280 ;
  assign n36066 = ~n26278 ;
  assign n26282 = n36066 & n26281 ;
  assign n36067 = ~n26281 ;
  assign n26283 = n26278 & n36067 ;
  assign n26284 = n26282 | n26283 ;
  assign n26285 = n9562 & n26284 ;
  assign n26295 = n10126 & n26039 ;
  assign n26296 = n10105 & n26278 ;
  assign n26297 = n26295 | n26296 ;
  assign n26298 = n26285 | n26297 ;
  assign n36068 = ~n26298 ;
  assign n26299 = x2 & n36068 ;
  assign n26300 = n30049 & n26298 ;
  assign n26301 = n26299 | n26300 ;
  assign n36069 = ~n25808 ;
  assign n26302 = n36069 & n26301 ;
  assign n36070 = ~n26254 ;
  assign n26303 = n36070 & n26302 ;
  assign n36071 = ~n26302 ;
  assign n26304 = n26254 & n36071 ;
  assign n26305 = n26303 | n26304 ;
  assign n26306 = n26012 | n26084 ;
  assign n26307 = n35999 & n26306 ;
  assign n36072 = ~n26305 ;
  assign n26308 = n36072 & n26307 ;
  assign n36073 = ~n26307 ;
  assign n26309 = n26305 & n36073 ;
  assign n26310 = n26308 | n26309 ;
  assign n36074 = ~n26310 ;
  assign n26311 = n26092 & n36074 ;
  assign n36075 = ~n26092 ;
  assign n26312 = n36075 & n26310 ;
  assign n29909 = n26311 | n26312 ;
  assign n26313 = n26250 | n26252 ;
  assign n26314 = n26172 | n26179 ;
  assign n36076 = ~n26184 ;
  assign n26315 = n26182 & n36076 ;
  assign n36077 = ~n26315 ;
  assign n26316 = n26314 & n36077 ;
  assign n26317 = n26157 | n26164 ;
  assign n36078 = ~n26169 ;
  assign n26318 = n26167 & n36078 ;
  assign n36079 = ~n26318 ;
  assign n26319 = n26317 & n36079 ;
  assign n36080 = ~n26140 ;
  assign n26320 = n26137 & n36080 ;
  assign n26321 = n26121 & n26125 ;
  assign n26322 = n26120 | n26321 ;
  assign n26323 = n338 | n833 ;
  assign n26324 = n2204 | n26323 ;
  assign n26325 = n623 | n916 ;
  assign n26326 = n26324 | n26325 ;
  assign n26327 = n521 | n1825 ;
  assign n26328 = n3031 | n26327 ;
  assign n26329 = n11239 | n26328 ;
  assign n26330 = n26326 | n26329 ;
  assign n26331 = n1620 | n1653 ;
  assign n26332 = n2305 | n26331 ;
  assign n26333 = n13213 | n26332 ;
  assign n26334 = n26330 | n26333 ;
  assign n26335 = n2120 | n26334 ;
  assign n36081 = ~n5546 ;
  assign n26336 = n36081 & n5603 ;
  assign n36082 = ~n26335 ;
  assign n26337 = n36082 & n26336 ;
  assign n26338 = n26322 & n26337 ;
  assign n26339 = n26322 | n26337 ;
  assign n36083 = ~n26338 ;
  assign n26340 = n36083 & n26339 ;
  assign n20497 = n889 & n20486 ;
  assign n19890 = n3329 & n19870 ;
  assign n19912 = n3311 & n19893 ;
  assign n26341 = n19890 | n19912 ;
  assign n26342 = n3343 & n19846 ;
  assign n26343 = n26341 | n26342 ;
  assign n26344 = n20497 | n26343 ;
  assign n26345 = n26340 | n26344 ;
  assign n26346 = n26340 & n26344 ;
  assign n36084 = ~n26346 ;
  assign n26347 = n26345 & n36084 ;
  assign n20517 = n895 & n34442 ;
  assign n20080 = n2861 & n20067 ;
  assign n20101 = n2849 & n34354 ;
  assign n26348 = n20080 | n20101 ;
  assign n26349 = n894 & n20527 ;
  assign n26350 = n26348 | n26349 ;
  assign n26351 = n20517 | n26350 ;
  assign n26352 = x29 | n26351 ;
  assign n26353 = x29 & n26351 ;
  assign n36085 = ~n26353 ;
  assign n26354 = n26352 & n36085 ;
  assign n36086 = ~n26347 ;
  assign n26355 = n36086 & n26354 ;
  assign n36087 = ~n26354 ;
  assign n26356 = n26347 & n36087 ;
  assign n26357 = n26355 | n26356 ;
  assign n36088 = ~n26357 ;
  assign n26358 = n26320 & n36088 ;
  assign n36089 = ~n26320 ;
  assign n26359 = n36089 & n26357 ;
  assign n26360 = n26358 | n26359 ;
  assign n20838 = n3791 & n20833 ;
  assign n19794 = n3802 & n34519 ;
  assign n19819 = n209 & n34355 ;
  assign n26361 = n19794 | n19819 ;
  assign n26362 = n3818 & n20845 ;
  assign n26363 = n26361 | n26362 ;
  assign n26364 = n20838 | n26363 ;
  assign n26365 = x26 | n26364 ;
  assign n26366 = x26 & n26364 ;
  assign n36090 = ~n26366 ;
  assign n26367 = n26365 & n36090 ;
  assign n36091 = ~n26360 ;
  assign n26368 = n36091 & n26367 ;
  assign n36092 = ~n26367 ;
  assign n26369 = n26360 & n36092 ;
  assign n26370 = n26368 | n26369 ;
  assign n26371 = n26142 | n26149 ;
  assign n36093 = ~n26155 ;
  assign n26372 = n36093 & n26371 ;
  assign n36094 = ~n26370 ;
  assign n26373 = n36094 & n26372 ;
  assign n36095 = ~n26372 ;
  assign n26374 = n26370 & n36095 ;
  assign n26375 = n26373 | n26374 ;
  assign n21079 = n4135 & n34598 ;
  assign n19716 = n4148 & n34363 ;
  assign n19743 = n4185 & n34520 ;
  assign n26376 = n19716 | n19743 ;
  assign n26377 = n4165 & n34349 ;
  assign n26378 = n26376 | n26377 ;
  assign n26379 = n21079 | n26378 ;
  assign n26380 = x23 | n26379 ;
  assign n26381 = x23 & n26379 ;
  assign n36096 = ~n26381 ;
  assign n26382 = n26380 & n36096 ;
  assign n36097 = ~n26375 ;
  assign n26383 = n36097 & n26382 ;
  assign n36098 = ~n26382 ;
  assign n26384 = n26375 & n36098 ;
  assign n26385 = n26383 | n26384 ;
  assign n36099 = ~n26385 ;
  assign n26386 = n26319 & n36099 ;
  assign n36100 = ~n26319 ;
  assign n26387 = n36100 & n26385 ;
  assign n26388 = n26386 | n26387 ;
  assign n21856 = n4686 & n21848 ;
  assign n19675 = n4726 & n34360 ;
  assign n21770 = n4706 & n34803 ;
  assign n26389 = n19675 | n21770 ;
  assign n26390 = n4748 & n21753 ;
  assign n26391 = n26389 | n26390 ;
  assign n26392 = n21856 | n26391 ;
  assign n26393 = x20 | n26392 ;
  assign n26394 = x20 & n26392 ;
  assign n36101 = ~n26394 ;
  assign n26395 = n26393 & n36101 ;
  assign n36102 = ~n26388 ;
  assign n26396 = n36102 & n26395 ;
  assign n36103 = ~n26395 ;
  assign n26397 = n26388 & n36103 ;
  assign n26398 = n26396 | n26397 ;
  assign n26399 = n26316 | n26398 ;
  assign n26400 = n26316 & n26398 ;
  assign n36104 = ~n26400 ;
  assign n26401 = n26399 & n36104 ;
  assign n22627 = n37300 & n35030 ;
  assign n21744 = n5166 & n21729 ;
  assign n22536 = n5144 & n35018 ;
  assign n26402 = n21744 | n22536 ;
  assign n26403 = n5191 & n22533 ;
  assign n26404 = n26402 | n26403 ;
  assign n26405 = n22627 | n26404 ;
  assign n26406 = x17 | n26405 ;
  assign n26407 = x17 & n26405 ;
  assign n36105 = ~n26407 ;
  assign n26408 = n26406 & n36105 ;
  assign n36106 = ~n26401 ;
  assign n26409 = n36106 & n26408 ;
  assign n36107 = ~n26408 ;
  assign n26410 = n26401 & n36107 ;
  assign n26411 = n26409 | n26410 ;
  assign n26412 = n26187 | n26194 ;
  assign n36108 = ~n26200 ;
  assign n26413 = n36108 & n26412 ;
  assign n36109 = ~n26411 ;
  assign n26414 = n36109 & n26413 ;
  assign n36110 = ~n26413 ;
  assign n26415 = n26411 & n36110 ;
  assign n26416 = n26414 | n26415 ;
  assign n23409 = n5937 & n35252 ;
  assign n22511 = n5994 & n35020 ;
  assign n23342 = n5970 & n23339 ;
  assign n26417 = n22511 | n23342 ;
  assign n26418 = n6018 & n35254 ;
  assign n26419 = n26417 | n26418 ;
  assign n26420 = n23409 | n26419 ;
  assign n26421 = x14 | n26420 ;
  assign n26422 = x14 & n26420 ;
  assign n36111 = ~n26422 ;
  assign n26423 = n26421 & n36111 ;
  assign n26424 = n26416 & n26423 ;
  assign n26425 = n26416 | n26423 ;
  assign n36112 = ~n26424 ;
  assign n26426 = n36112 & n26425 ;
  assign n26427 = n26099 | n26202 ;
  assign n36113 = ~n26208 ;
  assign n26428 = n36113 & n26427 ;
  assign n26429 = n26426 & n26428 ;
  assign n26430 = n26426 | n26428 ;
  assign n36114 = ~n26429 ;
  assign n26431 = n36114 & n26430 ;
  assign n24172 = n6272 & n24168 ;
  assign n23299 = n6244 & n35467 ;
  assign n24107 = n6190 & n35458 ;
  assign n26432 = n23299 | n24107 ;
  assign n26433 = n6217 & n24080 ;
  assign n26434 = n26432 | n26433 ;
  assign n26435 = n24172 | n26434 ;
  assign n26436 = x11 | n26435 ;
  assign n26437 = x11 & n26435 ;
  assign n36115 = ~n26437 ;
  assign n26438 = n26436 & n36115 ;
  assign n26439 = n26431 & n26438 ;
  assign n26440 = n26431 | n26438 ;
  assign n36116 = ~n26439 ;
  assign n26441 = n36116 & n26440 ;
  assign n26442 = n26210 | n26217 ;
  assign n36117 = ~n26223 ;
  assign n26443 = n36117 & n26442 ;
  assign n36118 = ~n26441 ;
  assign n26444 = n36118 & n26443 ;
  assign n36119 = ~n26443 ;
  assign n26445 = n26441 & n36119 ;
  assign n26446 = n26444 | n26445 ;
  assign n25321 = n7068 & n35670 ;
  assign n24066 = n7041 & n24057 ;
  assign n24679 = n69 & n24676 ;
  assign n26447 = n24066 | n24679 ;
  assign n26448 = n7017 & n35663 ;
  assign n26449 = n26447 | n26448 ;
  assign n26450 = n25321 | n26449 ;
  assign n26451 = x8 | n26450 ;
  assign n26452 = x8 & n26450 ;
  assign n36120 = ~n26452 ;
  assign n26453 = n26451 & n36120 ;
  assign n36121 = ~n26446 ;
  assign n26454 = n36121 & n26453 ;
  assign n36122 = ~n26453 ;
  assign n26455 = n26446 & n36122 ;
  assign n26456 = n26454 | n26455 ;
  assign n36123 = ~n26238 ;
  assign n26457 = n26234 & n36123 ;
  assign n26458 = n26456 & n26457 ;
  assign n26459 = n26456 | n26457 ;
  assign n36124 = ~n26458 ;
  assign n26460 = n36124 & n26459 ;
  assign n25827 = n8157 & n35910 ;
  assign n24823 = n8195 & n24815 ;
  assign n25406 = n740 & n35784 ;
  assign n26461 = n24823 | n25406 ;
  assign n26462 = n9052 & n25796 ;
  assign n26463 = n26461 | n26462 ;
  assign n26464 = n25827 | n26463 ;
  assign n26465 = x5 | n26464 ;
  assign n26466 = x5 & n26464 ;
  assign n36125 = ~n26466 ;
  assign n26467 = n26465 & n36125 ;
  assign n36126 = ~n26460 ;
  assign n26468 = n36126 & n26467 ;
  assign n36127 = ~n26467 ;
  assign n26469 = n26460 & n36127 ;
  assign n26470 = n26468 | n26469 ;
  assign n26471 = n26313 | n26470 ;
  assign n26472 = n26313 & n26470 ;
  assign n36128 = ~n26472 ;
  assign n26473 = n26471 & n36128 ;
  assign n26048 = n9552 & n26039 ;
  assign n26484 = n26039 | n26061 ;
  assign n26485 = n26059 & n36066 ;
  assign n36129 = ~n26485 ;
  assign n26486 = n26484 & n36129 ;
  assign n36130 = ~n26486 ;
  assign n26487 = n9562 & n36130 ;
  assign n26500 = n10126 & n26278 ;
  assign n26279 = n26039 | n26278 ;
  assign n36131 = ~n26279 ;
  assign n26501 = n10105 & n36131 ;
  assign n26502 = n26500 | n26501 ;
  assign n26503 = n26487 | n26502 ;
  assign n36132 = ~n26503 ;
  assign n26504 = x2 & n36132 ;
  assign n26505 = n30049 & n26503 ;
  assign n26506 = n26504 | n26505 ;
  assign n36133 = ~n26048 ;
  assign n26507 = n36133 & n26506 ;
  assign n26508 = n26473 & n26507 ;
  assign n26509 = n26473 | n26507 ;
  assign n36134 = ~n26508 ;
  assign n26510 = n36134 & n26509 ;
  assign n26511 = n26254 | n26302 ;
  assign n36135 = ~n26309 ;
  assign n26512 = n36135 & n26511 ;
  assign n26513 = n26510 | n26512 ;
  assign n26514 = n26510 & n26512 ;
  assign n36136 = ~n26514 ;
  assign n26515 = n26513 & n36136 ;
  assign n36137 = ~n26312 ;
  assign n26516 = n36137 & n26515 ;
  assign n36138 = ~n26515 ;
  assign n26517 = n26312 & n36138 ;
  assign n29908 = n26516 | n26517 ;
  assign n26067 = n8157 & n26065 ;
  assign n25396 = n8195 & n35784 ;
  assign n25801 = n740 & n25796 ;
  assign n26518 = n25396 | n25801 ;
  assign n26519 = n9052 & n26039 ;
  assign n26520 = n26518 | n26519 ;
  assign n26521 = n26067 | n26520 ;
  assign n26522 = x5 | n26521 ;
  assign n26523 = x5 & n26521 ;
  assign n36139 = ~n26523 ;
  assign n26524 = n26522 & n36139 ;
  assign n36140 = ~n26469 ;
  assign n26525 = n36140 & n26471 ;
  assign n26526 = n26524 & n26525 ;
  assign n26527 = n26524 | n26525 ;
  assign n36141 = ~n26526 ;
  assign n26528 = n36141 & n26527 ;
  assign n23377 = n5937 & n23372 ;
  assign n23320 = n5970 & n35244 ;
  assign n23343 = n5994 & n23339 ;
  assign n26529 = n23320 | n23343 ;
  assign n26530 = n6018 & n35246 ;
  assign n26531 = n26529 | n26530 ;
  assign n26532 = n23377 | n26531 ;
  assign n36142 = ~n26532 ;
  assign n26533 = x14 & n36142 ;
  assign n26534 = n30547 & n26532 ;
  assign n26535 = n26533 | n26534 ;
  assign n26536 = n1324 | n3750 ;
  assign n26537 = n4591 | n26536 ;
  assign n26538 = n245 | n534 ;
  assign n26539 = n684 | n695 ;
  assign n26540 = n26538 | n26539 ;
  assign n26541 = n723 | n26540 ;
  assign n26542 = n26537 | n26541 ;
  assign n26543 = n25872 | n26542 ;
  assign n26544 = n3729 | n4997 ;
  assign n26545 = n225 | n381 ;
  assign n26546 = n2029 | n26545 ;
  assign n36143 = ~n26546 ;
  assign n26547 = n147 & n36143 ;
  assign n36144 = ~n26544 ;
  assign n26548 = n36144 & n26547 ;
  assign n26549 = n1609 | n2154 ;
  assign n26550 = n4039 | n26549 ;
  assign n26551 = n214 | n811 ;
  assign n26552 = n845 | n26551 ;
  assign n26553 = n966 | n26552 ;
  assign n26554 = n1191 | n1583 ;
  assign n26555 = n26553 | n26554 ;
  assign n26556 = n26550 | n26555 ;
  assign n36145 = ~n26556 ;
  assign n26557 = n26548 & n36145 ;
  assign n36146 = ~n26543 ;
  assign n26558 = n36146 & n26557 ;
  assign n36147 = ~n12289 ;
  assign n26559 = n36147 & n26558 ;
  assign n26560 = n32141 & n26559 ;
  assign n20585 = n889 & n20579 ;
  assign n19856 = n3329 & n19846 ;
  assign n19891 = n3311 & n19870 ;
  assign n26561 = n19856 | n19891 ;
  assign n26562 = n3343 & n20067 ;
  assign n26563 = n26561 | n26562 ;
  assign n26564 = n20585 | n26563 ;
  assign n36148 = ~n26564 ;
  assign n26565 = n26560 & n36148 ;
  assign n36149 = ~n26560 ;
  assign n26566 = n36149 & n26564 ;
  assign n26567 = n26565 | n26566 ;
  assign n36150 = ~n26337 ;
  assign n26568 = n26322 & n36150 ;
  assign n36151 = ~n26340 ;
  assign n26569 = n36151 & n26344 ;
  assign n26570 = n26568 | n26569 ;
  assign n26571 = n26567 | n26570 ;
  assign n26572 = n26567 & n26570 ;
  assign n36152 = ~n26572 ;
  assign n26573 = n26571 & n36152 ;
  assign n20780 = n895 & n34511 ;
  assign n19843 = n2849 & n19824 ;
  assign n20113 = n2861 & n34354 ;
  assign n26574 = n19843 | n20113 ;
  assign n26575 = n894 & n34513 ;
  assign n26576 = n26574 | n26575 ;
  assign n26577 = n20780 | n26576 ;
  assign n26578 = x29 | n26577 ;
  assign n26579 = x29 & n26577 ;
  assign n36153 = ~n26579 ;
  assign n26580 = n26578 & n36153 ;
  assign n26581 = n26573 & n26580 ;
  assign n26582 = n26573 | n26580 ;
  assign n36154 = ~n26581 ;
  assign n26583 = n36154 & n26582 ;
  assign n26584 = n26355 | n26358 ;
  assign n26585 = n26583 | n26584 ;
  assign n26586 = n26583 & n26584 ;
  assign n36155 = ~n26586 ;
  assign n26587 = n26585 & n36155 ;
  assign n20811 = n3791 & n20805 ;
  assign n19769 = n3802 & n19752 ;
  assign n19786 = n209 & n34519 ;
  assign n26588 = n19769 | n19786 ;
  assign n26589 = n3818 & n34520 ;
  assign n26590 = n26588 | n26589 ;
  assign n26591 = n20811 | n26590 ;
  assign n26592 = x26 | n26591 ;
  assign n26593 = x26 & n26591 ;
  assign n36156 = ~n26593 ;
  assign n26594 = n26592 & n36156 ;
  assign n26595 = n26587 & n26594 ;
  assign n26596 = n26587 | n26594 ;
  assign n36157 = ~n26595 ;
  assign n26597 = n36157 & n26596 ;
  assign n26598 = n26368 | n26373 ;
  assign n26599 = n26597 | n26598 ;
  assign n26600 = n26597 & n26598 ;
  assign n36158 = ~n26600 ;
  assign n26601 = n26599 & n36158 ;
  assign n20155 = n4135 & n34362 ;
  assign n19698 = n4148 & n34349 ;
  assign n19725 = n4185 & n34363 ;
  assign n26602 = n19698 | n19725 ;
  assign n26603 = n4165 & n34365 ;
  assign n26604 = n26602 | n26603 ;
  assign n26605 = n20155 | n26604 ;
  assign n26606 = x23 | n26605 ;
  assign n26607 = x23 & n26605 ;
  assign n36159 = ~n26607 ;
  assign n26608 = n26606 & n36159 ;
  assign n26609 = n26601 & n26608 ;
  assign n26610 = n26601 | n26608 ;
  assign n36160 = ~n26609 ;
  assign n26611 = n36160 & n26610 ;
  assign n26612 = n26383 | n26386 ;
  assign n26613 = n26611 | n26612 ;
  assign n26614 = n26611 & n26612 ;
  assign n36161 = ~n26614 ;
  assign n26615 = n26613 & n36161 ;
  assign n21798 = n4686 & n34802 ;
  assign n21769 = n4726 & n34803 ;
  assign n21820 = n4706 & n21753 ;
  assign n26616 = n21769 | n21820 ;
  assign n26617 = n4748 & n21804 ;
  assign n26618 = n26616 | n26617 ;
  assign n26619 = n21798 | n26618 ;
  assign n26620 = x20 | n26619 ;
  assign n26621 = x20 & n26619 ;
  assign n36162 = ~n26621 ;
  assign n26622 = n26620 & n36162 ;
  assign n26623 = n26615 & n26622 ;
  assign n26624 = n26615 | n26622 ;
  assign n36163 = ~n26623 ;
  assign n26625 = n36163 & n26624 ;
  assign n36164 = ~n26398 ;
  assign n26626 = n26316 & n36164 ;
  assign n26627 = n26396 | n26626 ;
  assign n26628 = n26625 | n26627 ;
  assign n26629 = n26625 & n26627 ;
  assign n36165 = ~n26629 ;
  assign n26630 = n26628 & n36165 ;
  assign n22570 = n37300 & n35022 ;
  assign n22541 = n5166 & n35018 ;
  assign n22583 = n5144 & n22533 ;
  assign n26631 = n22541 | n22583 ;
  assign n26632 = n5191 & n35020 ;
  assign n26633 = n26631 | n26632 ;
  assign n26634 = n22570 | n26633 ;
  assign n26635 = x17 | n26634 ;
  assign n26636 = x17 & n26634 ;
  assign n36166 = ~n26636 ;
  assign n26637 = n26635 & n36166 ;
  assign n36167 = ~n26630 ;
  assign n26638 = n36167 & n26637 ;
  assign n36168 = ~n26637 ;
  assign n26639 = n26630 & n36168 ;
  assign n26640 = n26638 | n26639 ;
  assign n26641 = n26411 | n26413 ;
  assign n36169 = ~n26410 ;
  assign n26642 = n36169 & n26641 ;
  assign n26643 = n26640 & n26642 ;
  assign n26644 = n26640 | n26642 ;
  assign n36170 = ~n26643 ;
  assign n26645 = n36170 & n26644 ;
  assign n36171 = ~n26535 ;
  assign n26646 = n36171 & n26645 ;
  assign n36172 = ~n26645 ;
  assign n26647 = n26535 & n36172 ;
  assign n26648 = n26646 | n26647 ;
  assign n36173 = ~n26423 ;
  assign n26649 = n26416 & n36173 ;
  assign n36174 = ~n26649 ;
  assign n26650 = n26430 & n36174 ;
  assign n26651 = n26648 | n26650 ;
  assign n26652 = n26648 & n26650 ;
  assign n36175 = ~n26652 ;
  assign n26653 = n26651 & n36175 ;
  assign n24143 = n6272 & n35457 ;
  assign n24083 = n6190 & n24080 ;
  assign n24105 = n6244 & n35458 ;
  assign n26654 = n24083 | n24105 ;
  assign n26655 = n6217 & n24151 ;
  assign n26656 = n26654 | n26655 ;
  assign n26657 = n24143 | n26656 ;
  assign n26658 = x11 | n26657 ;
  assign n26659 = x11 & n26657 ;
  assign n36176 = ~n26659 ;
  assign n26660 = n26658 & n36176 ;
  assign n26661 = n26653 & n26660 ;
  assign n26662 = n26653 | n26660 ;
  assign n36177 = ~n26661 ;
  assign n26663 = n36177 & n26662 ;
  assign n36178 = ~n26438 ;
  assign n26664 = n26431 & n36178 ;
  assign n26665 = n26441 | n26443 ;
  assign n36179 = ~n26664 ;
  assign n26666 = n36179 & n26665 ;
  assign n36180 = ~n26663 ;
  assign n26667 = n36180 & n26666 ;
  assign n36181 = ~n26666 ;
  assign n26668 = n26663 & n36181 ;
  assign n26669 = n26667 | n26668 ;
  assign n24879 = n7068 & n35662 ;
  assign n24688 = n7041 & n24676 ;
  assign n24848 = n69 & n35663 ;
  assign n26670 = n24688 | n24848 ;
  assign n26671 = n7017 & n24815 ;
  assign n26672 = n26670 | n26671 ;
  assign n26673 = n24879 | n26672 ;
  assign n26674 = x8 | n26673 ;
  assign n26675 = x8 & n26673 ;
  assign n36182 = ~n26675 ;
  assign n26676 = n26674 & n36182 ;
  assign n26677 = n26669 & n26676 ;
  assign n26678 = n26669 | n26676 ;
  assign n36183 = ~n26677 ;
  assign n26679 = n36183 & n26678 ;
  assign n36184 = ~n26456 ;
  assign n26680 = n36184 & n26457 ;
  assign n26681 = n26454 | n26680 ;
  assign n36185 = ~n26679 ;
  assign n26682 = n36185 & n26681 ;
  assign n36186 = ~n26681 ;
  assign n26683 = n26679 & n36186 ;
  assign n26684 = n26682 | n26683 ;
  assign n26685 = n26528 | n26684 ;
  assign n26686 = n26528 & n26684 ;
  assign n36187 = ~n26686 ;
  assign n26687 = n26685 & n36187 ;
  assign n36188 = ~n26507 ;
  assign n26688 = n26473 & n36188 ;
  assign n36189 = ~n26688 ;
  assign n26689 = n26513 & n36189 ;
  assign n26690 = n26687 & n26689 ;
  assign n26691 = n26687 | n26689 ;
  assign n36190 = ~n26690 ;
  assign n26692 = n36190 & n26691 ;
  assign n26693 = n9552 & n26278 ;
  assign n26497 = n10126 & n36131 ;
  assign n26694 = n26278 & n26484 ;
  assign n36191 = ~n26694 ;
  assign n26695 = n26279 & n36191 ;
  assign n36192 = ~n26695 ;
  assign n26696 = n9562 & n36192 ;
  assign n26706 = n26497 | n26696 ;
  assign n36193 = ~n26706 ;
  assign n26707 = x2 & n36193 ;
  assign n26708 = n30049 & n26706 ;
  assign n26709 = n26707 | n26708 ;
  assign n36194 = ~n26693 ;
  assign n26710 = n36194 & n26709 ;
  assign n26711 = n26692 & n26710 ;
  assign n26712 = n26692 | n26710 ;
  assign n36195 = ~n26711 ;
  assign n26713 = n36195 & n26712 ;
  assign n26714 = n26517 & n26713 ;
  assign n29906 = n26517 | n26713 ;
  assign n36196 = ~n26714 ;
  assign n29907 = n36196 & n29906 ;
  assign n36197 = ~n26713 ;
  assign n26715 = n26517 & n36197 ;
  assign n26716 = n26527 & n36187 ;
  assign n36198 = ~n26580 ;
  assign n26717 = n26573 & n36198 ;
  assign n36199 = ~n26717 ;
  assign n26718 = n26585 & n36199 ;
  assign n26719 = n406 | n747 ;
  assign n26720 = n4056 | n5482 ;
  assign n26721 = n26719 | n26720 ;
  assign n26722 = n181 | n203 ;
  assign n26723 = n446 | n630 ;
  assign n26724 = n26722 | n26723 ;
  assign n26725 = n4890 | n26724 ;
  assign n26726 = n5854 | n26725 ;
  assign n26727 = n26721 | n26726 ;
  assign n26728 = n4783 | n11568 ;
  assign n26729 = n13345 | n26728 ;
  assign n26730 = n26727 | n26729 ;
  assign n26731 = n3148 | n26730 ;
  assign n36200 = ~n26731 ;
  assign n26732 = n13734 & n36200 ;
  assign n20555 = n889 & n34450 ;
  assign n19865 = n3311 & n19846 ;
  assign n20077 = n3329 & n20067 ;
  assign n26733 = n19865 | n20077 ;
  assign n26734 = n3343 & n34452 ;
  assign n26735 = n26733 | n26734 ;
  assign n26736 = n20555 | n26735 ;
  assign n26737 = n26732 | n26736 ;
  assign n26738 = n26732 & n26736 ;
  assign n36201 = ~n26738 ;
  assign n26739 = n26737 & n36201 ;
  assign n36202 = ~n26565 ;
  assign n26740 = n36202 & n26571 ;
  assign n36203 = ~n26739 ;
  assign n26741 = n36203 & n26740 ;
  assign n36204 = ~n26740 ;
  assign n26742 = n26739 & n36204 ;
  assign n26743 = n26741 | n26742 ;
  assign n20874 = n895 & n20863 ;
  assign n19820 = n2849 & n34355 ;
  assign n19844 = n2861 & n19824 ;
  assign n26744 = n19820 | n19844 ;
  assign n26745 = n894 & n34536 ;
  assign n26746 = n26744 | n26745 ;
  assign n26747 = n20874 | n26746 ;
  assign n26748 = x29 | n26747 ;
  assign n26749 = x29 & n26747 ;
  assign n36205 = ~n26749 ;
  assign n26750 = n26748 & n36205 ;
  assign n36206 = ~n26743 ;
  assign n26751 = n36206 & n26750 ;
  assign n36207 = ~n26750 ;
  assign n26752 = n26743 & n36207 ;
  assign n26753 = n26751 | n26752 ;
  assign n36208 = ~n26753 ;
  assign n26754 = n26718 & n36208 ;
  assign n36209 = ~n26718 ;
  assign n26755 = n36209 & n26753 ;
  assign n26756 = n26754 | n26755 ;
  assign n21104 = n3791 & n34603 ;
  assign n19740 = n3802 & n34520 ;
  assign n19770 = n209 & n19752 ;
  assign n26757 = n19740 | n19770 ;
  assign n26758 = n3818 & n34596 ;
  assign n26759 = n26757 | n26758 ;
  assign n26760 = n21104 | n26759 ;
  assign n26761 = x26 | n26760 ;
  assign n26762 = x26 & n26760 ;
  assign n36210 = ~n26762 ;
  assign n26763 = n26761 & n36210 ;
  assign n36211 = ~n26756 ;
  assign n26764 = n36211 & n26763 ;
  assign n36212 = ~n26763 ;
  assign n26765 = n26756 & n36212 ;
  assign n26766 = n26764 | n26765 ;
  assign n36213 = ~n26594 ;
  assign n26767 = n26587 & n36213 ;
  assign n36214 = ~n26767 ;
  assign n26768 = n26599 & n36214 ;
  assign n36215 = ~n26766 ;
  assign n26769 = n36215 & n26768 ;
  assign n36216 = ~n26768 ;
  assign n26770 = n26766 & n36216 ;
  assign n26771 = n26769 | n26770 ;
  assign n21879 = n4135 & n34817 ;
  assign n19676 = n4148 & n34360 ;
  assign n19699 = n4185 & n34349 ;
  assign n26772 = n19676 | n19699 ;
  assign n26773 = n4165 & n34803 ;
  assign n26774 = n26772 | n26773 ;
  assign n26775 = n21879 | n26774 ;
  assign n26776 = x23 | n26775 ;
  assign n26777 = x23 & n26775 ;
  assign n36217 = ~n26777 ;
  assign n26778 = n26776 & n36217 ;
  assign n36218 = ~n26771 ;
  assign n26779 = n36218 & n26778 ;
  assign n36219 = ~n26778 ;
  assign n26780 = n26771 & n36219 ;
  assign n26781 = n26779 | n26780 ;
  assign n36220 = ~n26608 ;
  assign n26782 = n26601 & n36220 ;
  assign n36221 = ~n26782 ;
  assign n26783 = n26613 & n36221 ;
  assign n36222 = ~n26781 ;
  assign n26784 = n36222 & n26783 ;
  assign n36223 = ~n26783 ;
  assign n26785 = n26781 & n36223 ;
  assign n26786 = n26784 | n26785 ;
  assign n22651 = n4686 & n35035 ;
  assign n21745 = n4706 & n21729 ;
  assign n21821 = n4726 & n21753 ;
  assign n26787 = n21745 | n21821 ;
  assign n26788 = n4748 & n35018 ;
  assign n26789 = n26787 | n26788 ;
  assign n26790 = n22651 | n26789 ;
  assign n26791 = x20 | n26790 ;
  assign n26792 = x20 & n26790 ;
  assign n36224 = ~n26792 ;
  assign n26793 = n26791 & n36224 ;
  assign n36225 = ~n26786 ;
  assign n26794 = n36225 & n26793 ;
  assign n36226 = ~n26793 ;
  assign n26795 = n26786 & n36226 ;
  assign n26796 = n26794 | n26795 ;
  assign n36227 = ~n26622 ;
  assign n26797 = n26615 & n36227 ;
  assign n36228 = ~n26797 ;
  assign n26798 = n26628 & n36228 ;
  assign n36229 = ~n26796 ;
  assign n26799 = n36229 & n26798 ;
  assign n36230 = ~n26798 ;
  assign n26800 = n26796 & n36230 ;
  assign n26801 = n26799 | n26800 ;
  assign n23434 = n37300 & n35262 ;
  assign n22512 = n5144 & n35020 ;
  assign n22578 = n5166 & n22533 ;
  assign n26802 = n22512 | n22578 ;
  assign n26803 = n5191 & n23444 ;
  assign n26804 = n26802 | n26803 ;
  assign n26805 = n23434 | n26804 ;
  assign n26806 = x17 | n26805 ;
  assign n26807 = x17 & n26805 ;
  assign n36231 = ~n26807 ;
  assign n26808 = n26806 & n36231 ;
  assign n26809 = n26638 | n26642 ;
  assign n36232 = ~n26639 ;
  assign n26810 = n36232 & n26809 ;
  assign n36233 = ~n26810 ;
  assign n26811 = n26808 & n36233 ;
  assign n36234 = ~n26808 ;
  assign n26812 = n36234 & n26810 ;
  assign n26813 = n26811 | n26812 ;
  assign n36235 = ~n26801 ;
  assign n26814 = n36235 & n26813 ;
  assign n36236 = ~n26813 ;
  assign n26815 = n26801 & n36236 ;
  assign n26816 = n26814 | n26815 ;
  assign n24198 = n5937 & n35472 ;
  assign n23293 = n5970 & n35467 ;
  assign n23318 = n5994 & n35244 ;
  assign n26817 = n23293 | n23318 ;
  assign n26818 = n6018 & n35465 ;
  assign n26819 = n26817 | n26818 ;
  assign n26820 = n24198 | n26819 ;
  assign n26821 = x14 | n26820 ;
  assign n26822 = x14 & n26820 ;
  assign n36237 = ~n26822 ;
  assign n26823 = n26821 & n36237 ;
  assign n36238 = ~n26646 ;
  assign n26824 = n36238 & n26651 ;
  assign n26825 = n26823 & n26824 ;
  assign n26826 = n26823 | n26824 ;
  assign n36239 = ~n26825 ;
  assign n26827 = n36239 & n26826 ;
  assign n36240 = ~n26816 ;
  assign n26828 = n36240 & n26827 ;
  assign n36241 = ~n26827 ;
  assign n26829 = n26816 & n36241 ;
  assign n26830 = n26828 | n26829 ;
  assign n25293 = n6272 & n25288 ;
  assign n24069 = n6190 & n24057 ;
  assign n24090 = n6244 & n24080 ;
  assign n26831 = n24069 | n24090 ;
  assign n26832 = n6217 & n24676 ;
  assign n26833 = n26831 | n26832 ;
  assign n26834 = n25293 | n26833 ;
  assign n26835 = x11 | n26834 ;
  assign n26836 = x11 & n26834 ;
  assign n36242 = ~n26836 ;
  assign n26837 = n26835 & n36242 ;
  assign n36243 = ~n26830 ;
  assign n26838 = n36243 & n26837 ;
  assign n36244 = ~n26837 ;
  assign n26839 = n26830 & n36244 ;
  assign n26840 = n26838 | n26839 ;
  assign n36245 = ~n26653 ;
  assign n26841 = n36245 & n26660 ;
  assign n26842 = n26667 | n26841 ;
  assign n36246 = ~n26842 ;
  assign n26843 = n26840 & n36246 ;
  assign n36247 = ~n26840 ;
  assign n26844 = n36247 & n26842 ;
  assign n26845 = n26843 | n26844 ;
  assign n25424 = n7068 & n35785 ;
  assign n24822 = n69 & n24815 ;
  assign n24847 = n7041 & n35663 ;
  assign n26846 = n24822 | n24847 ;
  assign n26847 = n7017 & n35784 ;
  assign n26848 = n26846 | n26847 ;
  assign n26849 = n25424 | n26848 ;
  assign n26850 = x8 | n26849 ;
  assign n26851 = x8 & n26849 ;
  assign n36248 = ~n26851 ;
  assign n26852 = n26850 & n36248 ;
  assign n36249 = ~n26845 ;
  assign n26853 = n36249 & n26852 ;
  assign n36250 = ~n26852 ;
  assign n26854 = n26845 & n36250 ;
  assign n26855 = n26853 | n26854 ;
  assign n36251 = ~n26669 ;
  assign n26856 = n36251 & n26676 ;
  assign n26857 = n26682 | n26856 ;
  assign n36252 = ~n26857 ;
  assign n26858 = n26855 & n36252 ;
  assign n36253 = ~n26855 ;
  assign n26859 = n36253 & n26857 ;
  assign n26860 = n26858 | n26859 ;
  assign n26287 = n8157 & n26284 ;
  assign n25805 = n8195 & n25796 ;
  assign n26052 = n740 & n26039 ;
  assign n26861 = n25805 | n26052 ;
  assign n26862 = n9052 & n26278 ;
  assign n26863 = n26861 | n26862 ;
  assign n26864 = n26287 | n26863 ;
  assign n26865 = x5 | n26864 ;
  assign n26866 = x5 & n26864 ;
  assign n36254 = ~n26866 ;
  assign n26867 = n26865 & n36254 ;
  assign n36255 = ~n26860 ;
  assign n26868 = n36255 & n26867 ;
  assign n36256 = ~n26867 ;
  assign n26869 = n26860 & n36256 ;
  assign n26870 = n26868 | n26869 ;
  assign n26871 = n26716 | n26870 ;
  assign n26872 = n26716 & n26870 ;
  assign n36257 = ~n26872 ;
  assign n26873 = n26871 & n36257 ;
  assign n26498 = n733 | n26279 ;
  assign n26874 = x2 & n26498 ;
  assign n36258 = ~n26873 ;
  assign n26875 = n36258 & n26874 ;
  assign n36259 = ~n26874 ;
  assign n26876 = n26873 & n36259 ;
  assign n26877 = n26875 | n26876 ;
  assign n36260 = ~n26687 ;
  assign n26878 = n36260 & n26689 ;
  assign n36261 = ~n26689 ;
  assign n26879 = n26687 & n36261 ;
  assign n36262 = ~n26879 ;
  assign n26880 = n26710 & n36262 ;
  assign n26881 = n26878 | n26880 ;
  assign n26882 = n26877 | n26881 ;
  assign n26883 = n26877 & n26881 ;
  assign n36263 = ~n26883 ;
  assign n26884 = n26882 & n36263 ;
  assign n36264 = ~n26715 ;
  assign n26885 = n36264 & n26884 ;
  assign n36265 = ~n26884 ;
  assign n26886 = n26715 & n36265 ;
  assign n29905 = n26885 | n26886 ;
  assign n36266 = ~n26870 ;
  assign n26887 = n26716 & n36266 ;
  assign n26888 = n26868 | n26887 ;
  assign n26889 = n26840 | n26842 ;
  assign n36267 = ~n26839 ;
  assign n26890 = n36267 & n26889 ;
  assign n26891 = n26816 & n26827 ;
  assign n36268 = ~n26891 ;
  assign n26892 = n26826 & n36268 ;
  assign n24173 = n5937 & n24168 ;
  assign n23291 = n5994 & n35467 ;
  assign n24120 = n5970 & n35458 ;
  assign n26893 = n23291 | n24120 ;
  assign n26894 = n6018 & n24080 ;
  assign n26895 = n26893 | n26894 ;
  assign n26896 = n24173 | n26895 ;
  assign n36269 = ~n26896 ;
  assign n26897 = x14 & n36269 ;
  assign n26898 = n30547 & n26896 ;
  assign n26899 = n26897 | n26898 ;
  assign n26900 = n131 | n870 ;
  assign n26901 = n3008 | n4964 ;
  assign n26902 = n26900 | n26901 ;
  assign n26903 = n2622 | n26902 ;
  assign n36270 = ~n684 ;
  assign n26904 = n145 & n36270 ;
  assign n26905 = n996 | n1252 ;
  assign n36271 = ~n26905 ;
  assign n26906 = n26904 & n36271 ;
  assign n26907 = n535 | n696 ;
  assign n36272 = ~n26907 ;
  assign n26908 = n26906 & n36272 ;
  assign n26909 = n853 | n1305 ;
  assign n36273 = ~n26909 ;
  assign n26910 = n26908 & n36273 ;
  assign n36274 = ~n166 ;
  assign n26911 = n36274 & n26910 ;
  assign n36275 = ~n26903 ;
  assign n26912 = n36275 & n26911 ;
  assign n26913 = n1110 | n1892 ;
  assign n26914 = n2282 | n26913 ;
  assign n26915 = n26328 | n26914 ;
  assign n26916 = n26544 | n26915 ;
  assign n26917 = n801 | n26916 ;
  assign n26918 = n2359 | n2965 ;
  assign n26919 = n26917 | n26918 ;
  assign n36276 = ~n26919 ;
  assign n26920 = n26912 & n36276 ;
  assign n20525 = n889 & n34442 ;
  assign n20071 = n3311 & n20067 ;
  assign n20114 = n3329 & n34354 ;
  assign n26921 = n20071 | n20114 ;
  assign n26922 = n3343 & n20527 ;
  assign n26923 = n26921 | n26922 ;
  assign n26924 = n20525 | n26923 ;
  assign n36277 = ~n26924 ;
  assign n26925 = n26920 & n36277 ;
  assign n36278 = ~n26920 ;
  assign n26926 = n36278 & n26924 ;
  assign n26927 = n26925 | n26926 ;
  assign n36279 = ~n26732 ;
  assign n26928 = n36279 & n26736 ;
  assign n26929 = n26741 | n26928 ;
  assign n26930 = n26927 | n26929 ;
  assign n26931 = n26927 & n26929 ;
  assign n36280 = ~n26931 ;
  assign n26932 = n26930 & n36280 ;
  assign n20843 = n895 & n20833 ;
  assign n19795 = n2849 & n34519 ;
  assign n19821 = n2861 & n34355 ;
  assign n26933 = n19795 | n19821 ;
  assign n26934 = n894 & n20845 ;
  assign n26935 = n26933 | n26934 ;
  assign n26936 = n20843 | n26935 ;
  assign n26937 = x29 | n26936 ;
  assign n26938 = x29 & n26936 ;
  assign n36281 = ~n26938 ;
  assign n26939 = n26937 & n36281 ;
  assign n26940 = n26932 & n26939 ;
  assign n26941 = n26932 | n26939 ;
  assign n36282 = ~n26940 ;
  assign n26942 = n36282 & n26941 ;
  assign n26943 = n26751 | n26754 ;
  assign n26944 = n26942 | n26943 ;
  assign n26945 = n26942 & n26943 ;
  assign n36283 = ~n26945 ;
  assign n26946 = n26944 & n36283 ;
  assign n21071 = n3791 & n34598 ;
  assign n19723 = n3802 & n34363 ;
  assign n19747 = n209 & n34520 ;
  assign n26947 = n19723 | n19747 ;
  assign n26948 = n3818 & n34349 ;
  assign n26949 = n26947 | n26948 ;
  assign n26950 = n21071 | n26949 ;
  assign n26951 = x26 | n26950 ;
  assign n26952 = x26 & n26950 ;
  assign n36284 = ~n26952 ;
  assign n26953 = n26951 & n36284 ;
  assign n26954 = n26946 & n26953 ;
  assign n26955 = n26946 | n26953 ;
  assign n36285 = ~n26954 ;
  assign n26956 = n36285 & n26955 ;
  assign n26957 = n26764 | n26769 ;
  assign n26958 = n26956 | n26957 ;
  assign n26959 = n26956 & n26957 ;
  assign n36286 = ~n26959 ;
  assign n26960 = n26958 & n36286 ;
  assign n21857 = n4135 & n21848 ;
  assign n19670 = n4185 & n34360 ;
  assign n21771 = n4148 & n34803 ;
  assign n26961 = n19670 | n21771 ;
  assign n26962 = n4165 & n21753 ;
  assign n26963 = n26961 | n26962 ;
  assign n26964 = n21857 | n26963 ;
  assign n26965 = x23 | n26964 ;
  assign n26966 = x23 & n26964 ;
  assign n36287 = ~n26966 ;
  assign n26967 = n26965 & n36287 ;
  assign n26968 = n26960 & n26967 ;
  assign n26969 = n26960 | n26967 ;
  assign n36288 = ~n26968 ;
  assign n26970 = n36288 & n26969 ;
  assign n26971 = n26779 | n26784 ;
  assign n26972 = n26970 | n26971 ;
  assign n26973 = n26970 & n26971 ;
  assign n36289 = ~n26973 ;
  assign n26974 = n26972 & n36289 ;
  assign n22623 = n4686 & n35030 ;
  assign n21734 = n4726 & n21729 ;
  assign n22542 = n4706 & n35018 ;
  assign n26975 = n21734 | n22542 ;
  assign n26976 = n4748 & n22533 ;
  assign n26977 = n26975 | n26976 ;
  assign n26978 = n22623 | n26977 ;
  assign n26979 = x20 | n26978 ;
  assign n26980 = x20 & n26978 ;
  assign n36290 = ~n26980 ;
  assign n26981 = n26979 & n36290 ;
  assign n36291 = ~n26974 ;
  assign n26982 = n36291 & n26981 ;
  assign n36292 = ~n26981 ;
  assign n26983 = n26974 & n36292 ;
  assign n26984 = n26982 | n26983 ;
  assign n26985 = n26796 | n26798 ;
  assign n36293 = ~n26795 ;
  assign n26986 = n36293 & n26985 ;
  assign n36294 = ~n26984 ;
  assign n26987 = n36294 & n26986 ;
  assign n36295 = ~n26986 ;
  assign n26988 = n26984 & n36295 ;
  assign n26989 = n26987 | n26988 ;
  assign n23410 = n37300 & n35252 ;
  assign n22524 = n5166 & n35020 ;
  assign n23355 = n5144 & n23339 ;
  assign n26990 = n22524 | n23355 ;
  assign n26991 = n5191 & n35254 ;
  assign n26992 = n26990 | n26991 ;
  assign n26993 = n23410 | n26992 ;
  assign n26994 = x17 | n26993 ;
  assign n26995 = x17 & n26993 ;
  assign n36296 = ~n26995 ;
  assign n26996 = n26994 & n36296 ;
  assign n36297 = ~n26989 ;
  assign n26997 = n36297 & n26996 ;
  assign n36298 = ~n26996 ;
  assign n26998 = n26989 & n36298 ;
  assign n26999 = n26997 | n26998 ;
  assign n27000 = n26808 & n26810 ;
  assign n27001 = n26814 | n27000 ;
  assign n27002 = n26999 | n27001 ;
  assign n27003 = n26999 & n27001 ;
  assign n36299 = ~n27003 ;
  assign n27004 = n27002 & n36299 ;
  assign n36300 = ~n26899 ;
  assign n27005 = n36300 & n27004 ;
  assign n36301 = ~n27004 ;
  assign n27006 = n26899 & n36301 ;
  assign n27007 = n27005 | n27006 ;
  assign n36302 = ~n27007 ;
  assign n27008 = n26892 & n36302 ;
  assign n36303 = ~n26892 ;
  assign n27009 = n36303 & n27007 ;
  assign n27010 = n27008 | n27009 ;
  assign n25323 = n6272 & n35670 ;
  assign n24064 = n6244 & n24057 ;
  assign n24694 = n6190 & n24676 ;
  assign n27011 = n24064 | n24694 ;
  assign n27012 = n6217 & n35663 ;
  assign n27013 = n27011 | n27012 ;
  assign n27014 = n25323 | n27013 ;
  assign n27015 = x11 | n27014 ;
  assign n27016 = x11 & n27014 ;
  assign n36304 = ~n27016 ;
  assign n27017 = n27015 & n36304 ;
  assign n36305 = ~n27010 ;
  assign n27018 = n36305 & n27017 ;
  assign n36306 = ~n27017 ;
  assign n27019 = n27010 & n36306 ;
  assign n27020 = n27018 | n27019 ;
  assign n36307 = ~n27020 ;
  assign n27021 = n26890 & n36307 ;
  assign n36308 = ~n26890 ;
  assign n27022 = n36308 & n27020 ;
  assign n27023 = n27021 | n27022 ;
  assign n25829 = n7068 & n35910 ;
  assign n24821 = n7041 & n24815 ;
  assign n25405 = n69 & n35784 ;
  assign n27024 = n24821 | n25405 ;
  assign n27025 = n7017 & n25796 ;
  assign n27026 = n27024 | n27025 ;
  assign n27027 = n25829 | n27026 ;
  assign n27028 = x8 | n27027 ;
  assign n27029 = x8 & n27027 ;
  assign n36309 = ~n27029 ;
  assign n27030 = n27028 & n36309 ;
  assign n36310 = ~n27023 ;
  assign n27031 = n36310 & n27030 ;
  assign n36311 = ~n27030 ;
  assign n27032 = n27023 & n36311 ;
  assign n27033 = n27031 | n27032 ;
  assign n27034 = n26855 | n26857 ;
  assign n36312 = ~n26854 ;
  assign n27035 = n36312 & n27034 ;
  assign n27036 = n27033 | n27035 ;
  assign n27037 = n27033 & n27035 ;
  assign n36313 = ~n27037 ;
  assign n27038 = n27036 & n36313 ;
  assign n26489 = n8157 & n36130 ;
  assign n26046 = n8195 & n26039 ;
  assign n26474 = n740 & n26278 ;
  assign n27039 = n26046 | n26474 ;
  assign n27040 = n9052 & n36131 ;
  assign n27041 = n27039 | n27040 ;
  assign n27042 = n26489 | n27041 ;
  assign n27043 = x5 | n27042 ;
  assign n27044 = x5 & n27042 ;
  assign n36314 = ~n27044 ;
  assign n27045 = n27043 & n36314 ;
  assign n27046 = x2 & n27045 ;
  assign n27047 = x2 | n27045 ;
  assign n36315 = ~n27046 ;
  assign n27048 = n36315 & n27047 ;
  assign n27049 = n27038 & n27048 ;
  assign n27050 = n27038 | n27048 ;
  assign n36316 = ~n27049 ;
  assign n27051 = n36316 & n27050 ;
  assign n27052 = n26888 & n27051 ;
  assign n27053 = n26888 | n27051 ;
  assign n36317 = ~n27052 ;
  assign n27054 = n36317 & n27053 ;
  assign n36318 = ~n26876 ;
  assign n27055 = n36318 & n26882 ;
  assign n27056 = n27054 & n27055 ;
  assign n27057 = n27054 | n27055 ;
  assign n36319 = ~n27056 ;
  assign n27058 = n36319 & n27057 ;
  assign n27059 = n26886 & n27058 ;
  assign n29903 = n26886 | n27058 ;
  assign n36320 = ~n27059 ;
  assign n29904 = n36320 & n29903 ;
  assign n36321 = ~n27058 ;
  assign n27060 = n26886 & n36321 ;
  assign n27061 = n1469 | n1497 ;
  assign n27062 = n2326 | n11643 ;
  assign n27063 = n27061 | n27062 ;
  assign n1974 = n249 | n312 ;
  assign n27064 = n334 | n377 ;
  assign n27065 = n1974 | n27064 ;
  assign n27066 = n15348 | n27065 ;
  assign n27067 = n27063 | n27066 ;
  assign n27068 = n1807 | n27067 ;
  assign n36322 = ~n27068 ;
  assign n27069 = n23113 & n36322 ;
  assign n27070 = n2004 | n5605 ;
  assign n27071 = n22977 | n27070 ;
  assign n27072 = n5834 | n27071 ;
  assign n36323 = ~n27072 ;
  assign n27073 = n27069 & n36323 ;
  assign n27074 = n30152 & n27073 ;
  assign n36324 = ~n4973 ;
  assign n27075 = n36324 & n27074 ;
  assign n27076 = n30049 & n27075 ;
  assign n36325 = ~n27075 ;
  assign n27077 = x2 & n36325 ;
  assign n27078 = n27076 | n27077 ;
  assign n20784 = n889 & n34511 ;
  assign n19845 = n3329 & n19824 ;
  assign n20115 = n3311 & n34354 ;
  assign n27079 = n19845 | n20115 ;
  assign n27080 = n3343 & n34513 ;
  assign n27081 = n27079 | n27080 ;
  assign n27082 = n20784 | n27081 ;
  assign n27083 = n27078 | n27082 ;
  assign n27084 = n27078 & n27082 ;
  assign n36326 = ~n27084 ;
  assign n27085 = n27083 & n36326 ;
  assign n20815 = n895 & n20805 ;
  assign n19771 = n2849 & n19752 ;
  assign n19796 = n2861 & n34519 ;
  assign n27086 = n19771 | n19796 ;
  assign n27087 = n894 & n34520 ;
  assign n27088 = n27086 | n27087 ;
  assign n27089 = n20815 | n27088 ;
  assign n27090 = x29 | n27089 ;
  assign n27091 = x29 & n27089 ;
  assign n36327 = ~n27091 ;
  assign n27092 = n27090 & n36327 ;
  assign n36328 = ~n26925 ;
  assign n27093 = n36328 & n26930 ;
  assign n27094 = n27092 & n27093 ;
  assign n27095 = n27092 | n27093 ;
  assign n36329 = ~n27094 ;
  assign n27096 = n36329 & n27095 ;
  assign n36330 = ~n27085 ;
  assign n27097 = n36330 & n27096 ;
  assign n36331 = ~n27096 ;
  assign n27099 = n27085 & n36331 ;
  assign n27100 = n27097 | n27099 ;
  assign n20156 = n3791 & n34362 ;
  assign n19700 = n3802 & n34349 ;
  assign n19726 = n209 & n34363 ;
  assign n27101 = n19700 | n19726 ;
  assign n27102 = n3818 & n34365 ;
  assign n27103 = n27101 | n27102 ;
  assign n27104 = n20156 | n27103 ;
  assign n27105 = x26 | n27104 ;
  assign n27106 = x26 & n27104 ;
  assign n36332 = ~n27106 ;
  assign n27107 = n27105 & n36332 ;
  assign n27108 = n27100 & n27107 ;
  assign n27109 = n27100 | n27107 ;
  assign n36333 = ~n27108 ;
  assign n27110 = n36333 & n27109 ;
  assign n36334 = ~n26939 ;
  assign n27111 = n26932 & n36334 ;
  assign n36335 = ~n27111 ;
  assign n27112 = n26944 & n36335 ;
  assign n36336 = ~n27110 ;
  assign n27113 = n36336 & n27112 ;
  assign n36337 = ~n27112 ;
  assign n27114 = n27110 & n36337 ;
  assign n27115 = n27113 | n27114 ;
  assign n21793 = n4135 & n34802 ;
  assign n21772 = n4185 & n34803 ;
  assign n21806 = n4148 & n21753 ;
  assign n27116 = n21772 | n21806 ;
  assign n27117 = n4165 & n21804 ;
  assign n27118 = n27116 | n27117 ;
  assign n27119 = n21793 | n27118 ;
  assign n27120 = x23 | n27119 ;
  assign n27121 = x23 & n27119 ;
  assign n36338 = ~n27121 ;
  assign n27122 = n27120 & n36338 ;
  assign n36339 = ~n27115 ;
  assign n27123 = n36339 & n27122 ;
  assign n36340 = ~n27122 ;
  assign n27124 = n27115 & n36340 ;
  assign n27125 = n27123 | n27124 ;
  assign n36341 = ~n26953 ;
  assign n27126 = n26946 & n36341 ;
  assign n36342 = ~n27126 ;
  assign n27127 = n26958 & n36342 ;
  assign n36343 = ~n27125 ;
  assign n27128 = n36343 & n27127 ;
  assign n36344 = ~n27127 ;
  assign n27129 = n27125 & n36344 ;
  assign n27130 = n27128 | n27129 ;
  assign n22572 = n4686 & n35022 ;
  assign n22547 = n4726 & n35018 ;
  assign n22593 = n4706 & n22533 ;
  assign n27131 = n22547 | n22593 ;
  assign n27132 = n4748 & n35020 ;
  assign n27133 = n27131 | n27132 ;
  assign n27134 = n22572 | n27133 ;
  assign n27135 = x20 | n27134 ;
  assign n27136 = x20 & n27134 ;
  assign n36345 = ~n27136 ;
  assign n27137 = n27135 & n36345 ;
  assign n36346 = ~n27130 ;
  assign n27138 = n36346 & n27137 ;
  assign n36347 = ~n27137 ;
  assign n27139 = n27130 & n36347 ;
  assign n27140 = n27138 | n27139 ;
  assign n36348 = ~n26960 ;
  assign n27141 = n36348 & n26967 ;
  assign n36349 = ~n26970 ;
  assign n27142 = n36349 & n26971 ;
  assign n27143 = n27141 | n27142 ;
  assign n27144 = n27140 | n27143 ;
  assign n27145 = n27140 & n27143 ;
  assign n36350 = ~n27145 ;
  assign n27146 = n27144 & n36350 ;
  assign n23378 = n37300 & n23372 ;
  assign n23317 = n5144 & n35244 ;
  assign n23356 = n5166 & n23339 ;
  assign n27147 = n23317 | n23356 ;
  assign n27148 = n5191 & n35246 ;
  assign n27149 = n27147 | n27148 ;
  assign n27150 = n23378 | n27149 ;
  assign n27151 = x17 | n27150 ;
  assign n27152 = x17 & n27150 ;
  assign n36351 = ~n27152 ;
  assign n27153 = n27151 & n36351 ;
  assign n27154 = n27146 & n27153 ;
  assign n27155 = n27146 | n27153 ;
  assign n36352 = ~n27154 ;
  assign n27156 = n36352 & n27155 ;
  assign n27157 = n26982 | n26987 ;
  assign n27158 = n27156 | n27157 ;
  assign n27159 = n27156 & n27157 ;
  assign n36353 = ~n27159 ;
  assign n27160 = n27158 & n36353 ;
  assign n24144 = n5937 & n35457 ;
  assign n24089 = n5970 & n24080 ;
  assign n24110 = n5994 & n35458 ;
  assign n27161 = n24089 | n24110 ;
  assign n27162 = n6018 & n24151 ;
  assign n27163 = n27161 | n27162 ;
  assign n27164 = n24144 | n27163 ;
  assign n27165 = x14 | n27164 ;
  assign n27166 = x14 & n27164 ;
  assign n36354 = ~n27166 ;
  assign n27167 = n27165 & n36354 ;
  assign n36355 = ~n27160 ;
  assign n27168 = n36355 & n27167 ;
  assign n36356 = ~n27167 ;
  assign n27169 = n27160 & n36356 ;
  assign n27170 = n27168 | n27169 ;
  assign n36357 = ~n26998 ;
  assign n27171 = n36357 & n27002 ;
  assign n36358 = ~n27170 ;
  assign n27172 = n36358 & n27171 ;
  assign n36359 = ~n27171 ;
  assign n27173 = n27170 & n36359 ;
  assign n27174 = n27172 | n27173 ;
  assign n24875 = n6272 & n35662 ;
  assign n24692 = n6244 & n24676 ;
  assign n24844 = n6190 & n35663 ;
  assign n27175 = n24692 | n24844 ;
  assign n27176 = n6217 & n24815 ;
  assign n27177 = n27175 | n27176 ;
  assign n27178 = n24875 | n27177 ;
  assign n27179 = x11 | n27178 ;
  assign n27180 = x11 & n27178 ;
  assign n36360 = ~n27180 ;
  assign n27181 = n27179 & n36360 ;
  assign n36361 = ~n27174 ;
  assign n27182 = n36361 & n27181 ;
  assign n36362 = ~n27181 ;
  assign n27183 = n27174 & n36362 ;
  assign n27184 = n27182 | n27183 ;
  assign n27185 = n27006 | n27008 ;
  assign n36363 = ~n27185 ;
  assign n27186 = n27184 & n36363 ;
  assign n36364 = ~n27184 ;
  assign n27187 = n36364 & n27185 ;
  assign n27188 = n27186 | n27187 ;
  assign n26070 = n7068 & n26065 ;
  assign n25395 = n7041 & n35784 ;
  assign n25807 = n69 & n25796 ;
  assign n27189 = n25395 | n25807 ;
  assign n27190 = n7017 & n26039 ;
  assign n27191 = n27189 | n27190 ;
  assign n27192 = n26070 | n27191 ;
  assign n27193 = x8 | n27192 ;
  assign n27194 = x8 & n27192 ;
  assign n36365 = ~n27194 ;
  assign n27195 = n27193 & n36365 ;
  assign n27196 = n27188 & n27195 ;
  assign n27197 = n27188 | n27195 ;
  assign n36366 = ~n27196 ;
  assign n27198 = n36366 & n27197 ;
  assign n27199 = n27018 | n27021 ;
  assign n36367 = ~n27199 ;
  assign n27200 = n27198 & n36367 ;
  assign n36368 = ~n27198 ;
  assign n27201 = n36368 & n27199 ;
  assign n27202 = n27200 | n27201 ;
  assign n26697 = n8157 & n36192 ;
  assign n27203 = n8195 & n26278 ;
  assign n27204 = n740 & n36131 ;
  assign n27205 = n27203 | n27204 ;
  assign n27206 = n26697 | n27205 ;
  assign n36369 = ~n27206 ;
  assign n27207 = x5 & n36369 ;
  assign n27208 = n30053 & n27206 ;
  assign n27209 = n27207 | n27208 ;
  assign n27210 = n27202 | n27209 ;
  assign n27211 = n27202 & n27209 ;
  assign n36370 = ~n27211 ;
  assign n27212 = n27210 & n36370 ;
  assign n36371 = ~n27032 ;
  assign n27213 = n36371 & n27036 ;
  assign n27214 = n27212 | n27213 ;
  assign n27215 = n27212 & n27213 ;
  assign n36372 = ~n27215 ;
  assign n27216 = n27214 & n36372 ;
  assign n27217 = n27047 & n36316 ;
  assign n36373 = ~n27216 ;
  assign n27218 = n36373 & n27217 ;
  assign n36374 = ~n27217 ;
  assign n27219 = n27216 & n36374 ;
  assign n27220 = n27218 | n27219 ;
  assign n36375 = ~n26888 ;
  assign n27221 = n36375 & n27051 ;
  assign n36376 = ~n27221 ;
  assign n27222 = n27055 & n36376 ;
  assign n36377 = ~n27051 ;
  assign n27223 = n26888 & n36377 ;
  assign n27224 = n27222 | n27223 ;
  assign n27225 = n27220 | n27224 ;
  assign n27226 = n27220 & n27224 ;
  assign n36378 = ~n27226 ;
  assign n27227 = n27225 & n36378 ;
  assign n27228 = n27060 & n27227 ;
  assign n29901 = n27060 | n27227 ;
  assign n36379 = ~n27228 ;
  assign n29902 = n36379 & n29901 ;
  assign n36380 = ~n27227 ;
  assign n27229 = n27060 & n36380 ;
  assign n36381 = ~n27195 ;
  assign n27230 = n27188 & n36381 ;
  assign n27231 = n27198 | n27199 ;
  assign n36382 = ~n27230 ;
  assign n27232 = n36382 & n27231 ;
  assign n36383 = ~n27146 ;
  assign n27233 = n36383 & n27153 ;
  assign n36384 = ~n27156 ;
  assign n27234 = n36384 & n27157 ;
  assign n27235 = n27233 | n27234 ;
  assign n23442 = n4686 & n35262 ;
  assign n22525 = n4706 & n35020 ;
  assign n22594 = n4726 & n22533 ;
  assign n27236 = n22525 | n22594 ;
  assign n27237 = n4748 & n23444 ;
  assign n27238 = n27236 | n27237 ;
  assign n27239 = n23442 | n27238 ;
  assign n27240 = x20 | n27239 ;
  assign n27241 = x20 & n27239 ;
  assign n36385 = ~n27241 ;
  assign n27242 = n27240 & n36385 ;
  assign n27243 = n1211 | n1230 ;
  assign n27244 = n1718 | n3016 ;
  assign n27245 = n27243 | n27244 ;
  assign n27246 = n235 | n439 ;
  assign n27247 = n141 | n27246 ;
  assign n27248 = n949 | n27247 ;
  assign n27249 = n1726 | n2305 ;
  assign n27250 = n27248 | n27249 ;
  assign n27251 = n27245 | n27250 ;
  assign n27252 = n348 | n501 ;
  assign n27253 = n2174 | n27252 ;
  assign n27254 = n13605 | n27253 ;
  assign n27255 = n2394 | n3493 ;
  assign n27256 = n3682 | n20450 ;
  assign n27257 = n27255 | n27256 ;
  assign n27258 = n1098 | n27257 ;
  assign n27259 = n27254 | n27258 ;
  assign n27260 = n27251 | n27259 ;
  assign n27261 = n2001 | n27260 ;
  assign n27262 = n13568 | n27261 ;
  assign n27263 = x2 | n27262 ;
  assign n27264 = x2 & n27262 ;
  assign n36386 = ~n27264 ;
  assign n27265 = n27263 & n36386 ;
  assign n36387 = ~n27078 ;
  assign n27266 = n36387 & n27082 ;
  assign n27267 = n27077 | n27266 ;
  assign n36388 = ~n27267 ;
  assign n27268 = n27265 & n36388 ;
  assign n36389 = ~n27265 ;
  assign n27269 = n36389 & n27267 ;
  assign n27270 = n27268 | n27269 ;
  assign n20873 = n889 & n20863 ;
  assign n19822 = n3329 & n34355 ;
  assign n19836 = n3311 & n19824 ;
  assign n27271 = n19822 | n19836 ;
  assign n27272 = n3343 & n34536 ;
  assign n27273 = n27271 | n27272 ;
  assign n27274 = n20873 | n27273 ;
  assign n36390 = ~n27274 ;
  assign n27275 = n27270 & n36390 ;
  assign n36391 = ~n27270 ;
  assign n27276 = n36391 & n27274 ;
  assign n27277 = n27275 | n27276 ;
  assign n27098 = n27085 & n27096 ;
  assign n36392 = ~n27098 ;
  assign n27278 = n27095 & n36392 ;
  assign n27279 = n27277 & n27278 ;
  assign n27280 = n27277 | n27278 ;
  assign n36393 = ~n27279 ;
  assign n27281 = n36393 & n27280 ;
  assign n21105 = n895 & n34603 ;
  assign n19748 = n2849 & n34520 ;
  assign n19772 = n2861 & n19752 ;
  assign n27282 = n19748 | n19772 ;
  assign n27283 = n894 & n34596 ;
  assign n27284 = n27282 | n27283 ;
  assign n27285 = n21105 | n27284 ;
  assign n27286 = x29 | n27285 ;
  assign n27287 = x29 & n27285 ;
  assign n36394 = ~n27287 ;
  assign n27288 = n27286 & n36394 ;
  assign n36395 = ~n27281 ;
  assign n27289 = n36395 & n27288 ;
  assign n36396 = ~n27288 ;
  assign n27290 = n27281 & n36396 ;
  assign n27291 = n27289 | n27290 ;
  assign n21880 = n3791 & n34817 ;
  assign n19677 = n3802 & n34360 ;
  assign n19701 = n209 & n34349 ;
  assign n27292 = n19677 | n19701 ;
  assign n27293 = n3818 & n34803 ;
  assign n27294 = n27292 | n27293 ;
  assign n27295 = n21880 | n27294 ;
  assign n36397 = ~n27295 ;
  assign n27296 = x26 & n36397 ;
  assign n27297 = n30019 & n27295 ;
  assign n27298 = n27296 | n27297 ;
  assign n36398 = ~n27298 ;
  assign n27299 = n27291 & n36398 ;
  assign n36399 = ~n27291 ;
  assign n27300 = n36399 & n27298 ;
  assign n27301 = n27299 | n27300 ;
  assign n36400 = ~n27107 ;
  assign n27302 = n27100 & n36400 ;
  assign n27303 = n27110 | n27112 ;
  assign n36401 = ~n27302 ;
  assign n27304 = n36401 & n27303 ;
  assign n36402 = ~n27301 ;
  assign n27305 = n36402 & n27304 ;
  assign n36403 = ~n27304 ;
  assign n27306 = n27301 & n36403 ;
  assign n27307 = n27305 | n27306 ;
  assign n22646 = n4135 & n35035 ;
  assign n21731 = n4148 & n21729 ;
  assign n21809 = n4185 & n21753 ;
  assign n27308 = n21731 | n21809 ;
  assign n27309 = n4165 & n35018 ;
  assign n27310 = n27308 | n27309 ;
  assign n27311 = n22646 | n27310 ;
  assign n36404 = ~n27311 ;
  assign n27312 = x23 & n36404 ;
  assign n27313 = n30030 & n27311 ;
  assign n27314 = n27312 | n27313 ;
  assign n36405 = ~n27314 ;
  assign n27315 = n27307 & n36405 ;
  assign n36406 = ~n27307 ;
  assign n27316 = n36406 & n27314 ;
  assign n27317 = n27315 | n27316 ;
  assign n27318 = n27123 | n27128 ;
  assign n27319 = n27317 | n27318 ;
  assign n27320 = n27317 & n27318 ;
  assign n36407 = ~n27320 ;
  assign n27321 = n27319 & n36407 ;
  assign n27322 = n27242 & n27321 ;
  assign n27323 = n27242 | n27321 ;
  assign n36408 = ~n27322 ;
  assign n27324 = n36408 & n27323 ;
  assign n24200 = n37300 & n35472 ;
  assign n23307 = n5144 & n35467 ;
  assign n23323 = n5166 & n35244 ;
  assign n27325 = n23307 | n23323 ;
  assign n27326 = n5191 & n35465 ;
  assign n27327 = n27325 | n27326 ;
  assign n27328 = n24200 | n27327 ;
  assign n27329 = x17 | n27328 ;
  assign n27330 = x17 & n27328 ;
  assign n36409 = ~n27330 ;
  assign n27331 = n27329 & n36409 ;
  assign n27332 = n27324 & n27331 ;
  assign n27333 = n27324 | n27331 ;
  assign n36410 = ~n27332 ;
  assign n27334 = n36410 & n27333 ;
  assign n36411 = ~n27139 ;
  assign n27335 = n36411 & n27144 ;
  assign n27336 = n27334 & n27335 ;
  assign n27337 = n27334 | n27335 ;
  assign n36412 = ~n27336 ;
  assign n27338 = n36412 & n27337 ;
  assign n25292 = n5937 & n25288 ;
  assign n24062 = n5970 & n24057 ;
  assign n24092 = n5994 & n24080 ;
  assign n27339 = n24062 | n24092 ;
  assign n27340 = n6018 & n24676 ;
  assign n27341 = n27339 | n27340 ;
  assign n27342 = n25292 | n27341 ;
  assign n27343 = x14 | n27342 ;
  assign n27344 = x14 & n27342 ;
  assign n36413 = ~n27344 ;
  assign n27345 = n27343 & n36413 ;
  assign n27346 = n27338 & n27345 ;
  assign n27347 = n27338 | n27345 ;
  assign n36414 = ~n27346 ;
  assign n27348 = n36414 & n27347 ;
  assign n36415 = ~n27235 ;
  assign n27349 = n36415 & n27348 ;
  assign n36416 = ~n27348 ;
  assign n27350 = n27235 & n36416 ;
  assign n27351 = n27349 | n27350 ;
  assign n25425 = n6272 & n35785 ;
  assign n24818 = n6190 & n24815 ;
  assign n24843 = n6244 & n35663 ;
  assign n27352 = n24818 | n24843 ;
  assign n27353 = n6217 & n35784 ;
  assign n27354 = n27352 | n27353 ;
  assign n27355 = n25425 | n27354 ;
  assign n27356 = x11 | n27355 ;
  assign n27357 = x11 & n27355 ;
  assign n36417 = ~n27357 ;
  assign n27358 = n27356 & n36417 ;
  assign n36418 = ~n27351 ;
  assign n27359 = n36418 & n27358 ;
  assign n36419 = ~n27358 ;
  assign n27360 = n27351 & n36419 ;
  assign n27361 = n27359 | n27360 ;
  assign n27362 = n27168 | n27172 ;
  assign n36420 = ~n27362 ;
  assign n27363 = n27361 & n36420 ;
  assign n36421 = ~n27361 ;
  assign n27364 = n36421 & n27362 ;
  assign n27365 = n27363 | n27364 ;
  assign n26288 = n7068 & n26284 ;
  assign n25800 = n7041 & n25796 ;
  assign n26051 = n69 & n26039 ;
  assign n27366 = n25800 | n26051 ;
  assign n27367 = n7017 & n26278 ;
  assign n27368 = n27366 | n27367 ;
  assign n27369 = n26288 | n27368 ;
  assign n27370 = x8 | n27369 ;
  assign n27371 = x8 & n27369 ;
  assign n36422 = ~n27371 ;
  assign n27372 = n27370 & n36422 ;
  assign n36423 = ~n27365 ;
  assign n27373 = n36423 & n27372 ;
  assign n36424 = ~n27372 ;
  assign n27374 = n27365 & n36424 ;
  assign n27375 = n27373 | n27374 ;
  assign n27376 = n27184 | n27185 ;
  assign n36425 = ~n27183 ;
  assign n27377 = n36425 & n27376 ;
  assign n27378 = n27375 & n27377 ;
  assign n27379 = n27375 | n27377 ;
  assign n36426 = ~n27378 ;
  assign n27380 = n36426 & n27379 ;
  assign n26499 = n735 & n36131 ;
  assign n27381 = n741 | n26279 ;
  assign n27382 = x5 & n27381 ;
  assign n27383 = n26499 | n27382 ;
  assign n27384 = n27380 | n27383 ;
  assign n27385 = n27380 & n27383 ;
  assign n36427 = ~n27385 ;
  assign n27386 = n27384 & n36427 ;
  assign n36428 = ~n27232 ;
  assign n27387 = n36428 & n27386 ;
  assign n36429 = ~n27386 ;
  assign n27388 = n27232 & n36429 ;
  assign n27389 = n27387 | n27388 ;
  assign n36430 = ~n27209 ;
  assign n27390 = n27202 & n36430 ;
  assign n36431 = ~n27390 ;
  assign n27391 = n27214 & n36431 ;
  assign n27392 = n27389 & n27391 ;
  assign n27393 = n27389 | n27391 ;
  assign n36432 = ~n27392 ;
  assign n27394 = n36432 & n27393 ;
  assign n36433 = ~n27219 ;
  assign n27395 = n36433 & n27224 ;
  assign n27396 = n27218 | n27395 ;
  assign n36434 = ~n27394 ;
  assign n27397 = n36434 & n27396 ;
  assign n36435 = ~n27396 ;
  assign n27398 = n27394 & n36435 ;
  assign n27399 = n27397 | n27398 ;
  assign n36436 = ~n27399 ;
  assign n27400 = n27229 & n36436 ;
  assign n36437 = ~n27229 ;
  assign n29899 = n36437 & n27399 ;
  assign n41 = n27400 | n29899 ;
  assign n27401 = n27229 & n27399 ;
  assign n27402 = n27392 | n27396 ;
  assign n27403 = n27393 & n27402 ;
  assign n25830 = n6272 & n35910 ;
  assign n24828 = n6244 & n24815 ;
  assign n25403 = n6190 & n35784 ;
  assign n27404 = n24828 | n25403 ;
  assign n27405 = n6217 & n25796 ;
  assign n27406 = n27404 | n27405 ;
  assign n27407 = n25830 | n27406 ;
  assign n27408 = x11 | n27407 ;
  assign n27409 = x11 & n27407 ;
  assign n36438 = ~n27409 ;
  assign n27410 = n27408 & n36438 ;
  assign n27411 = n921 | n1246 ;
  assign n27412 = n2426 | n27411 ;
  assign n27413 = n472 | n27412 ;
  assign n27414 = n11602 | n12954 ;
  assign n27415 = n27413 | n27414 ;
  assign n27416 = n270 | n320 ;
  assign n27417 = n383 | n2311 ;
  assign n27418 = n27416 | n27417 ;
  assign n27419 = n916 | n27418 ;
  assign n27420 = n1032 | n27419 ;
  assign n27421 = n3284 | n27420 ;
  assign n27422 = n27415 | n27421 ;
  assign n27423 = n4008 | n27422 ;
  assign n27424 = n2077 | n27423 ;
  assign n27425 = n3074 | n27424 ;
  assign n27426 = x2 | n27425 ;
  assign n27427 = x2 & n27425 ;
  assign n36439 = ~n27427 ;
  assign n27428 = n27426 & n36439 ;
  assign n27429 = n27263 & n27267 ;
  assign n27430 = n27264 | n27429 ;
  assign n36440 = ~n27430 ;
  assign n27431 = n27428 & n36440 ;
  assign n36441 = ~n27428 ;
  assign n27432 = n36441 & n27430 ;
  assign n27433 = n27431 | n27432 ;
  assign n20844 = n889 & n20833 ;
  assign n19797 = n3329 & n34519 ;
  assign n19802 = n3311 & n34355 ;
  assign n27434 = n19797 | n19802 ;
  assign n27435 = n3343 & n20845 ;
  assign n27436 = n27434 | n27435 ;
  assign n27437 = n20844 | n27436 ;
  assign n27438 = n27433 | n27437 ;
  assign n27439 = n27433 & n27437 ;
  assign n36442 = ~n27439 ;
  assign n27440 = n27438 & n36442 ;
  assign n27441 = n27270 | n27274 ;
  assign n36443 = ~n27278 ;
  assign n27442 = n27277 & n36443 ;
  assign n36444 = ~n27442 ;
  assign n27443 = n27441 & n36444 ;
  assign n27444 = n27440 & n27443 ;
  assign n27445 = n27440 | n27443 ;
  assign n36445 = ~n27444 ;
  assign n27446 = n36445 & n27445 ;
  assign n21075 = n895 & n34598 ;
  assign n19717 = n2849 & n34363 ;
  assign n19749 = n2861 & n34520 ;
  assign n27447 = n19717 | n19749 ;
  assign n27448 = n894 & n34349 ;
  assign n27449 = n27447 | n27448 ;
  assign n27450 = n21075 | n27449 ;
  assign n27451 = x29 | n27450 ;
  assign n27452 = x29 & n27450 ;
  assign n36446 = ~n27452 ;
  assign n27453 = n27451 & n36446 ;
  assign n36447 = ~n27446 ;
  assign n27454 = n36447 & n27453 ;
  assign n36448 = ~n27453 ;
  assign n27455 = n27446 & n36448 ;
  assign n27456 = n27454 | n27455 ;
  assign n21851 = n3791 & n21848 ;
  assign n19678 = n209 & n34360 ;
  assign n21764 = n3802 & n34803 ;
  assign n27457 = n19678 | n21764 ;
  assign n27458 = n3818 & n21753 ;
  assign n27459 = n27457 | n27458 ;
  assign n27460 = n21851 | n27459 ;
  assign n36449 = ~n27460 ;
  assign n27461 = x26 & n36449 ;
  assign n27462 = n30019 & n27460 ;
  assign n27463 = n27461 | n27462 ;
  assign n36450 = ~n27463 ;
  assign n27464 = n27456 & n36450 ;
  assign n36451 = ~n27456 ;
  assign n27465 = n36451 & n27463 ;
  assign n27466 = n27464 | n27465 ;
  assign n27467 = n27281 | n27288 ;
  assign n36452 = ~n27299 ;
  assign n27468 = n36452 & n27467 ;
  assign n36453 = ~n27466 ;
  assign n27469 = n36453 & n27468 ;
  assign n36454 = ~n27468 ;
  assign n27470 = n27466 & n36454 ;
  assign n27471 = n27469 | n27470 ;
  assign n22628 = n4135 & n35030 ;
  assign n21747 = n4185 & n21729 ;
  assign n22553 = n4148 & n35018 ;
  assign n27472 = n21747 | n22553 ;
  assign n27473 = n4165 & n22533 ;
  assign n27474 = n27472 | n27473 ;
  assign n27475 = n22628 | n27474 ;
  assign n36455 = ~n27475 ;
  assign n27476 = x23 & n36455 ;
  assign n27477 = n30030 & n27475 ;
  assign n27478 = n27476 | n27477 ;
  assign n36456 = ~n27478 ;
  assign n27479 = n27471 & n36456 ;
  assign n36457 = ~n27471 ;
  assign n27480 = n36457 & n27478 ;
  assign n27481 = n27479 | n27480 ;
  assign n27482 = n27301 | n27304 ;
  assign n36458 = ~n27315 ;
  assign n27483 = n36458 & n27482 ;
  assign n36459 = ~n27481 ;
  assign n27484 = n36459 & n27483 ;
  assign n36460 = ~n27483 ;
  assign n27485 = n27481 & n36460 ;
  assign n27486 = n27484 | n27485 ;
  assign n23411 = n4686 & n35252 ;
  assign n22527 = n4726 & n35020 ;
  assign n23357 = n4706 & n23339 ;
  assign n27487 = n22527 | n23357 ;
  assign n27488 = n4748 & n35254 ;
  assign n27489 = n27487 | n27488 ;
  assign n27490 = n23411 | n27489 ;
  assign n36461 = ~n27490 ;
  assign n27491 = x20 & n36461 ;
  assign n27492 = n30374 & n27490 ;
  assign n27493 = n27491 | n27492 ;
  assign n36462 = ~n27493 ;
  assign n27494 = n27486 & n36462 ;
  assign n36463 = ~n27486 ;
  assign n27495 = n36463 & n27493 ;
  assign n27496 = n27494 | n27495 ;
  assign n27497 = n27320 | n27322 ;
  assign n27498 = n27496 | n27497 ;
  assign n27499 = n27496 & n27497 ;
  assign n36464 = ~n27499 ;
  assign n27500 = n27498 & n36464 ;
  assign n24174 = n37300 & n24168 ;
  assign n23305 = n5166 & n35467 ;
  assign n24104 = n5144 & n35458 ;
  assign n27501 = n23305 | n24104 ;
  assign n27502 = n5191 & n24080 ;
  assign n27503 = n27501 | n27502 ;
  assign n27504 = n24174 | n27503 ;
  assign n36465 = ~n27504 ;
  assign n27505 = x17 & n36465 ;
  assign n27506 = n30580 & n27504 ;
  assign n27507 = n27505 | n27506 ;
  assign n36466 = ~n27507 ;
  assign n27508 = n27500 & n36466 ;
  assign n36467 = ~n27500 ;
  assign n27509 = n36467 & n27507 ;
  assign n27510 = n27508 | n27509 ;
  assign n25324 = n5937 & n35670 ;
  assign n24061 = n5994 & n24057 ;
  assign n24678 = n5970 & n24676 ;
  assign n27511 = n24061 | n24678 ;
  assign n27512 = n6018 & n35663 ;
  assign n27513 = n27511 | n27512 ;
  assign n27514 = n25324 | n27513 ;
  assign n27515 = x14 | n27514 ;
  assign n27516 = x14 & n27514 ;
  assign n36468 = ~n27516 ;
  assign n27517 = n27515 & n36468 ;
  assign n36469 = ~n27510 ;
  assign n27518 = n36469 & n27517 ;
  assign n36470 = ~n27517 ;
  assign n27519 = n27510 & n36470 ;
  assign n27520 = n27518 | n27519 ;
  assign n27521 = n27332 | n27336 ;
  assign n27522 = n27520 | n27521 ;
  assign n27523 = n27520 & n27521 ;
  assign n36471 = ~n27523 ;
  assign n27524 = n27522 & n36471 ;
  assign n27525 = n27410 & n27524 ;
  assign n27526 = n27410 | n27524 ;
  assign n36472 = ~n27525 ;
  assign n27527 = n36472 & n27526 ;
  assign n36473 = ~n27349 ;
  assign n27528 = n27347 & n36473 ;
  assign n27529 = n27527 & n27528 ;
  assign n27530 = n27527 | n27528 ;
  assign n36474 = ~n27529 ;
  assign n27531 = n36474 & n27530 ;
  assign n26491 = n7068 & n36130 ;
  assign n26045 = n7041 & n26039 ;
  assign n26476 = n69 & n26278 ;
  assign n27532 = n26045 | n26476 ;
  assign n27533 = n7017 & n36131 ;
  assign n27534 = n27532 | n27533 ;
  assign n27535 = n26491 | n27534 ;
  assign n27536 = x8 | n27535 ;
  assign n27537 = x8 & n27535 ;
  assign n36475 = ~n27537 ;
  assign n27538 = n27536 & n36475 ;
  assign n27539 = n27351 | n27358 ;
  assign n36476 = ~n27363 ;
  assign n27540 = n36476 & n27539 ;
  assign n27541 = n27538 & n27540 ;
  assign n27542 = n27538 | n27540 ;
  assign n36477 = ~n27541 ;
  assign n27543 = n36477 & n27542 ;
  assign n36478 = ~n27531 ;
  assign n27544 = n36478 & n27543 ;
  assign n36479 = ~n27543 ;
  assign n27545 = n27531 & n36479 ;
  assign n27546 = n27544 | n27545 ;
  assign n27547 = n27365 | n27372 ;
  assign n36480 = ~n27377 ;
  assign n27548 = n27375 & n36480 ;
  assign n36481 = ~n27548 ;
  assign n27549 = n27547 & n36481 ;
  assign n27550 = x5 | n27549 ;
  assign n27551 = x5 & n27549 ;
  assign n36482 = ~n27551 ;
  assign n27552 = n27550 & n36482 ;
  assign n36483 = ~n27546 ;
  assign n27553 = n36483 & n27552 ;
  assign n36484 = ~n27552 ;
  assign n27554 = n27546 & n36484 ;
  assign n27555 = n27553 | n27554 ;
  assign n27556 = n27232 & n27386 ;
  assign n27557 = n27385 | n27556 ;
  assign n27558 = n27555 | n27557 ;
  assign n27559 = n27555 & n27557 ;
  assign n36485 = ~n27559 ;
  assign n27560 = n27558 & n36485 ;
  assign n36486 = ~n27403 ;
  assign n27561 = n36486 & n27560 ;
  assign n36487 = ~n27560 ;
  assign n27562 = n27403 & n36487 ;
  assign n27563 = n27561 | n27562 ;
  assign n27564 = n27401 | n27563 ;
  assign n27565 = n27401 & n27563 ;
  assign n36488 = ~n27565 ;
  assign n42 = n27564 & n36488 ;
  assign n24145 = n37300 & n35457 ;
  assign n24081 = n5144 & n24080 ;
  assign n24119 = n5166 & n35458 ;
  assign n27566 = n24081 | n24119 ;
  assign n27567 = n5191 & n24151 ;
  assign n27568 = n27566 | n27567 ;
  assign n27569 = n24145 | n27568 ;
  assign n27570 = x17 | n27569 ;
  assign n27571 = x17 & n27569 ;
  assign n36489 = ~n27571 ;
  assign n27572 = n27570 & n36489 ;
  assign n36490 = ~n27431 ;
  assign n27573 = n27426 & n36490 ;
  assign n27574 = n2154 | n2962 ;
  assign n27575 = n4274 | n27574 ;
  assign n27576 = n356 | n1662 ;
  assign n27577 = n2768 | n2951 ;
  assign n27578 = n27576 | n27577 ;
  assign n27579 = n200 | n221 ;
  assign n27580 = n224 | n399 ;
  assign n27581 = n27579 | n27580 ;
  assign n27582 = n1411 | n27581 ;
  assign n27583 = n27578 | n27582 ;
  assign n27584 = n27575 | n27583 ;
  assign n27585 = n22246 | n27584 ;
  assign n27586 = n20256 | n27585 ;
  assign n27587 = n12836 | n27586 ;
  assign n27588 = n1680 | n27587 ;
  assign n36491 = ~n27588 ;
  assign n27589 = n4369 & n36491 ;
  assign n27590 = n30306 & n27588 ;
  assign n27591 = n27589 | n27590 ;
  assign n27592 = n27573 & n27591 ;
  assign n27593 = n27573 | n27591 ;
  assign n36492 = ~n27592 ;
  assign n27594 = n36492 & n27593 ;
  assign n20816 = n889 & n20805 ;
  assign n19755 = n3329 & n19752 ;
  assign n19798 = n3311 & n34519 ;
  assign n27595 = n19755 | n19798 ;
  assign n27596 = n3343 & n34520 ;
  assign n27597 = n27595 | n27596 ;
  assign n27598 = n20816 | n27597 ;
  assign n36493 = ~n27598 ;
  assign n27599 = n27594 & n36493 ;
  assign n36494 = ~n27594 ;
  assign n27600 = n36494 & n27598 ;
  assign n27601 = n27599 | n27600 ;
  assign n20150 = n895 & n34362 ;
  assign n19702 = n2849 & n34349 ;
  assign n19727 = n2861 & n34363 ;
  assign n27602 = n19702 | n19727 ;
  assign n27603 = n894 & n34365 ;
  assign n27604 = n27602 | n27603 ;
  assign n27605 = n20150 | n27604 ;
  assign n36495 = ~n27605 ;
  assign n27606 = x29 & n36495 ;
  assign n27607 = n30024 & n27605 ;
  assign n27608 = n27606 | n27607 ;
  assign n36496 = ~n27608 ;
  assign n27609 = n27601 & n36496 ;
  assign n36497 = ~n27601 ;
  assign n27610 = n36497 & n27608 ;
  assign n27611 = n27609 | n27610 ;
  assign n36498 = ~n27443 ;
  assign n27612 = n27440 & n36498 ;
  assign n36499 = ~n27612 ;
  assign n27613 = n27438 & n36499 ;
  assign n27614 = n27611 & n27613 ;
  assign n27615 = n27611 | n27613 ;
  assign n36500 = ~n27614 ;
  assign n27616 = n36500 & n27615 ;
  assign n21799 = n3791 & n34802 ;
  assign n21773 = n209 & n34803 ;
  assign n21822 = n3802 & n21753 ;
  assign n27617 = n21773 | n21822 ;
  assign n27618 = n3818 & n21804 ;
  assign n27619 = n27617 | n27618 ;
  assign n27620 = n21799 | n27619 ;
  assign n36501 = ~n27620 ;
  assign n27621 = x26 & n36501 ;
  assign n27622 = n30019 & n27620 ;
  assign n27623 = n27621 | n27622 ;
  assign n36502 = ~n27623 ;
  assign n27624 = n27616 & n36502 ;
  assign n36503 = ~n27616 ;
  assign n27625 = n36503 & n27623 ;
  assign n27626 = n27624 | n27625 ;
  assign n27627 = n27446 | n27453 ;
  assign n36504 = ~n27464 ;
  assign n27628 = n36504 & n27627 ;
  assign n27629 = n27626 & n27628 ;
  assign n27630 = n27626 | n27628 ;
  assign n36505 = ~n27629 ;
  assign n27631 = n36505 & n27630 ;
  assign n27632 = n27466 | n27468 ;
  assign n36506 = ~n27479 ;
  assign n27633 = n36506 & n27632 ;
  assign n27634 = n27631 & n27633 ;
  assign n27635 = n27631 | n27633 ;
  assign n36507 = ~n27634 ;
  assign n27636 = n36507 & n27635 ;
  assign n22573 = n4135 & n35022 ;
  assign n22554 = n4185 & n35018 ;
  assign n22595 = n4148 & n22533 ;
  assign n27637 = n22554 | n22595 ;
  assign n27638 = n4165 & n35020 ;
  assign n27639 = n27637 | n27638 ;
  assign n27640 = n22573 | n27639 ;
  assign n36508 = ~n27640 ;
  assign n27641 = x23 & n36508 ;
  assign n27642 = n30030 & n27640 ;
  assign n27643 = n27641 | n27642 ;
  assign n36509 = ~n27643 ;
  assign n27644 = n27636 & n36509 ;
  assign n36510 = ~n27636 ;
  assign n27645 = n36510 & n27643 ;
  assign n27646 = n27644 | n27645 ;
  assign n27647 = n27481 | n27483 ;
  assign n36511 = ~n27494 ;
  assign n27648 = n36511 & n27647 ;
  assign n23380 = n4686 & n23372 ;
  assign n23331 = n4706 & n35244 ;
  assign n23358 = n4726 & n23339 ;
  assign n27649 = n23331 | n23358 ;
  assign n27650 = n4748 & n35246 ;
  assign n27651 = n27649 | n27650 ;
  assign n27652 = n23380 | n27651 ;
  assign n36512 = ~n27652 ;
  assign n27653 = x20 & n36512 ;
  assign n27654 = n30374 & n27652 ;
  assign n27655 = n27653 | n27654 ;
  assign n27656 = n27648 | n27655 ;
  assign n27657 = n27648 & n27655 ;
  assign n36513 = ~n27657 ;
  assign n27658 = n27656 & n36513 ;
  assign n27659 = n27646 & n27658 ;
  assign n27660 = n27646 | n27658 ;
  assign n36514 = ~n27659 ;
  assign n27661 = n36514 & n27660 ;
  assign n36515 = ~n27508 ;
  assign n27662 = n27498 & n36515 ;
  assign n27663 = n27661 & n27662 ;
  assign n27664 = n27661 | n27662 ;
  assign n36516 = ~n27663 ;
  assign n27665 = n36516 & n27664 ;
  assign n27666 = n27572 & n27665 ;
  assign n27667 = n27572 | n27665 ;
  assign n36517 = ~n27666 ;
  assign n27668 = n36517 & n27667 ;
  assign n24880 = n5937 & n35662 ;
  assign n24677 = n5994 & n24676 ;
  assign n24841 = n5970 & n35663 ;
  assign n27669 = n24677 | n24841 ;
  assign n27670 = n6018 & n24815 ;
  assign n27671 = n27669 | n27670 ;
  assign n27672 = n24880 | n27671 ;
  assign n27673 = x14 | n27672 ;
  assign n27674 = x14 & n27672 ;
  assign n36518 = ~n27674 ;
  assign n27675 = n27673 & n36518 ;
  assign n27676 = n27668 & n27675 ;
  assign n27677 = n27668 | n27675 ;
  assign n36519 = ~n27676 ;
  assign n27678 = n36519 & n27677 ;
  assign n27679 = n27510 & n27517 ;
  assign n27680 = n27523 | n27679 ;
  assign n36520 = ~n27680 ;
  assign n27681 = n27678 & n36520 ;
  assign n36521 = ~n27678 ;
  assign n27682 = n36521 & n27680 ;
  assign n27683 = n27681 | n27682 ;
  assign n26072 = n6272 & n26065 ;
  assign n25400 = n6244 & n35784 ;
  assign n25799 = n6190 & n25796 ;
  assign n27684 = n25400 | n25799 ;
  assign n27685 = n6217 & n26039 ;
  assign n27686 = n27684 | n27685 ;
  assign n27687 = n26072 | n27686 ;
  assign n27688 = x11 | n27687 ;
  assign n27689 = x11 & n27687 ;
  assign n36522 = ~n27689 ;
  assign n27690 = n27688 & n36522 ;
  assign n27691 = n27683 & n27690 ;
  assign n27692 = n27683 | n27690 ;
  assign n36523 = ~n27691 ;
  assign n27693 = n36523 & n27692 ;
  assign n36524 = ~n27528 ;
  assign n27694 = n27527 & n36524 ;
  assign n36525 = ~n27694 ;
  assign n27695 = n27526 & n36525 ;
  assign n27696 = n27693 & n27695 ;
  assign n27697 = n27693 | n27695 ;
  assign n36526 = ~n27696 ;
  assign n27698 = n36526 & n27697 ;
  assign n26698 = n7068 & n36192 ;
  assign n27699 = n7041 & n26278 ;
  assign n27700 = n69 & n36131 ;
  assign n27701 = n27699 | n27700 ;
  assign n27702 = n26698 | n27701 ;
  assign n27703 = x8 | n27702 ;
  assign n27704 = x8 & n27702 ;
  assign n36527 = ~n27704 ;
  assign n27705 = n27703 & n36527 ;
  assign n36528 = ~n27698 ;
  assign n27706 = n36528 & n27705 ;
  assign n36529 = ~n27705 ;
  assign n27707 = n27698 & n36529 ;
  assign n27708 = n27706 | n27707 ;
  assign n36530 = ~n27544 ;
  assign n27709 = n27542 & n36530 ;
  assign n27710 = n27708 & n27709 ;
  assign n27711 = n27708 | n27709 ;
  assign n36531 = ~n27710 ;
  assign n27712 = n36531 & n27711 ;
  assign n27713 = n27546 & n27552 ;
  assign n27714 = n27551 | n27713 ;
  assign n27715 = n27712 | n27714 ;
  assign n27716 = n27712 & n27714 ;
  assign n36532 = ~n27716 ;
  assign n27717 = n27715 & n36532 ;
  assign n36533 = ~n27561 ;
  assign n27718 = n27558 & n36533 ;
  assign n36534 = ~n27717 ;
  assign n27719 = n36534 & n27718 ;
  assign n36535 = ~n27718 ;
  assign n27720 = n27717 & n36535 ;
  assign n27721 = n27719 | n27720 ;
  assign n27722 = n27565 | n27721 ;
  assign n27723 = n27565 & n27721 ;
  assign n36536 = ~n27723 ;
  assign n43 = n27722 & n36536 ;
  assign n27724 = n30223 & n27588 ;
  assign n36537 = ~n27724 ;
  assign n27725 = n3479 & n36537 ;
  assign n27726 = n1109 | n1210 ;
  assign n27727 = n5073 | n27726 ;
  assign n27728 = n4298 | n27727 ;
  assign n27729 = n5610 | n27728 ;
  assign n27730 = n510 | n946 ;
  assign n27731 = n988 | n27730 ;
  assign n27732 = n3682 | n15458 ;
  assign n27733 = n27731 | n27732 ;
  assign n27734 = n4633 | n27733 ;
  assign n27735 = n27729 | n27734 ;
  assign n27736 = n4049 | n13714 ;
  assign n27737 = n25871 | n27736 ;
  assign n27738 = n181 | n353 ;
  assign n27739 = n765 | n27738 ;
  assign n27740 = n291 | n27739 ;
  assign n27741 = n5528 | n27740 ;
  assign n27742 = n1635 | n1766 ;
  assign n27743 = n2203 | n12816 ;
  assign n27744 = n27742 | n27743 ;
  assign n27745 = n2453 | n27744 ;
  assign n27746 = n27741 | n27745 ;
  assign n27747 = n27737 | n27746 ;
  assign n27748 = n1316 | n27747 ;
  assign n27749 = n27735 | n27748 ;
  assign n27750 = n3978 | n27749 ;
  assign n27751 = n27725 | n27750 ;
  assign n27752 = n27725 & n27750 ;
  assign n36538 = ~n27752 ;
  assign n27753 = n27751 & n36538 ;
  assign n21100 = n889 & n34603 ;
  assign n19750 = n3329 & n34520 ;
  assign n19773 = n3311 & n19752 ;
  assign n27754 = n19750 | n19773 ;
  assign n27755 = n3343 & n34596 ;
  assign n27756 = n27754 | n27755 ;
  assign n27757 = n21100 | n27756 ;
  assign n36539 = ~n27757 ;
  assign n27758 = n27753 & n36539 ;
  assign n36540 = ~n27753 ;
  assign n27759 = n36540 & n27757 ;
  assign n27760 = n27758 | n27759 ;
  assign n27761 = n27594 & n27598 ;
  assign n27762 = n27592 | n27761 ;
  assign n27763 = n27760 | n27762 ;
  assign n27764 = n27760 & n27762 ;
  assign n36541 = ~n27764 ;
  assign n27765 = n27763 & n36541 ;
  assign n21881 = n895 & n34817 ;
  assign n19680 = n2849 & n34360 ;
  assign n19694 = n2861 & n34349 ;
  assign n27766 = n19680 | n19694 ;
  assign n27767 = n894 & n34803 ;
  assign n27768 = n27766 | n27767 ;
  assign n27769 = n21881 | n27768 ;
  assign n36542 = ~n27769 ;
  assign n27770 = x29 & n36542 ;
  assign n27771 = n30024 & n27769 ;
  assign n27772 = n27770 | n27771 ;
  assign n36543 = ~n27772 ;
  assign n27773 = n27765 & n36543 ;
  assign n36544 = ~n27765 ;
  assign n27774 = n36544 & n27772 ;
  assign n27775 = n27773 | n27774 ;
  assign n27776 = n27601 & n27608 ;
  assign n27777 = n27614 | n27776 ;
  assign n27778 = n27775 | n27777 ;
  assign n27779 = n27775 & n27777 ;
  assign n36545 = ~n27779 ;
  assign n27780 = n27778 & n36545 ;
  assign n22652 = n3791 & n35035 ;
  assign n21748 = n3802 & n21729 ;
  assign n21823 = n209 & n21753 ;
  assign n27781 = n21748 | n21823 ;
  assign n27782 = n3818 & n35018 ;
  assign n27783 = n27781 | n27782 ;
  assign n27784 = n22652 | n27783 ;
  assign n36546 = ~n27784 ;
  assign n27785 = x26 & n36546 ;
  assign n27786 = n30019 & n27784 ;
  assign n27787 = n27785 | n27786 ;
  assign n36547 = ~n27787 ;
  assign n27788 = n27780 & n36547 ;
  assign n36548 = ~n27780 ;
  assign n27789 = n36548 & n27787 ;
  assign n27790 = n27788 | n27789 ;
  assign n27791 = n27616 & n27623 ;
  assign n27792 = n27629 | n27791 ;
  assign n27793 = n27790 | n27792 ;
  assign n27794 = n27790 & n27792 ;
  assign n36549 = ~n27794 ;
  assign n27795 = n27793 & n36549 ;
  assign n23439 = n4135 & n35262 ;
  assign n22526 = n4148 & n35020 ;
  assign n22597 = n4185 & n22533 ;
  assign n27796 = n22526 | n22597 ;
  assign n27797 = n4165 & n23444 ;
  assign n27798 = n27796 | n27797 ;
  assign n27799 = n23439 | n27798 ;
  assign n36550 = ~n27799 ;
  assign n27800 = x23 & n36550 ;
  assign n27801 = n30030 & n27799 ;
  assign n27802 = n27800 | n27801 ;
  assign n36551 = ~n27802 ;
  assign n27803 = n27795 & n36551 ;
  assign n36552 = ~n27795 ;
  assign n27804 = n36552 & n27802 ;
  assign n27805 = n27803 | n27804 ;
  assign n27806 = n27636 & n27643 ;
  assign n27807 = n27634 | n27806 ;
  assign n27808 = n27805 | n27807 ;
  assign n27809 = n27805 & n27807 ;
  assign n36553 = ~n27809 ;
  assign n27810 = n27808 & n36553 ;
  assign n24203 = n4686 & n35472 ;
  assign n23296 = n4706 & n35467 ;
  assign n23332 = n4726 & n35244 ;
  assign n27811 = n23296 | n23332 ;
  assign n27812 = n4748 & n35465 ;
  assign n27813 = n27811 | n27812 ;
  assign n27814 = n24203 | n27813 ;
  assign n36554 = ~n27814 ;
  assign n27815 = x20 & n36554 ;
  assign n27816 = n30374 & n27814 ;
  assign n27817 = n27815 | n27816 ;
  assign n36555 = ~n27817 ;
  assign n27818 = n27810 & n36555 ;
  assign n36556 = ~n27810 ;
  assign n27819 = n36556 & n27817 ;
  assign n27820 = n27818 | n27819 ;
  assign n27821 = n27657 | n27659 ;
  assign n27822 = n27820 | n27821 ;
  assign n27823 = n27820 & n27821 ;
  assign n36557 = ~n27823 ;
  assign n27824 = n27822 & n36557 ;
  assign n25295 = n37300 & n25288 ;
  assign n24060 = n5144 & n24057 ;
  assign n24087 = n5166 & n24080 ;
  assign n27825 = n24060 | n24087 ;
  assign n27826 = n5191 & n24676 ;
  assign n27827 = n27825 | n27826 ;
  assign n27828 = n25295 | n27827 ;
  assign n36558 = ~n27828 ;
  assign n27829 = x17 & n36558 ;
  assign n27830 = n30580 & n27828 ;
  assign n27831 = n27829 | n27830 ;
  assign n36559 = ~n27831 ;
  assign n27832 = n27824 & n36559 ;
  assign n36560 = ~n27824 ;
  assign n27833 = n36560 & n27831 ;
  assign n27834 = n27832 | n27833 ;
  assign n27835 = n27663 | n27666 ;
  assign n36561 = ~n27835 ;
  assign n27836 = n27834 & n36561 ;
  assign n36562 = ~n27834 ;
  assign n27837 = n36562 & n27835 ;
  assign n27838 = n27836 | n27837 ;
  assign n25426 = n5937 & n35785 ;
  assign n24820 = n5970 & n24815 ;
  assign n24840 = n5994 & n35663 ;
  assign n27839 = n24820 | n24840 ;
  assign n27840 = n6018 & n35784 ;
  assign n27841 = n27839 | n27840 ;
  assign n27842 = n25426 | n27841 ;
  assign n36563 = ~n27842 ;
  assign n27843 = x14 & n36563 ;
  assign n27844 = n30547 & n27842 ;
  assign n27845 = n27843 | n27844 ;
  assign n36564 = ~n27845 ;
  assign n27846 = n27838 & n36564 ;
  assign n36565 = ~n27838 ;
  assign n27847 = n36565 & n27845 ;
  assign n27848 = n27846 | n27847 ;
  assign n26290 = n6272 & n26284 ;
  assign n25798 = n6244 & n25796 ;
  assign n26043 = n6190 & n26039 ;
  assign n27849 = n25798 | n26043 ;
  assign n27850 = n6217 & n26278 ;
  assign n27851 = n27849 | n27850 ;
  assign n27852 = n26290 | n27851 ;
  assign n27853 = x11 | n27852 ;
  assign n27854 = x11 & n27852 ;
  assign n36566 = ~n27854 ;
  assign n27855 = n27853 & n36566 ;
  assign n27856 = n27848 & n27855 ;
  assign n27857 = n27848 | n27855 ;
  assign n36567 = ~n27856 ;
  assign n27858 = n36567 & n27857 ;
  assign n27859 = n27678 & n27680 ;
  assign n27860 = n27676 | n27859 ;
  assign n36568 = ~n27860 ;
  assign n27861 = n27858 & n36568 ;
  assign n36569 = ~n27858 ;
  assign n27862 = n36569 & n27860 ;
  assign n27863 = n27861 | n27862 ;
  assign n27864 = n70 | n26279 ;
  assign n27865 = n30185 & n27864 ;
  assign n27866 = x7 | n27864 ;
  assign n36570 = ~n27865 ;
  assign n27867 = n36570 & n27866 ;
  assign n36571 = ~n27867 ;
  assign n27868 = n27863 & n36571 ;
  assign n36572 = ~n27863 ;
  assign n27869 = n36572 & n27867 ;
  assign n27870 = n27868 | n27869 ;
  assign n36573 = ~n27695 ;
  assign n27871 = n27693 & n36573 ;
  assign n36574 = ~n27871 ;
  assign n27872 = n27692 & n36574 ;
  assign n27873 = n27870 & n27872 ;
  assign n27874 = n27870 | n27872 ;
  assign n36575 = ~n27873 ;
  assign n27875 = n36575 & n27874 ;
  assign n27876 = n27698 | n27705 ;
  assign n36576 = ~n27709 ;
  assign n27877 = n27708 & n36576 ;
  assign n36577 = ~n27877 ;
  assign n27878 = n27876 & n36577 ;
  assign n27879 = n27875 & n27878 ;
  assign n27880 = n27875 | n27878 ;
  assign n36578 = ~n27879 ;
  assign n27881 = n36578 & n27880 ;
  assign n36579 = ~n27720 ;
  assign n27882 = n27715 & n36579 ;
  assign n27883 = n27881 | n27882 ;
  assign n27885 = n27881 & n27882 ;
  assign n36580 = ~n27885 ;
  assign n27886 = n27883 & n36580 ;
  assign n27887 = n27723 | n27886 ;
  assign n27888 = n27723 & n27886 ;
  assign n36581 = ~n27888 ;
  assign n44 = n27887 & n36581 ;
  assign n27889 = n27858 & n27860 ;
  assign n27890 = n27856 | n27889 ;
  assign n27891 = x8 | n27890 ;
  assign n27892 = x8 & n27890 ;
  assign n36582 = ~n27892 ;
  assign n27893 = n27891 & n36582 ;
  assign n27894 = n160 | n354 ;
  assign n27895 = n833 | n846 ;
  assign n27896 = n27894 | n27895 ;
  assign n27897 = n3852 | n11127 ;
  assign n27898 = n27896 | n27897 ;
  assign n27899 = n2746 | n4618 ;
  assign n27900 = n13255 | n13434 ;
  assign n27901 = n27899 | n27900 ;
  assign n27902 = n3689 | n27901 ;
  assign n27903 = n27898 | n27902 ;
  assign n36583 = ~n27903 ;
  assign n27904 = n2309 & n36583 ;
  assign n27905 = n194 | n401 ;
  assign n27906 = n480 | n540 ;
  assign n27907 = n27905 | n27906 ;
  assign n27908 = n384 | n3099 ;
  assign n27909 = n27907 | n27908 ;
  assign n27910 = n5371 | n27909 ;
  assign n27911 = n22986 | n27910 ;
  assign n27912 = n418 | n489 ;
  assign n27913 = n713 | n27912 ;
  assign n27914 = n269 | n279 ;
  assign n27915 = n3240 | n27914 ;
  assign n27916 = n13501 | n27915 ;
  assign n27917 = n27913 | n27916 ;
  assign n27918 = n12800 | n27917 ;
  assign n27919 = n27911 | n27918 ;
  assign n27920 = n13891 | n27919 ;
  assign n36584 = ~n27920 ;
  assign n27921 = n27904 & n36584 ;
  assign n36585 = ~n21508 ;
  assign n27922 = n36585 & n27921 ;
  assign n36586 = ~n27750 ;
  assign n27923 = n36586 & n27922 ;
  assign n36587 = ~n27922 ;
  assign n27924 = n27750 & n36587 ;
  assign n27925 = n27923 | n27924 ;
  assign n27926 = n27752 | n27758 ;
  assign n36588 = ~n27926 ;
  assign n27927 = n27925 & n36588 ;
  assign n36589 = ~n27925 ;
  assign n27928 = n36589 & n27926 ;
  assign n27929 = n27927 | n27928 ;
  assign n21080 = n889 & n34598 ;
  assign n19722 = n3329 & n34363 ;
  assign n19737 = n3311 & n34520 ;
  assign n27930 = n19722 | n19737 ;
  assign n27931 = n3343 & n34349 ;
  assign n27932 = n27930 | n27931 ;
  assign n27933 = n21080 | n27932 ;
  assign n36590 = ~n27933 ;
  assign n27934 = n27929 & n36590 ;
  assign n36591 = ~n27929 ;
  assign n27935 = n36591 & n27933 ;
  assign n27936 = n27934 | n27935 ;
  assign n36592 = ~n27773 ;
  assign n27937 = n27763 & n36592 ;
  assign n36593 = ~n27936 ;
  assign n27938 = n36593 & n27937 ;
  assign n36594 = ~n27937 ;
  assign n27939 = n27936 & n36594 ;
  assign n27940 = n27938 | n27939 ;
  assign n21858 = n895 & n21848 ;
  assign n19673 = n2861 & n34360 ;
  assign n21774 = n2849 & n34803 ;
  assign n27941 = n19673 | n21774 ;
  assign n27942 = n894 & n21753 ;
  assign n27943 = n27941 | n27942 ;
  assign n27944 = n21858 | n27943 ;
  assign n27945 = x29 | n27944 ;
  assign n27946 = x29 & n27944 ;
  assign n36595 = ~n27946 ;
  assign n27947 = n27945 & n36595 ;
  assign n27948 = n27940 & n27947 ;
  assign n27949 = n27940 | n27947 ;
  assign n36596 = ~n27948 ;
  assign n27950 = n36596 & n27949 ;
  assign n22630 = n3791 & n35030 ;
  assign n21749 = n209 & n21729 ;
  assign n22555 = n3802 & n35018 ;
  assign n27951 = n21749 | n22555 ;
  assign n27952 = n3818 & n22533 ;
  assign n27953 = n27951 | n27952 ;
  assign n27954 = n22630 | n27953 ;
  assign n36597 = ~n27954 ;
  assign n27955 = x26 & n36597 ;
  assign n27956 = n30019 & n27954 ;
  assign n27957 = n27955 | n27956 ;
  assign n36598 = ~n27957 ;
  assign n27958 = n27950 & n36598 ;
  assign n36599 = ~n27950 ;
  assign n27959 = n36599 & n27957 ;
  assign n27960 = n27958 | n27959 ;
  assign n36600 = ~n27788 ;
  assign n27961 = n27778 & n36600 ;
  assign n36601 = ~n27960 ;
  assign n27962 = n36601 & n27961 ;
  assign n36602 = ~n27961 ;
  assign n27963 = n27960 & n36602 ;
  assign n27964 = n27962 | n27963 ;
  assign n23412 = n4135 & n35252 ;
  assign n22528 = n4185 & n35020 ;
  assign n23359 = n4148 & n23339 ;
  assign n27965 = n22528 | n23359 ;
  assign n27966 = n4165 & n35254 ;
  assign n27967 = n27965 | n27966 ;
  assign n27968 = n23412 | n27967 ;
  assign n36603 = ~n27968 ;
  assign n27969 = x23 & n36603 ;
  assign n27970 = n30030 & n27968 ;
  assign n27971 = n27969 | n27970 ;
  assign n27972 = n27964 | n27971 ;
  assign n27973 = n27964 & n27971 ;
  assign n36604 = ~n27973 ;
  assign n27974 = n27972 & n36604 ;
  assign n36605 = ~n27803 ;
  assign n27975 = n27793 & n36605 ;
  assign n36606 = ~n27974 ;
  assign n27976 = n36606 & n27975 ;
  assign n36607 = ~n27975 ;
  assign n27977 = n27974 & n36607 ;
  assign n27978 = n27976 | n27977 ;
  assign n24175 = n4686 & n24168 ;
  assign n23302 = n4726 & n35467 ;
  assign n24115 = n4706 & n35458 ;
  assign n27979 = n23302 | n24115 ;
  assign n27980 = n4748 & n24080 ;
  assign n27981 = n27979 | n27980 ;
  assign n27982 = n24175 | n27981 ;
  assign n36608 = ~n27982 ;
  assign n27983 = x20 & n36608 ;
  assign n27984 = n30374 & n27982 ;
  assign n27985 = n27983 | n27984 ;
  assign n27986 = n27978 | n27985 ;
  assign n27987 = n27978 & n27985 ;
  assign n36609 = ~n27987 ;
  assign n27988 = n27986 & n36609 ;
  assign n36610 = ~n27818 ;
  assign n27989 = n27808 & n36610 ;
  assign n27990 = n27988 & n27989 ;
  assign n27991 = n27988 | n27989 ;
  assign n36611 = ~n27990 ;
  assign n27992 = n36611 & n27991 ;
  assign n25325 = n37300 & n35670 ;
  assign n24058 = n5166 & n24057 ;
  assign n24687 = n5144 & n24676 ;
  assign n27993 = n24058 | n24687 ;
  assign n27994 = n5191 & n35663 ;
  assign n27995 = n27993 | n27994 ;
  assign n27996 = n25325 | n27995 ;
  assign n36612 = ~n27996 ;
  assign n27997 = x17 & n36612 ;
  assign n27998 = n30580 & n27996 ;
  assign n27999 = n27997 | n27998 ;
  assign n28000 = n27992 | n27999 ;
  assign n28001 = n27992 & n27999 ;
  assign n36613 = ~n28001 ;
  assign n28002 = n28000 & n36613 ;
  assign n36614 = ~n27832 ;
  assign n28003 = n27822 & n36614 ;
  assign n28004 = n28002 & n28003 ;
  assign n28005 = n28002 | n28003 ;
  assign n36615 = ~n28004 ;
  assign n28006 = n36615 & n28005 ;
  assign n25828 = n5937 & n35910 ;
  assign n24817 = n5994 & n24815 ;
  assign n25398 = n5970 & n35784 ;
  assign n28007 = n24817 | n25398 ;
  assign n28008 = n6018 & n25796 ;
  assign n28009 = n28007 | n28008 ;
  assign n28010 = n25828 | n28009 ;
  assign n36616 = ~n28010 ;
  assign n28011 = x14 & n36616 ;
  assign n28012 = n30547 & n28010 ;
  assign n28013 = n28011 | n28012 ;
  assign n28014 = n28006 | n28013 ;
  assign n28015 = n28006 & n28013 ;
  assign n36617 = ~n28015 ;
  assign n28016 = n28014 & n36617 ;
  assign n26490 = n6272 & n36130 ;
  assign n26041 = n6244 & n26039 ;
  assign n26477 = n6190 & n26278 ;
  assign n28017 = n26041 | n26477 ;
  assign n28018 = n6217 & n36131 ;
  assign n28019 = n28017 | n28018 ;
  assign n28020 = n26490 | n28019 ;
  assign n28021 = x11 | n28020 ;
  assign n28022 = x11 & n28020 ;
  assign n36618 = ~n28022 ;
  assign n28023 = n28021 & n36618 ;
  assign n28024 = n27834 & n27835 ;
  assign n28025 = n27838 & n27845 ;
  assign n28026 = n28024 | n28025 ;
  assign n36619 = ~n28026 ;
  assign n28027 = n28023 & n36619 ;
  assign n36620 = ~n28023 ;
  assign n28028 = n36620 & n28026 ;
  assign n28029 = n28027 | n28028 ;
  assign n36621 = ~n28016 ;
  assign n28030 = n36621 & n28029 ;
  assign n36622 = ~n28029 ;
  assign n28031 = n28016 & n36622 ;
  assign n28032 = n28030 | n28031 ;
  assign n36623 = ~n28032 ;
  assign n28033 = n27893 & n36623 ;
  assign n36624 = ~n27893 ;
  assign n28034 = n36624 & n28032 ;
  assign n28035 = n28033 | n28034 ;
  assign n28036 = n27863 & n27867 ;
  assign n28037 = n27873 | n28036 ;
  assign n36625 = ~n28037 ;
  assign n28038 = n28035 & n36625 ;
  assign n36626 = ~n28035 ;
  assign n28039 = n36626 & n28037 ;
  assign n28040 = n28038 | n28039 ;
  assign n36627 = ~n27882 ;
  assign n27884 = n27881 & n36627 ;
  assign n36628 = ~n27884 ;
  assign n28041 = n27880 & n36628 ;
  assign n28042 = n28040 & n28041 ;
  assign n28043 = n28040 | n28041 ;
  assign n36629 = ~n28042 ;
  assign n28044 = n36629 & n28043 ;
  assign n28045 = n36581 & n28044 ;
  assign n36630 = ~n28044 ;
  assign n28046 = n27888 & n36630 ;
  assign n29895 = n28045 | n28046 ;
  assign n28047 = n658 | n688 ;
  assign n28048 = n1825 | n2748 ;
  assign n28049 = n28047 | n28048 ;
  assign n28050 = n955 | n22204 ;
  assign n28051 = n28049 | n28050 ;
  assign n28052 = n1319 | n1412 ;
  assign n28053 = n4625 | n22183 ;
  assign n28054 = n28052 | n28053 ;
  assign n28055 = n28051 | n28054 ;
  assign n28056 = n1905 | n28055 ;
  assign n28057 = n4563 | n28056 ;
  assign n36631 = ~n28057 ;
  assign n28058 = n2402 & n36631 ;
  assign n28059 = n36586 & n28058 ;
  assign n36632 = ~n28058 ;
  assign n28060 = n27750 & n36632 ;
  assign n28061 = n28059 | n28060 ;
  assign n28062 = x8 | n28061 ;
  assign n28063 = x8 & n28061 ;
  assign n36633 = ~n28063 ;
  assign n28064 = n28062 & n36633 ;
  assign n20158 = n889 & n34362 ;
  assign n19692 = n3329 & n34349 ;
  assign n19710 = n3311 & n34363 ;
  assign n28065 = n19692 | n19710 ;
  assign n28066 = n3343 & n34365 ;
  assign n28067 = n28065 | n28066 ;
  assign n28068 = n20158 | n28067 ;
  assign n28069 = n28064 | n28068 ;
  assign n28070 = n28064 & n28068 ;
  assign n36634 = ~n28070 ;
  assign n28071 = n28069 & n36634 ;
  assign n28072 = n27750 & n27922 ;
  assign n28073 = n27925 & n27926 ;
  assign n28074 = n28072 | n28073 ;
  assign n36635 = ~n28074 ;
  assign n28075 = n28071 & n36635 ;
  assign n36636 = ~n28071 ;
  assign n28076 = n36636 & n28074 ;
  assign n28077 = n28075 | n28076 ;
  assign n21800 = n895 & n34802 ;
  assign n21775 = n2861 & n34803 ;
  assign n21824 = n2849 & n21753 ;
  assign n28078 = n21775 | n21824 ;
  assign n28079 = n894 & n21804 ;
  assign n28080 = n28078 | n28079 ;
  assign n28081 = n21800 | n28080 ;
  assign n36637 = ~n28081 ;
  assign n28082 = x29 & n36637 ;
  assign n28083 = n30024 & n28081 ;
  assign n28084 = n28082 | n28083 ;
  assign n36638 = ~n28084 ;
  assign n28085 = n28077 & n36638 ;
  assign n36639 = ~n28077 ;
  assign n28086 = n36639 & n28084 ;
  assign n28087 = n28085 | n28086 ;
  assign n28088 = n27936 | n27937 ;
  assign n36640 = ~n27934 ;
  assign n28089 = n36640 & n28088 ;
  assign n36641 = ~n28087 ;
  assign n28090 = n36641 & n28089 ;
  assign n36642 = ~n28089 ;
  assign n28091 = n28087 & n36642 ;
  assign n28092 = n28090 | n28091 ;
  assign n22574 = n3791 & n35022 ;
  assign n22550 = n209 & n35018 ;
  assign n22579 = n3802 & n22533 ;
  assign n28093 = n22550 | n22579 ;
  assign n28094 = n3818 & n35020 ;
  assign n28095 = n28093 | n28094 ;
  assign n28096 = n22574 | n28095 ;
  assign n36643 = ~n28096 ;
  assign n28097 = x26 & n36643 ;
  assign n28098 = n30019 & n28096 ;
  assign n28099 = n28097 | n28098 ;
  assign n36644 = ~n28099 ;
  assign n28100 = n28092 & n36644 ;
  assign n36645 = ~n28092 ;
  assign n28101 = n36645 & n28099 ;
  assign n28102 = n28100 | n28101 ;
  assign n36646 = ~n27947 ;
  assign n28103 = n27940 & n36646 ;
  assign n28104 = n27950 | n27957 ;
  assign n36647 = ~n28103 ;
  assign n28105 = n36647 & n28104 ;
  assign n36648 = ~n28102 ;
  assign n28106 = n36648 & n28105 ;
  assign n36649 = ~n28105 ;
  assign n28107 = n28102 & n36649 ;
  assign n28108 = n28106 | n28107 ;
  assign n36650 = ~n27964 ;
  assign n28109 = n36650 & n27971 ;
  assign n28110 = n27962 | n28109 ;
  assign n23381 = n4135 & n23372 ;
  assign n23333 = n4148 & n35244 ;
  assign n23360 = n4185 & n23339 ;
  assign n28111 = n23333 | n23360 ;
  assign n28112 = n4165 & n35246 ;
  assign n28113 = n28111 | n28112 ;
  assign n28114 = n23381 | n28113 ;
  assign n36651 = ~n28114 ;
  assign n28115 = x23 & n36651 ;
  assign n28116 = n30030 & n28114 ;
  assign n28117 = n28115 | n28116 ;
  assign n28118 = n28110 | n28117 ;
  assign n28119 = n28110 & n28117 ;
  assign n36652 = ~n28119 ;
  assign n28120 = n28118 & n36652 ;
  assign n28121 = n28108 & n28120 ;
  assign n28122 = n28108 | n28120 ;
  assign n36653 = ~n28121 ;
  assign n28123 = n36653 & n28122 ;
  assign n24146 = n4686 & n35457 ;
  assign n24095 = n4706 & n24080 ;
  assign n24122 = n4726 & n35458 ;
  assign n28124 = n24095 | n24122 ;
  assign n28125 = n4748 & n24151 ;
  assign n28126 = n28124 | n28125 ;
  assign n28127 = n24146 | n28126 ;
  assign n28128 = x20 | n28127 ;
  assign n28129 = x20 & n28127 ;
  assign n36654 = ~n28129 ;
  assign n28130 = n28128 & n36654 ;
  assign n36655 = ~n27977 ;
  assign n28131 = n36655 & n27986 ;
  assign n28132 = n28130 & n28131 ;
  assign n28133 = n28130 | n28131 ;
  assign n36656 = ~n28132 ;
  assign n28134 = n36656 & n28133 ;
  assign n28135 = n28123 & n28134 ;
  assign n28136 = n28123 | n28134 ;
  assign n36657 = ~n28135 ;
  assign n28137 = n36657 & n28136 ;
  assign n24881 = n37300 & n35662 ;
  assign n24689 = n5166 & n24676 ;
  assign n24839 = n5144 & n35663 ;
  assign n28138 = n24689 | n24839 ;
  assign n28139 = n5191 & n24815 ;
  assign n28140 = n28138 | n28139 ;
  assign n28141 = n24881 | n28140 ;
  assign n36658 = ~n28141 ;
  assign n28142 = x17 & n36658 ;
  assign n28143 = n30580 & n28141 ;
  assign n28144 = n28142 | n28143 ;
  assign n28145 = n28137 | n28144 ;
  assign n28146 = n28137 & n28144 ;
  assign n36659 = ~n28146 ;
  assign n28147 = n28145 & n36659 ;
  assign n36660 = ~n27989 ;
  assign n28148 = n27988 & n36660 ;
  assign n36661 = ~n28148 ;
  assign n28149 = n28000 & n36661 ;
  assign n36662 = ~n28147 ;
  assign n28150 = n36662 & n28149 ;
  assign n36663 = ~n28149 ;
  assign n28151 = n28147 & n36663 ;
  assign n28152 = n28150 | n28151 ;
  assign n26071 = n5937 & n26065 ;
  assign n25404 = n5994 & n35784 ;
  assign n25797 = n5970 & n25796 ;
  assign n28153 = n25404 | n25797 ;
  assign n28154 = n6018 & n26039 ;
  assign n28155 = n28153 | n28154 ;
  assign n28156 = n26071 | n28155 ;
  assign n28157 = x14 | n28156 ;
  assign n28158 = x14 & n28156 ;
  assign n36664 = ~n28158 ;
  assign n28159 = n28157 & n36664 ;
  assign n36665 = ~n28003 ;
  assign n28160 = n28002 & n36665 ;
  assign n36666 = ~n28160 ;
  assign n28161 = n28014 & n36666 ;
  assign n28162 = n28159 & n28161 ;
  assign n28163 = n28159 | n28161 ;
  assign n36667 = ~n28162 ;
  assign n28164 = n36667 & n28163 ;
  assign n28165 = n28152 & n28164 ;
  assign n28166 = n28152 | n28164 ;
  assign n36668 = ~n28165 ;
  assign n28167 = n36668 & n28166 ;
  assign n26699 = n6272 & n36192 ;
  assign n28168 = n6244 & n26278 ;
  assign n28169 = n6190 & n36131 ;
  assign n28170 = n28168 | n28169 ;
  assign n28171 = n26699 | n28170 ;
  assign n28172 = x11 | n28171 ;
  assign n28173 = x11 & n28171 ;
  assign n36669 = ~n28173 ;
  assign n28174 = n28172 & n36669 ;
  assign n28175 = n28023 & n28026 ;
  assign n28176 = n28030 | n28175 ;
  assign n36670 = ~n28176 ;
  assign n28177 = n28174 & n36670 ;
  assign n36671 = ~n28174 ;
  assign n28178 = n36671 & n28176 ;
  assign n28179 = n28177 | n28178 ;
  assign n28180 = n28167 & n28179 ;
  assign n28182 = n28167 | n28179 ;
  assign n36672 = ~n28180 ;
  assign n28183 = n36672 & n28182 ;
  assign n28184 = n27893 & n28032 ;
  assign n36673 = ~n28184 ;
  assign n28185 = n27891 & n36673 ;
  assign n36674 = ~n28183 ;
  assign n28186 = n36674 & n28185 ;
  assign n36675 = ~n28185 ;
  assign n28187 = n28183 & n36675 ;
  assign n28188 = n28186 | n28187 ;
  assign n36676 = ~n26692 ;
  assign n28189 = n36676 & n26710 ;
  assign n28190 = n26878 | n28189 ;
  assign n28191 = n26875 | n28190 ;
  assign n28192 = n36318 & n28191 ;
  assign n36677 = ~n27054 ;
  assign n28193 = n36677 & n28192 ;
  assign n28194 = n27223 | n28193 ;
  assign n36678 = ~n27220 ;
  assign n28195 = n36678 & n28194 ;
  assign n28196 = n27218 | n28195 ;
  assign n28197 = n27392 | n28196 ;
  assign n28198 = n27393 & n28197 ;
  assign n28199 = n27559 | n28198 ;
  assign n28200 = n27558 & n28199 ;
  assign n28201 = n27716 | n28200 ;
  assign n28202 = n27715 & n28201 ;
  assign n36679 = ~n28202 ;
  assign n28203 = n27881 & n36679 ;
  assign n36680 = ~n28203 ;
  assign n28204 = n27880 & n36680 ;
  assign n28205 = n28040 | n28204 ;
  assign n36681 = ~n28038 ;
  assign n28206 = n36681 & n28205 ;
  assign n28207 = n28188 & n28206 ;
  assign n28208 = n28188 | n28206 ;
  assign n36682 = ~n28207 ;
  assign n28209 = n36682 & n28208 ;
  assign n36683 = ~n28046 ;
  assign n28210 = n36683 & n28209 ;
  assign n36684 = ~n28209 ;
  assign n28211 = n28046 & n36684 ;
  assign n29894 = n28210 | n28211 ;
  assign n36685 = ~n28060 ;
  assign n28212 = n36685 & n28062 ;
  assign n28213 = n602 | n2606 ;
  assign n28214 = n4255 | n11658 ;
  assign n28215 = n28213 | n28214 ;
  assign n28216 = n490 | n687 ;
  assign n28217 = n1355 | n28216 ;
  assign n28218 = n2407 | n13402 ;
  assign n28219 = n28217 | n28218 ;
  assign n28220 = n28215 | n28219 ;
  assign n28221 = n11207 | n21358 ;
  assign n28222 = n28220 | n28221 ;
  assign n28223 = n4809 | n28222 ;
  assign n36686 = ~n28223 ;
  assign n28224 = n1613 & n36686 ;
  assign n28225 = n28212 | n28224 ;
  assign n28226 = n28212 & n28224 ;
  assign n36687 = ~n28226 ;
  assign n28227 = n28225 & n36687 ;
  assign n21882 = n889 & n34817 ;
  assign n19663 = n3329 & n34360 ;
  assign n19703 = n3311 & n34349 ;
  assign n28228 = n19663 | n19703 ;
  assign n28229 = n3343 & n34803 ;
  assign n28230 = n28228 | n28229 ;
  assign n28231 = n21882 | n28230 ;
  assign n28232 = n28227 | n28231 ;
  assign n28233 = n28227 & n28231 ;
  assign n36688 = ~n28233 ;
  assign n28234 = n28232 & n36688 ;
  assign n28235 = n28071 & n28074 ;
  assign n36689 = ~n28235 ;
  assign n28236 = n28069 & n36689 ;
  assign n36690 = ~n28234 ;
  assign n28237 = n36690 & n28236 ;
  assign n36691 = ~n28236 ;
  assign n28238 = n28234 & n36691 ;
  assign n28239 = n28237 | n28238 ;
  assign n22653 = n895 & n35035 ;
  assign n21746 = n2849 & n21729 ;
  assign n21825 = n2861 & n21753 ;
  assign n28240 = n21746 | n21825 ;
  assign n28241 = n894 & n35018 ;
  assign n28242 = n28240 | n28241 ;
  assign n28243 = n22653 | n28242 ;
  assign n36692 = ~n28243 ;
  assign n28244 = x29 & n36692 ;
  assign n28245 = n30024 & n28243 ;
  assign n28246 = n28244 | n28245 ;
  assign n28247 = n28239 | n28246 ;
  assign n28248 = n28239 & n28246 ;
  assign n36693 = ~n28248 ;
  assign n28249 = n28247 & n36693 ;
  assign n28250 = n28087 | n28089 ;
  assign n36694 = ~n28085 ;
  assign n28251 = n36694 & n28250 ;
  assign n36695 = ~n28249 ;
  assign n28252 = n36695 & n28251 ;
  assign n36696 = ~n28251 ;
  assign n28253 = n28249 & n36696 ;
  assign n28254 = n28252 | n28253 ;
  assign n23435 = n3791 & n35262 ;
  assign n22520 = n3802 & n35020 ;
  assign n22598 = n209 & n22533 ;
  assign n28255 = n22520 | n22598 ;
  assign n28256 = n3818 & n23444 ;
  assign n28257 = n28255 | n28256 ;
  assign n28258 = n23435 | n28257 ;
  assign n36697 = ~n28258 ;
  assign n28259 = x26 & n36697 ;
  assign n28260 = n30019 & n28258 ;
  assign n28261 = n28259 | n28260 ;
  assign n28262 = n28254 | n28261 ;
  assign n28263 = n28254 & n28261 ;
  assign n36698 = ~n28263 ;
  assign n28264 = n28262 & n36698 ;
  assign n28265 = n28102 | n28105 ;
  assign n36699 = ~n28100 ;
  assign n28266 = n36699 & n28265 ;
  assign n28267 = n28264 & n28266 ;
  assign n28268 = n28264 | n28266 ;
  assign n36700 = ~n28267 ;
  assign n28269 = n36700 & n28268 ;
  assign n24201 = n4135 & n35472 ;
  assign n23308 = n4148 & n35467 ;
  assign n23334 = n4185 & n35244 ;
  assign n28270 = n23308 | n23334 ;
  assign n28271 = n4165 & n35465 ;
  assign n28272 = n28270 | n28271 ;
  assign n28273 = n24201 | n28272 ;
  assign n36701 = ~n28273 ;
  assign n28274 = x23 & n36701 ;
  assign n28275 = n30030 & n28273 ;
  assign n28276 = n28274 | n28275 ;
  assign n28277 = n28269 | n28276 ;
  assign n28278 = n28269 & n28276 ;
  assign n36702 = ~n28278 ;
  assign n28279 = n28277 & n36702 ;
  assign n28280 = n28118 & n36653 ;
  assign n28281 = n28279 & n28280 ;
  assign n28282 = n28279 | n28280 ;
  assign n36703 = ~n28281 ;
  assign n28283 = n36703 & n28282 ;
  assign n25294 = n4686 & n25288 ;
  assign n24070 = n4706 & n24057 ;
  assign n24082 = n4726 & n24080 ;
  assign n28284 = n24070 | n24082 ;
  assign n28285 = n4748 & n24676 ;
  assign n28286 = n28284 | n28285 ;
  assign n28287 = n25294 | n28286 ;
  assign n36704 = ~n28287 ;
  assign n28288 = x20 & n36704 ;
  assign n28289 = n30374 & n28287 ;
  assign n28290 = n28288 | n28289 ;
  assign n28291 = n28283 | n28290 ;
  assign n28292 = n28283 & n28290 ;
  assign n36705 = ~n28292 ;
  assign n28293 = n28291 & n36705 ;
  assign n36706 = ~n28123 ;
  assign n28294 = n36706 & n28134 ;
  assign n28295 = n28132 | n28294 ;
  assign n36707 = ~n28295 ;
  assign n28296 = n28293 & n36707 ;
  assign n36708 = ~n28293 ;
  assign n28297 = n36708 & n28295 ;
  assign n28298 = n28296 | n28297 ;
  assign n25427 = n37300 & n35785 ;
  assign n24824 = n5144 & n24815 ;
  assign n24846 = n5166 & n35663 ;
  assign n28299 = n24824 | n24846 ;
  assign n28300 = n5191 & n35784 ;
  assign n28301 = n28299 | n28300 ;
  assign n28302 = n25427 | n28301 ;
  assign n36709 = ~n28302 ;
  assign n28303 = x17 & n36709 ;
  assign n28304 = n30580 & n28302 ;
  assign n28305 = n28303 | n28304 ;
  assign n28306 = n28298 | n28305 ;
  assign n28307 = n28298 & n28305 ;
  assign n36710 = ~n28307 ;
  assign n28308 = n28306 & n36710 ;
  assign n36711 = ~n28137 ;
  assign n28309 = n36711 & n28144 ;
  assign n28310 = n28150 | n28309 ;
  assign n36712 = ~n28310 ;
  assign n28311 = n28308 & n36712 ;
  assign n36713 = ~n28308 ;
  assign n28312 = n36713 & n28310 ;
  assign n28313 = n28311 | n28312 ;
  assign n26292 = n5937 & n26284 ;
  assign n25806 = n5994 & n25796 ;
  assign n26053 = n5970 & n26039 ;
  assign n28314 = n25806 | n26053 ;
  assign n28315 = n6018 & n26278 ;
  assign n28316 = n28314 | n28315 ;
  assign n28317 = n26292 | n28316 ;
  assign n36714 = ~n28317 ;
  assign n28318 = x14 & n36714 ;
  assign n28319 = n30547 & n28317 ;
  assign n28320 = n28318 | n28319 ;
  assign n28321 = n28313 | n28320 ;
  assign n28322 = n28313 & n28320 ;
  assign n36715 = ~n28322 ;
  assign n28323 = n28321 & n36715 ;
  assign n28324 = n6213 | n26279 ;
  assign n28325 = n30180 & n28324 ;
  assign n28326 = x10 | n28324 ;
  assign n36716 = ~n28325 ;
  assign n28327 = n36716 & n28326 ;
  assign n28328 = n28163 & n36668 ;
  assign n36717 = ~n28327 ;
  assign n28329 = n36717 & n28328 ;
  assign n36718 = ~n28328 ;
  assign n28330 = n28327 & n36718 ;
  assign n28331 = n28329 | n28330 ;
  assign n28332 = n28323 & n28331 ;
  assign n28333 = n28323 | n28331 ;
  assign n36719 = ~n28332 ;
  assign n28334 = n36719 & n28333 ;
  assign n36720 = ~n28167 ;
  assign n28181 = n36720 & n28179 ;
  assign n28335 = n28174 & n28176 ;
  assign n28336 = n28181 | n28335 ;
  assign n36721 = ~n28336 ;
  assign n28337 = n28334 & n36721 ;
  assign n36722 = ~n28334 ;
  assign n28338 = n36722 & n28336 ;
  assign n28339 = n28337 | n28338 ;
  assign n28340 = n36681 & n28043 ;
  assign n28341 = n28188 | n28340 ;
  assign n36723 = ~n28187 ;
  assign n28342 = n36723 & n28341 ;
  assign n28343 = n28339 & n28342 ;
  assign n28344 = n28339 | n28342 ;
  assign n36724 = ~n28343 ;
  assign n28345 = n36724 & n28344 ;
  assign n36725 = ~n28211 ;
  assign n28346 = n36725 & n28345 ;
  assign n36726 = ~n28345 ;
  assign n28347 = n28211 & n36726 ;
  assign n29893 = n28346 | n28347 ;
  assign n36727 = ~n28313 ;
  assign n28348 = n36727 & n28320 ;
  assign n28349 = n28312 | n28348 ;
  assign n28350 = x11 | n28349 ;
  assign n28351 = x11 & n28349 ;
  assign n36728 = ~n28351 ;
  assign n28352 = n28350 & n36728 ;
  assign n28353 = n751 | n1010 ;
  assign n28354 = n1100 | n28353 ;
  assign n28355 = n2547 | n4602 ;
  assign n28356 = n28354 | n28355 ;
  assign n28357 = n1859 | n2427 ;
  assign n28358 = n2901 | n28357 ;
  assign n28359 = n1101 | n1160 ;
  assign n28360 = n1209 | n1694 ;
  assign n28361 = n28359 | n28360 ;
  assign n28362 = n28358 | n28361 ;
  assign n28363 = n28356 | n28362 ;
  assign n28364 = n11634 | n28363 ;
  assign n28365 = n22201 | n28364 ;
  assign n28366 = n27735 | n28365 ;
  assign n28367 = n3148 | n28366 ;
  assign n28368 = n28224 | n28367 ;
  assign n28369 = n28224 & n28367 ;
  assign n36729 = ~n28369 ;
  assign n28370 = n28368 & n36729 ;
  assign n36730 = ~n28212 ;
  assign n28371 = n36730 & n28224 ;
  assign n36731 = ~n28227 ;
  assign n28372 = n36731 & n28231 ;
  assign n28373 = n28371 | n28372 ;
  assign n36732 = ~n28373 ;
  assign n28374 = n28370 & n36732 ;
  assign n36733 = ~n28370 ;
  assign n28376 = n36733 & n28373 ;
  assign n28377 = n28374 | n28376 ;
  assign n21853 = n889 & n21848 ;
  assign n19679 = n3311 & n34360 ;
  assign n21776 = n3329 & n34803 ;
  assign n28378 = n19679 | n21776 ;
  assign n28379 = n3343 & n21753 ;
  assign n28380 = n28378 | n28379 ;
  assign n28381 = n21853 | n28380 ;
  assign n28382 = n28377 | n28381 ;
  assign n28383 = n28377 & n28381 ;
  assign n36734 = ~n28383 ;
  assign n28384 = n28382 & n36734 ;
  assign n22631 = n895 & n35030 ;
  assign n21750 = n2861 & n21729 ;
  assign n22544 = n2849 & n35018 ;
  assign n28385 = n21750 | n22544 ;
  assign n28386 = n894 & n22533 ;
  assign n28387 = n28385 | n28386 ;
  assign n28388 = n22631 | n28387 ;
  assign n36735 = ~n28388 ;
  assign n28389 = x29 & n36735 ;
  assign n28390 = n30024 & n28388 ;
  assign n28391 = n28389 | n28390 ;
  assign n36736 = ~n28391 ;
  assign n28392 = n28384 & n36736 ;
  assign n36737 = ~n28384 ;
  assign n28393 = n36737 & n28391 ;
  assign n28394 = n28392 | n28393 ;
  assign n36738 = ~n28239 ;
  assign n28395 = n36738 & n28246 ;
  assign n28396 = n28237 | n28395 ;
  assign n28397 = n28394 | n28396 ;
  assign n28398 = n28394 & n28396 ;
  assign n36739 = ~n28398 ;
  assign n28399 = n28397 & n36739 ;
  assign n23408 = n3791 & n35252 ;
  assign n22530 = n209 & n35020 ;
  assign n23344 = n3802 & n23339 ;
  assign n28400 = n22530 | n23344 ;
  assign n28401 = n3818 & n35254 ;
  assign n28402 = n28400 | n28401 ;
  assign n28403 = n23408 | n28402 ;
  assign n36740 = ~n28403 ;
  assign n28404 = x26 & n36740 ;
  assign n28405 = n30019 & n28403 ;
  assign n28406 = n28404 | n28405 ;
  assign n36741 = ~n28406 ;
  assign n28407 = n28399 & n36741 ;
  assign n36742 = ~n28399 ;
  assign n28408 = n36742 & n28406 ;
  assign n28409 = n28407 | n28408 ;
  assign n36743 = ~n28254 ;
  assign n28410 = n36743 & n28261 ;
  assign n28411 = n28252 | n28410 ;
  assign n36744 = ~n28411 ;
  assign n28412 = n28409 & n36744 ;
  assign n36745 = ~n28409 ;
  assign n28413 = n36745 & n28411 ;
  assign n28414 = n28412 | n28413 ;
  assign n24176 = n4135 & n24168 ;
  assign n23306 = n4185 & n35467 ;
  assign n24123 = n4148 & n35458 ;
  assign n28415 = n23306 | n24123 ;
  assign n28416 = n4165 & n24080 ;
  assign n28417 = n28415 | n28416 ;
  assign n28418 = n24176 | n28417 ;
  assign n36746 = ~n28418 ;
  assign n28419 = x23 & n36746 ;
  assign n28420 = n30030 & n28418 ;
  assign n28421 = n28419 | n28420 ;
  assign n36747 = ~n28421 ;
  assign n28422 = n28414 & n36747 ;
  assign n36748 = ~n28414 ;
  assign n28423 = n36748 & n28421 ;
  assign n28424 = n28422 | n28423 ;
  assign n36749 = ~n28266 ;
  assign n28425 = n28264 & n36749 ;
  assign n36750 = ~n28425 ;
  assign n28426 = n28277 & n36750 ;
  assign n36751 = ~n28424 ;
  assign n28427 = n36751 & n28426 ;
  assign n36752 = ~n28426 ;
  assign n28428 = n28424 & n36752 ;
  assign n28429 = n28427 | n28428 ;
  assign n25326 = n4686 & n35670 ;
  assign n24074 = n4726 & n24057 ;
  assign n24695 = n4706 & n24676 ;
  assign n28430 = n24074 | n24695 ;
  assign n28431 = n4748 & n35663 ;
  assign n28432 = n28430 | n28431 ;
  assign n28433 = n25326 | n28432 ;
  assign n36753 = ~n28433 ;
  assign n28434 = x20 & n36753 ;
  assign n28435 = n30374 & n28433 ;
  assign n28436 = n28434 | n28435 ;
  assign n36754 = ~n28436 ;
  assign n28437 = n28429 & n36754 ;
  assign n36755 = ~n28429 ;
  assign n28438 = n36755 & n28436 ;
  assign n28439 = n28437 | n28438 ;
  assign n36756 = ~n28280 ;
  assign n28440 = n28279 & n36756 ;
  assign n36757 = ~n28440 ;
  assign n28441 = n28291 & n36757 ;
  assign n36758 = ~n28439 ;
  assign n28442 = n36758 & n28441 ;
  assign n36759 = ~n28441 ;
  assign n28443 = n28439 & n36759 ;
  assign n28444 = n28442 | n28443 ;
  assign n25831 = n37300 & n35910 ;
  assign n24816 = n5166 & n24815 ;
  assign n25394 = n5144 & n35784 ;
  assign n28445 = n24816 | n25394 ;
  assign n28446 = n5191 & n25796 ;
  assign n28447 = n28445 | n28446 ;
  assign n28448 = n25831 | n28447 ;
  assign n36760 = ~n28448 ;
  assign n28449 = x17 & n36760 ;
  assign n28450 = n30580 & n28448 ;
  assign n28451 = n28449 | n28450 ;
  assign n28452 = n28444 | n28451 ;
  assign n28453 = n28444 & n28451 ;
  assign n36761 = ~n28453 ;
  assign n28454 = n28452 & n36761 ;
  assign n26492 = n5937 & n36130 ;
  assign n26049 = n5994 & n26039 ;
  assign n26475 = n5970 & n26278 ;
  assign n28455 = n26049 | n26475 ;
  assign n28456 = n6018 & n36131 ;
  assign n28457 = n28455 | n28456 ;
  assign n28458 = n26492 | n28457 ;
  assign n28459 = x14 | n28458 ;
  assign n28460 = x14 & n28458 ;
  assign n36762 = ~n28460 ;
  assign n28461 = n28459 & n36762 ;
  assign n36763 = ~n28296 ;
  assign n28462 = n36763 & n28306 ;
  assign n28463 = n28461 & n28462 ;
  assign n28464 = n28461 | n28462 ;
  assign n36764 = ~n28463 ;
  assign n28465 = n36764 & n28464 ;
  assign n28466 = n28454 & n28465 ;
  assign n28467 = n28454 | n28465 ;
  assign n36765 = ~n28466 ;
  assign n28468 = n36765 & n28467 ;
  assign n28469 = n28352 & n28468 ;
  assign n28470 = n28352 | n28468 ;
  assign n36766 = ~n28469 ;
  assign n28471 = n36766 & n28470 ;
  assign n28472 = n28327 | n28328 ;
  assign n28473 = n36719 & n28472 ;
  assign n36767 = ~n28471 ;
  assign n28474 = n36767 & n28473 ;
  assign n36768 = ~n28473 ;
  assign n28475 = n28471 & n36768 ;
  assign n28476 = n28474 | n28475 ;
  assign n28477 = n36723 & n28208 ;
  assign n28478 = n28339 | n28477 ;
  assign n36769 = ~n28337 ;
  assign n28479 = n36769 & n28478 ;
  assign n36770 = ~n28476 ;
  assign n28480 = n36770 & n28479 ;
  assign n36771 = ~n28479 ;
  assign n28481 = n28476 & n36771 ;
  assign n28482 = n28480 | n28481 ;
  assign n28483 = n28347 | n28482 ;
  assign n28484 = n28347 & n28482 ;
  assign n36772 = ~n28484 ;
  assign n48 = n28483 & n36772 ;
  assign n24148 = n4135 & n35457 ;
  assign n24096 = n4148 & n24080 ;
  assign n24106 = n4185 & n35458 ;
  assign n28485 = n24096 | n24106 ;
  assign n28486 = n4165 & n24151 ;
  assign n28487 = n28485 | n28486 ;
  assign n28488 = n24148 | n28487 ;
  assign n36773 = ~n28488 ;
  assign n28489 = x23 & n36773 ;
  assign n28490 = n30030 & n28488 ;
  assign n28491 = n28489 | n28490 ;
  assign n28492 = n931 | n2559 ;
  assign n28493 = n2951 | n28492 ;
  assign n28494 = n2079 | n28493 ;
  assign n28495 = n23805 | n28494 ;
  assign n28496 = n439 | n540 ;
  assign n28497 = n630 | n841 ;
  assign n28498 = n28496 | n28497 ;
  assign n28499 = n488 | n858 ;
  assign n28500 = n28498 | n28499 ;
  assign n28501 = n2987 | n28500 ;
  assign n28502 = n3012 | n28501 ;
  assign n28503 = n28495 | n28502 ;
  assign n28504 = n1237 | n28503 ;
  assign n36774 = ~n28504 ;
  assign n28505 = n1291 & n36774 ;
  assign n36775 = ~n4607 ;
  assign n28506 = n36775 & n28505 ;
  assign n28507 = x11 & n28506 ;
  assign n28508 = x11 | n28506 ;
  assign n36776 = ~n28507 ;
  assign n28509 = n36776 & n28508 ;
  assign n36777 = ~n28224 ;
  assign n28510 = n36777 & n28509 ;
  assign n36778 = ~n28509 ;
  assign n28511 = n28224 & n36778 ;
  assign n28512 = n28510 | n28511 ;
  assign n28375 = n28369 | n28373 ;
  assign n28513 = n28368 & n28375 ;
  assign n36779 = ~n28512 ;
  assign n28514 = n36779 & n28513 ;
  assign n36780 = ~n28513 ;
  assign n28515 = n28512 & n36780 ;
  assign n28516 = n28514 | n28515 ;
  assign n21801 = n889 & n34802 ;
  assign n21758 = n3311 & n34803 ;
  assign n21826 = n3329 & n21753 ;
  assign n28517 = n21758 | n21826 ;
  assign n28518 = n3343 & n21804 ;
  assign n28519 = n28517 | n28518 ;
  assign n28520 = n21801 | n28519 ;
  assign n28521 = n28516 | n28520 ;
  assign n28522 = n28516 & n28520 ;
  assign n36781 = ~n28522 ;
  assign n28523 = n28521 & n36781 ;
  assign n36782 = ~n28392 ;
  assign n28524 = n28382 & n36782 ;
  assign n28525 = n28523 & n28524 ;
  assign n28526 = n28523 | n28524 ;
  assign n36783 = ~n28525 ;
  assign n28527 = n36783 & n28526 ;
  assign n22575 = n895 & n35022 ;
  assign n22556 = n2861 & n35018 ;
  assign n22600 = n2849 & n22533 ;
  assign n28528 = n22556 | n22600 ;
  assign n28529 = n894 & n35020 ;
  assign n28530 = n28528 | n28529 ;
  assign n28531 = n22575 | n28530 ;
  assign n36784 = ~n28531 ;
  assign n28532 = x29 & n36784 ;
  assign n28533 = n30024 & n28531 ;
  assign n28534 = n28532 | n28533 ;
  assign n28535 = n28527 | n28534 ;
  assign n28536 = n28527 & n28534 ;
  assign n36785 = ~n28536 ;
  assign n28537 = n28535 & n36785 ;
  assign n23379 = n3791 & n23372 ;
  assign n23329 = n3802 & n35244 ;
  assign n23361 = n209 & n23339 ;
  assign n28538 = n23329 | n23361 ;
  assign n28539 = n3818 & n35246 ;
  assign n28540 = n28538 | n28539 ;
  assign n28541 = n23379 | n28540 ;
  assign n36786 = ~n28541 ;
  assign n28542 = x26 & n36786 ;
  assign n28543 = n30019 & n28541 ;
  assign n28544 = n28542 | n28543 ;
  assign n28545 = n28399 & n28406 ;
  assign n28546 = n28398 | n28545 ;
  assign n28547 = n28544 | n28546 ;
  assign n28548 = n28544 & n28546 ;
  assign n36787 = ~n28548 ;
  assign n28549 = n28547 & n36787 ;
  assign n28550 = n28537 & n28549 ;
  assign n28551 = n28537 | n28549 ;
  assign n36788 = ~n28550 ;
  assign n28552 = n36788 & n28551 ;
  assign n28553 = n28409 | n28411 ;
  assign n36789 = ~n28422 ;
  assign n28554 = n36789 & n28553 ;
  assign n28555 = n28552 & n28554 ;
  assign n28556 = n28552 | n28554 ;
  assign n36790 = ~n28555 ;
  assign n28557 = n36790 & n28556 ;
  assign n28558 = n28491 | n28557 ;
  assign n28559 = n28491 & n28557 ;
  assign n36791 = ~n28559 ;
  assign n28560 = n28558 & n36791 ;
  assign n24882 = n4686 & n35662 ;
  assign n24696 = n4726 & n24676 ;
  assign n24853 = n4706 & n35663 ;
  assign n28561 = n24696 | n24853 ;
  assign n28562 = n4748 & n24815 ;
  assign n28563 = n28561 | n28562 ;
  assign n28564 = n24882 | n28563 ;
  assign n36792 = ~n28564 ;
  assign n28565 = x20 & n36792 ;
  assign n28566 = n30374 & n28564 ;
  assign n28567 = n28565 | n28566 ;
  assign n36793 = ~n28567 ;
  assign n28568 = n28560 & n36793 ;
  assign n36794 = ~n28560 ;
  assign n28569 = n36794 & n28567 ;
  assign n28570 = n28568 | n28569 ;
  assign n28571 = n28424 | n28426 ;
  assign n36795 = ~n28437 ;
  assign n28572 = n36795 & n28571 ;
  assign n36796 = ~n28570 ;
  assign n28573 = n36796 & n28572 ;
  assign n36797 = ~n28572 ;
  assign n28574 = n28570 & n36797 ;
  assign n28575 = n28573 | n28574 ;
  assign n26068 = n37300 & n26065 ;
  assign n25399 = n5166 & n35784 ;
  assign n25804 = n5144 & n25796 ;
  assign n28576 = n25399 | n25804 ;
  assign n28577 = n5191 & n26039 ;
  assign n28578 = n28576 | n28577 ;
  assign n28579 = n26068 | n28578 ;
  assign n36798 = ~n28579 ;
  assign n28580 = x17 & n36798 ;
  assign n28581 = n30580 & n28579 ;
  assign n28582 = n28580 | n28581 ;
  assign n36799 = ~n28582 ;
  assign n28583 = n28575 & n36799 ;
  assign n36800 = ~n28575 ;
  assign n28584 = n36800 & n28582 ;
  assign n28585 = n28583 | n28584 ;
  assign n28586 = n28439 | n28441 ;
  assign n36801 = ~n28451 ;
  assign n28587 = n28444 & n36801 ;
  assign n36802 = ~n28587 ;
  assign n28588 = n28586 & n36802 ;
  assign n36803 = ~n28585 ;
  assign n28589 = n36803 & n28588 ;
  assign n36804 = ~n28588 ;
  assign n28590 = n28585 & n36804 ;
  assign n28591 = n28589 | n28590 ;
  assign n26700 = n5937 & n36192 ;
  assign n28592 = n5994 & n26278 ;
  assign n28593 = n5970 & n36131 ;
  assign n28594 = n28592 | n28593 ;
  assign n28595 = n26700 | n28594 ;
  assign n36805 = ~n28595 ;
  assign n28596 = x14 & n36805 ;
  assign n28597 = n30547 & n28595 ;
  assign n28598 = n28596 | n28597 ;
  assign n28599 = n28463 | n28466 ;
  assign n28600 = n28598 | n28599 ;
  assign n28601 = n28598 & n28599 ;
  assign n36806 = ~n28601 ;
  assign n28602 = n28600 & n36806 ;
  assign n28603 = n28591 & n28602 ;
  assign n28605 = n28591 | n28602 ;
  assign n36807 = ~n28603 ;
  assign n28606 = n36807 & n28605 ;
  assign n36808 = ~n28468 ;
  assign n28607 = n28352 & n36808 ;
  assign n36809 = ~n28607 ;
  assign n28608 = n28350 & n36809 ;
  assign n36810 = ~n28606 ;
  assign n28609 = n36810 & n28608 ;
  assign n36811 = ~n28608 ;
  assign n28610 = n28606 & n36811 ;
  assign n28611 = n28609 | n28610 ;
  assign n28612 = n28471 | n28473 ;
  assign n28613 = n36769 & n28344 ;
  assign n36812 = ~n28613 ;
  assign n28614 = n28476 & n36812 ;
  assign n36813 = ~n28614 ;
  assign n28615 = n28612 & n36813 ;
  assign n28616 = n28611 & n28615 ;
  assign n28617 = n28611 | n28615 ;
  assign n36814 = ~n28616 ;
  assign n28618 = n36814 & n28617 ;
  assign n28619 = n36772 & n28618 ;
  assign n36815 = ~n28618 ;
  assign n28620 = n28484 & n36815 ;
  assign n29891 = n28619 | n28620 ;
  assign n36816 = ~n28515 ;
  assign n28621 = n36816 & n28521 ;
  assign n36817 = ~n28510 ;
  assign n28622 = n28508 & n36817 ;
  assign n28623 = n1271 | n2203 ;
  assign n28624 = n107 | n263 ;
  assign n28625 = n446 | n28624 ;
  assign n28626 = n590 | n1982 ;
  assign n28627 = n28625 | n28626 ;
  assign n28628 = n23178 | n28627 ;
  assign n28629 = n28623 | n28628 ;
  assign n28630 = n1363 | n3449 ;
  assign n28631 = n5839 | n28630 ;
  assign n28632 = n26903 | n28631 ;
  assign n28633 = n28629 | n28632 ;
  assign n28634 = n26543 | n28633 ;
  assign n28635 = n11636 | n23811 ;
  assign n28636 = n28634 | n28635 ;
  assign n28637 = n28622 & n28636 ;
  assign n28638 = n28622 | n28636 ;
  assign n36818 = ~n28637 ;
  assign n28639 = n36818 & n28638 ;
  assign n22654 = n889 & n35035 ;
  assign n21751 = n3329 & n21729 ;
  assign n21827 = n3311 & n21753 ;
  assign n28640 = n21751 | n21827 ;
  assign n28641 = n3343 & n35018 ;
  assign n28642 = n28640 | n28641 ;
  assign n28643 = n22654 | n28642 ;
  assign n36819 = ~n28643 ;
  assign n28644 = n28639 & n36819 ;
  assign n36820 = ~n28639 ;
  assign n28646 = n36820 & n28643 ;
  assign n28647 = n28644 | n28646 ;
  assign n28648 = n28621 & n28647 ;
  assign n28649 = n28621 | n28647 ;
  assign n36821 = ~n28648 ;
  assign n28650 = n36821 & n28649 ;
  assign n23437 = n895 & n35262 ;
  assign n22513 = n2849 & n35020 ;
  assign n22592 = n2861 & n22533 ;
  assign n28651 = n22513 | n22592 ;
  assign n28652 = n894 & n23444 ;
  assign n28653 = n28651 | n28652 ;
  assign n28654 = n23437 | n28653 ;
  assign n36822 = ~n28654 ;
  assign n28655 = x29 & n36822 ;
  assign n28656 = n30024 & n28654 ;
  assign n28657 = n28655 | n28656 ;
  assign n36823 = ~n28657 ;
  assign n28658 = n28650 & n36823 ;
  assign n36824 = ~n28650 ;
  assign n28659 = n36824 & n28657 ;
  assign n28660 = n28658 | n28659 ;
  assign n36825 = ~n28524 ;
  assign n28661 = n28523 & n36825 ;
  assign n36826 = ~n28661 ;
  assign n28662 = n28535 & n36826 ;
  assign n36827 = ~n28660 ;
  assign n28663 = n36827 & n28662 ;
  assign n36828 = ~n28662 ;
  assign n28664 = n28660 & n36828 ;
  assign n28665 = n28663 | n28664 ;
  assign n24204 = n3791 & n35472 ;
  assign n23309 = n3802 & n35467 ;
  assign n23335 = n209 & n35244 ;
  assign n28666 = n23309 | n23335 ;
  assign n28667 = n3818 & n35465 ;
  assign n28668 = n28666 | n28667 ;
  assign n28669 = n24204 | n28668 ;
  assign n36829 = ~n28669 ;
  assign n28670 = x26 & n36829 ;
  assign n28671 = n30019 & n28669 ;
  assign n28672 = n28670 | n28671 ;
  assign n36830 = ~n28672 ;
  assign n28673 = n28665 & n36830 ;
  assign n36831 = ~n28665 ;
  assign n28674 = n36831 & n28672 ;
  assign n28675 = n28673 | n28674 ;
  assign n28676 = n28547 & n36788 ;
  assign n36832 = ~n28675 ;
  assign n28677 = n36832 & n28676 ;
  assign n36833 = ~n28676 ;
  assign n28678 = n28675 & n36833 ;
  assign n28679 = n28677 | n28678 ;
  assign n25296 = n4135 & n25288 ;
  assign n24068 = n4148 & n24057 ;
  assign n24097 = n4185 & n24080 ;
  assign n28680 = n24068 | n24097 ;
  assign n28681 = n4165 & n24676 ;
  assign n28682 = n28680 | n28681 ;
  assign n28683 = n25296 | n28682 ;
  assign n36834 = ~n28683 ;
  assign n28684 = x23 & n36834 ;
  assign n28685 = n30030 & n28683 ;
  assign n28686 = n28684 | n28685 ;
  assign n36835 = ~n28686 ;
  assign n28687 = n28679 & n36835 ;
  assign n36836 = ~n28679 ;
  assign n28688 = n36836 & n28686 ;
  assign n28689 = n28687 | n28688 ;
  assign n36837 = ~n28552 ;
  assign n28690 = n36837 & n28554 ;
  assign n36838 = ~n28557 ;
  assign n28691 = n28491 & n36838 ;
  assign n28692 = n28690 | n28691 ;
  assign n28693 = n28689 | n28692 ;
  assign n28694 = n28689 & n28692 ;
  assign n36839 = ~n28694 ;
  assign n28695 = n28693 & n36839 ;
  assign n25428 = n4686 & n35785 ;
  assign n24826 = n4706 & n24815 ;
  assign n24854 = n4726 & n35663 ;
  assign n28696 = n24826 | n24854 ;
  assign n28697 = n4748 & n35784 ;
  assign n28698 = n28696 | n28697 ;
  assign n28699 = n25428 | n28698 ;
  assign n36840 = ~n28699 ;
  assign n28700 = x20 & n36840 ;
  assign n28701 = n30374 & n28699 ;
  assign n28702 = n28700 | n28701 ;
  assign n36841 = ~n28702 ;
  assign n28703 = n28695 & n36841 ;
  assign n36842 = ~n28695 ;
  assign n28704 = n36842 & n28702 ;
  assign n28705 = n28703 | n28704 ;
  assign n28706 = n28570 | n28572 ;
  assign n36843 = ~n28568 ;
  assign n28707 = n36843 & n28706 ;
  assign n36844 = ~n28705 ;
  assign n28708 = n36844 & n28707 ;
  assign n36845 = ~n28707 ;
  assign n28709 = n28705 & n36845 ;
  assign n28710 = n28708 | n28709 ;
  assign n26289 = n37300 & n26284 ;
  assign n25803 = n5166 & n25796 ;
  assign n26042 = n5144 & n26039 ;
  assign n28711 = n25803 | n26042 ;
  assign n28712 = n5191 & n26278 ;
  assign n28713 = n28711 | n28712 ;
  assign n28714 = n26289 | n28713 ;
  assign n36846 = ~n28714 ;
  assign n28715 = x17 & n36846 ;
  assign n28716 = n30580 & n28714 ;
  assign n28717 = n28715 | n28716 ;
  assign n36847 = ~n28717 ;
  assign n28718 = n28710 & n36847 ;
  assign n36848 = ~n28710 ;
  assign n28719 = n36848 & n28717 ;
  assign n28720 = n28718 | n28719 ;
  assign n28721 = n5992 | n26279 ;
  assign n28722 = n30547 & n28721 ;
  assign n28723 = x13 | n28721 ;
  assign n36849 = ~n28722 ;
  assign n28724 = n36849 & n28723 ;
  assign n28725 = n28585 | n28588 ;
  assign n36850 = ~n28583 ;
  assign n28726 = n36850 & n28725 ;
  assign n28727 = n28724 & n28726 ;
  assign n28728 = n28724 | n28726 ;
  assign n36851 = ~n28727 ;
  assign n28729 = n36851 & n28728 ;
  assign n36852 = ~n28720 ;
  assign n28730 = n36852 & n28729 ;
  assign n36853 = ~n28729 ;
  assign n28731 = n28720 & n36853 ;
  assign n28732 = n28730 | n28731 ;
  assign n36854 = ~n28591 ;
  assign n28604 = n36854 & n28602 ;
  assign n28733 = n28601 | n28604 ;
  assign n28734 = n28732 & n28733 ;
  assign n28735 = n28732 | n28733 ;
  assign n36855 = ~n28734 ;
  assign n28736 = n36855 & n28735 ;
  assign n36856 = ~n28481 ;
  assign n28737 = n36856 & n28612 ;
  assign n28738 = n28611 | n28737 ;
  assign n36857 = ~n28610 ;
  assign n28739 = n36857 & n28738 ;
  assign n36858 = ~n28736 ;
  assign n28740 = n36858 & n28739 ;
  assign n36859 = ~n28739 ;
  assign n28741 = n28736 & n36859 ;
  assign n28742 = n28740 | n28741 ;
  assign n28743 = n28620 | n28742 ;
  assign n28744 = n28620 & n28742 ;
  assign n36860 = ~n28744 ;
  assign n50 = n28743 & n36860 ;
  assign n28745 = n3292 & n30400 ;
  assign n36861 = ~n13951 ;
  assign n28746 = n36861 & n28745 ;
  assign n28747 = n220 | n253 ;
  assign n28748 = n354 | n660 ;
  assign n28749 = n28747 | n28748 ;
  assign n28750 = n124 | n242 ;
  assign n28751 = n28749 | n28750 ;
  assign n28752 = n1641 | n28751 ;
  assign n28753 = n666 | n1894 ;
  assign n28754 = n5816 | n28753 ;
  assign n28755 = n2081 | n28754 ;
  assign n28756 = n28752 | n28755 ;
  assign n28757 = n2753 | n28756 ;
  assign n28758 = n14325 | n28757 ;
  assign n36862 = ~n28758 ;
  assign n28759 = n28746 & n36862 ;
  assign n28760 = n34912 & n28759 ;
  assign n28761 = n28636 | n28760 ;
  assign n28762 = n28636 & n28760 ;
  assign n36863 = ~n28762 ;
  assign n28763 = n28761 & n36863 ;
  assign n22629 = n889 & n35030 ;
  assign n21743 = n3311 & n21729 ;
  assign n22538 = n3329 & n35018 ;
  assign n28764 = n21743 | n22538 ;
  assign n28765 = n3343 & n22533 ;
  assign n28766 = n28764 | n28765 ;
  assign n28767 = n22629 | n28766 ;
  assign n36864 = ~n28767 ;
  assign n28768 = n28763 & n36864 ;
  assign n36865 = ~n28763 ;
  assign n28770 = n36865 & n28767 ;
  assign n28771 = n28768 | n28770 ;
  assign n28645 = n28638 & n36819 ;
  assign n28772 = n28637 | n28645 ;
  assign n36866 = ~n28772 ;
  assign n28773 = n28771 & n36866 ;
  assign n36867 = ~n28771 ;
  assign n28774 = n36867 & n28772 ;
  assign n28775 = n28773 | n28774 ;
  assign n28776 = n28650 & n28657 ;
  assign n28777 = n28648 | n28776 ;
  assign n36868 = ~n28777 ;
  assign n28778 = n28775 & n36868 ;
  assign n36869 = ~n28775 ;
  assign n28779 = n36869 & n28777 ;
  assign n28780 = n28778 | n28779 ;
  assign n23413 = n895 & n35252 ;
  assign n22529 = n2861 & n35020 ;
  assign n23345 = n2849 & n23339 ;
  assign n28781 = n22529 | n23345 ;
  assign n28782 = n894 & n35254 ;
  assign n28783 = n28781 | n28782 ;
  assign n28784 = n23413 | n28783 ;
  assign n28785 = x29 | n28784 ;
  assign n28786 = x29 & n28784 ;
  assign n36870 = ~n28786 ;
  assign n28787 = n28785 & n36870 ;
  assign n36871 = ~n28780 ;
  assign n28788 = n36871 & n28787 ;
  assign n36872 = ~n28787 ;
  assign n28789 = n28780 & n36872 ;
  assign n28790 = n28788 | n28789 ;
  assign n24177 = n3791 & n24168 ;
  assign n23310 = n209 & n35467 ;
  assign n24108 = n3802 & n35458 ;
  assign n28791 = n23310 | n24108 ;
  assign n28792 = n3818 & n24080 ;
  assign n28793 = n28791 | n28792 ;
  assign n28794 = n24177 | n28793 ;
  assign n36873 = ~n28794 ;
  assign n28795 = x26 & n36873 ;
  assign n28796 = n30019 & n28794 ;
  assign n28797 = n28795 | n28796 ;
  assign n28798 = n28790 | n28797 ;
  assign n28799 = n28790 & n28797 ;
  assign n36874 = ~n28799 ;
  assign n28800 = n28798 & n36874 ;
  assign n28801 = n28660 | n28662 ;
  assign n36875 = ~n28673 ;
  assign n28802 = n36875 & n28801 ;
  assign n36876 = ~n28800 ;
  assign n28803 = n36876 & n28802 ;
  assign n36877 = ~n28802 ;
  assign n28804 = n28800 & n36877 ;
  assign n28805 = n28803 | n28804 ;
  assign n25327 = n4135 & n35670 ;
  assign n24063 = n4185 & n24057 ;
  assign n24686 = n4148 & n24676 ;
  assign n28806 = n24063 | n24686 ;
  assign n28807 = n4165 & n35663 ;
  assign n28808 = n28806 | n28807 ;
  assign n28809 = n25327 | n28808 ;
  assign n36878 = ~n28809 ;
  assign n28810 = x23 & n36878 ;
  assign n28811 = n30030 & n28809 ;
  assign n28812 = n28810 | n28811 ;
  assign n28813 = n28805 | n28812 ;
  assign n28814 = n28805 & n28812 ;
  assign n36879 = ~n28814 ;
  assign n28815 = n28813 & n36879 ;
  assign n28816 = n28675 | n28676 ;
  assign n36880 = ~n28687 ;
  assign n28817 = n36880 & n28816 ;
  assign n28818 = n28815 & n28817 ;
  assign n28819 = n28815 | n28817 ;
  assign n36881 = ~n28818 ;
  assign n28820 = n36881 & n28819 ;
  assign n25833 = n4686 & n35910 ;
  assign n24819 = n4726 & n24815 ;
  assign n25402 = n4706 & n35784 ;
  assign n28821 = n24819 | n25402 ;
  assign n28822 = n4748 & n25796 ;
  assign n28823 = n28821 | n28822 ;
  assign n28824 = n25833 | n28823 ;
  assign n36882 = ~n28824 ;
  assign n28825 = x20 & n36882 ;
  assign n28826 = n30374 & n28824 ;
  assign n28827 = n28825 | n28826 ;
  assign n36883 = ~n28827 ;
  assign n28828 = n28820 & n36883 ;
  assign n36884 = ~n28820 ;
  assign n28829 = n36884 & n28827 ;
  assign n28830 = n28828 | n28829 ;
  assign n26493 = n37300 & n36130 ;
  assign n26040 = n5166 & n26039 ;
  assign n26478 = n5144 & n26278 ;
  assign n28831 = n26040 | n26478 ;
  assign n28832 = n5191 & n36131 ;
  assign n28833 = n28831 | n28832 ;
  assign n28834 = n26493 | n28833 ;
  assign n28835 = x17 | n28834 ;
  assign n28836 = x17 & n28834 ;
  assign n36885 = ~n28836 ;
  assign n28837 = n28835 & n36885 ;
  assign n36886 = ~n28703 ;
  assign n28838 = n28693 & n36886 ;
  assign n28839 = n28837 & n28838 ;
  assign n28840 = n28837 | n28838 ;
  assign n36887 = ~n28839 ;
  assign n28841 = n36887 & n28840 ;
  assign n36888 = ~n28830 ;
  assign n28842 = n36888 & n28841 ;
  assign n36889 = ~n28841 ;
  assign n28843 = n28830 & n36889 ;
  assign n28844 = n28842 | n28843 ;
  assign n28845 = n28705 | n28707 ;
  assign n36890 = ~n28718 ;
  assign n28846 = n36890 & n28845 ;
  assign n28847 = x14 & n28846 ;
  assign n28848 = x14 | n28846 ;
  assign n36891 = ~n28847 ;
  assign n28849 = n36891 & n28848 ;
  assign n28850 = n28844 & n28849 ;
  assign n28851 = n28844 | n28849 ;
  assign n36892 = ~n28850 ;
  assign n28852 = n36892 & n28851 ;
  assign n28853 = n28720 & n28729 ;
  assign n28854 = n28727 | n28853 ;
  assign n36893 = ~n28854 ;
  assign n28855 = n28852 & n36893 ;
  assign n36894 = ~n28852 ;
  assign n28856 = n36894 & n28854 ;
  assign n28857 = n28855 | n28856 ;
  assign n28858 = n36857 & n28617 ;
  assign n28859 = n28734 | n28858 ;
  assign n28860 = n28735 & n28859 ;
  assign n28861 = n28857 & n28860 ;
  assign n28862 = n28857 | n28860 ;
  assign n36895 = ~n28861 ;
  assign n28863 = n36895 & n28862 ;
  assign n28864 = n28744 & n28863 ;
  assign n29888 = n28744 | n28863 ;
  assign n36896 = ~n28864 ;
  assign n29889 = n36896 & n29888 ;
  assign n36897 = ~n28863 ;
  assign n28865 = n28744 & n36897 ;
  assign n28866 = n2678 | n12830 ;
  assign n28867 = n13595 | n28866 ;
  assign n1299 = n683 | n698 ;
  assign n28868 = n200 | n220 ;
  assign n28869 = n495 | n28868 ;
  assign n28870 = n1299 | n28869 ;
  assign n28871 = n2147 | n28870 ;
  assign n28872 = n3756 | n28871 ;
  assign n36898 = ~n28872 ;
  assign n28873 = n5586 & n36898 ;
  assign n36899 = ~n28867 ;
  assign n28874 = n36899 & n28873 ;
  assign n36900 = ~n21602 ;
  assign n28875 = n36900 & n28874 ;
  assign n36901 = ~n1173 ;
  assign n28876 = n36901 & n28875 ;
  assign n36902 = ~n28636 ;
  assign n28877 = n36902 & n28876 ;
  assign n36903 = ~n28876 ;
  assign n28878 = n28636 & n36903 ;
  assign n28879 = n28877 | n28878 ;
  assign n28880 = x14 | n28879 ;
  assign n28881 = x14 & n28879 ;
  assign n36904 = ~n28881 ;
  assign n28882 = n28880 & n36904 ;
  assign n28769 = n28761 & n36864 ;
  assign n28883 = n28762 | n28769 ;
  assign n36905 = ~n28883 ;
  assign n28884 = n28882 & n36905 ;
  assign n36906 = ~n28882 ;
  assign n28885 = n36906 & n28883 ;
  assign n28886 = n28884 | n28885 ;
  assign n22576 = n889 & n35022 ;
  assign n22552 = n3311 & n35018 ;
  assign n22596 = n3329 & n22533 ;
  assign n28887 = n22552 | n22596 ;
  assign n28888 = n3343 & n35020 ;
  assign n28889 = n28887 | n28888 ;
  assign n28890 = n22576 | n28889 ;
  assign n28891 = n28886 | n28890 ;
  assign n28892 = n28886 & n28890 ;
  assign n36907 = ~n28892 ;
  assign n28893 = n28891 & n36907 ;
  assign n23382 = n895 & n23372 ;
  assign n23336 = n2849 & n35244 ;
  assign n23347 = n2861 & n23339 ;
  assign n28894 = n23336 | n23347 ;
  assign n28895 = n894 & n35246 ;
  assign n28896 = n28894 | n28895 ;
  assign n28897 = n23382 | n28896 ;
  assign n28898 = x29 | n28897 ;
  assign n28899 = x29 & n28897 ;
  assign n36908 = ~n28899 ;
  assign n28900 = n28898 & n36908 ;
  assign n28901 = n28893 & n28900 ;
  assign n28902 = n28893 | n28900 ;
  assign n36909 = ~n28901 ;
  assign n28903 = n36909 & n28902 ;
  assign n28904 = n28775 | n28777 ;
  assign n36910 = ~n28774 ;
  assign n28905 = n36910 & n28904 ;
  assign n36911 = ~n28903 ;
  assign n28906 = n36911 & n28905 ;
  assign n36912 = ~n28905 ;
  assign n28907 = n28903 & n36912 ;
  assign n28908 = n28906 | n28907 ;
  assign n24149 = n3791 & n35457 ;
  assign n24093 = n3802 & n24080 ;
  assign n24117 = n209 & n35458 ;
  assign n28909 = n24093 | n24117 ;
  assign n28910 = n3818 & n24151 ;
  assign n28911 = n28909 | n28910 ;
  assign n28912 = n24149 | n28911 ;
  assign n28913 = x26 | n28912 ;
  assign n28914 = x26 & n28912 ;
  assign n36913 = ~n28914 ;
  assign n28915 = n28913 & n36913 ;
  assign n36914 = ~n28790 ;
  assign n28916 = n36914 & n28797 ;
  assign n28917 = n28788 | n28916 ;
  assign n36915 = ~n28917 ;
  assign n28918 = n28915 & n36915 ;
  assign n36916 = ~n28915 ;
  assign n28919 = n36916 & n28917 ;
  assign n28920 = n28918 | n28919 ;
  assign n28921 = n28908 & n28920 ;
  assign n28922 = n28908 | n28920 ;
  assign n36917 = ~n28921 ;
  assign n28923 = n36917 & n28922 ;
  assign n24877 = n4135 & n35662 ;
  assign n24684 = n4185 & n24676 ;
  assign n24856 = n4148 & n35663 ;
  assign n28924 = n24684 | n24856 ;
  assign n28925 = n4165 & n24815 ;
  assign n28926 = n28924 | n28925 ;
  assign n28927 = n24877 | n28926 ;
  assign n36918 = ~n28927 ;
  assign n28928 = x23 & n36918 ;
  assign n28929 = n30030 & n28927 ;
  assign n28930 = n28928 | n28929 ;
  assign n36919 = ~n28930 ;
  assign n28931 = n28923 & n36919 ;
  assign n36920 = ~n28923 ;
  assign n28932 = n36920 & n28930 ;
  assign n28933 = n28931 | n28932 ;
  assign n36921 = ~n28804 ;
  assign n28934 = n36921 & n28813 ;
  assign n36922 = ~n28933 ;
  assign n28935 = n36922 & n28934 ;
  assign n36923 = ~n28934 ;
  assign n28936 = n28933 & n36923 ;
  assign n28937 = n28935 | n28936 ;
  assign n26073 = n4686 & n26065 ;
  assign n25410 = n4726 & n35784 ;
  assign n25802 = n4706 & n25796 ;
  assign n28938 = n25410 | n25802 ;
  assign n28939 = n4748 & n26039 ;
  assign n28940 = n28938 | n28939 ;
  assign n28941 = n26073 | n28940 ;
  assign n36924 = ~n28941 ;
  assign n28942 = x20 & n36924 ;
  assign n28943 = n30374 & n28941 ;
  assign n28944 = n28942 | n28943 ;
  assign n36925 = ~n28944 ;
  assign n28945 = n28937 & n36925 ;
  assign n36926 = ~n28937 ;
  assign n28946 = n36926 & n28944 ;
  assign n28947 = n28945 | n28946 ;
  assign n36927 = ~n28817 ;
  assign n28948 = n28815 & n36927 ;
  assign n28949 = n28820 | n28827 ;
  assign n36928 = ~n28948 ;
  assign n28950 = n36928 & n28949 ;
  assign n36929 = ~n28947 ;
  assign n28951 = n36929 & n28950 ;
  assign n36930 = ~n28950 ;
  assign n28952 = n28947 & n36930 ;
  assign n28953 = n28951 | n28952 ;
  assign n26703 = n37300 & n36192 ;
  assign n28954 = n5166 & n26278 ;
  assign n28955 = n5144 & n36131 ;
  assign n28956 = n28954 | n28955 ;
  assign n28957 = n26703 | n28956 ;
  assign n28958 = x17 | n28957 ;
  assign n28959 = x17 & n28957 ;
  assign n36931 = ~n28959 ;
  assign n28960 = n28958 & n36931 ;
  assign n28961 = n28839 | n28842 ;
  assign n36932 = ~n28961 ;
  assign n28962 = n28960 & n36932 ;
  assign n36933 = ~n28960 ;
  assign n28963 = n36933 & n28961 ;
  assign n28964 = n28962 | n28963 ;
  assign n28965 = n28953 & n28964 ;
  assign n28967 = n28953 | n28964 ;
  assign n36934 = ~n28965 ;
  assign n28968 = n36934 & n28967 ;
  assign n28969 = n28848 & n36892 ;
  assign n36935 = ~n28968 ;
  assign n28970 = n36935 & n28969 ;
  assign n36936 = ~n28969 ;
  assign n28971 = n28968 & n36936 ;
  assign n28972 = n28970 | n28971 ;
  assign n28973 = n28734 | n28739 ;
  assign n28974 = n28735 & n28973 ;
  assign n28975 = n28856 | n28974 ;
  assign n36937 = ~n28855 ;
  assign n28976 = n36937 & n28975 ;
  assign n28977 = n28972 & n28976 ;
  assign n28978 = n28972 | n28976 ;
  assign n36938 = ~n28977 ;
  assign n28979 = n36938 & n28978 ;
  assign n36939 = ~n28865 ;
  assign n28980 = n36939 & n28979 ;
  assign n36940 = ~n28979 ;
  assign n28981 = n28865 & n36940 ;
  assign n29887 = n28980 | n28981 ;
  assign n36941 = ~n28885 ;
  assign n28982 = n36941 & n28891 ;
  assign n36942 = ~n28878 ;
  assign n28983 = n36942 & n28880 ;
  assign n28984 = n221 | n540 ;
  assign n28985 = n662 | n28984 ;
  assign n28986 = n1310 | n28985 ;
  assign n28987 = n4020 | n20723 ;
  assign n28988 = n28986 | n28987 ;
  assign n28989 = n1718 | n2243 ;
  assign n28990 = n4596 | n13562 ;
  assign n28991 = n28989 | n28990 ;
  assign n28992 = n5029 | n28991 ;
  assign n28993 = n28988 | n28992 ;
  assign n28994 = n505 | n3571 ;
  assign n28995 = n28993 | n28994 ;
  assign n28996 = n3027 | n28995 ;
  assign n36943 = ~n28996 ;
  assign n28997 = n2402 & n36943 ;
  assign n36944 = ~n28983 ;
  assign n28998 = n36944 & n28997 ;
  assign n36945 = ~n28997 ;
  assign n28999 = n28983 & n36945 ;
  assign n29000 = n28998 | n28999 ;
  assign n23443 = n889 & n35262 ;
  assign n22523 = n3329 & n35020 ;
  assign n22599 = n3311 & n22533 ;
  assign n29001 = n22523 | n22599 ;
  assign n29002 = n3343 & n23444 ;
  assign n29003 = n29001 | n29002 ;
  assign n29004 = n23443 | n29003 ;
  assign n36946 = ~n29004 ;
  assign n29005 = n29000 & n36946 ;
  assign n36947 = ~n29000 ;
  assign n29007 = n36947 & n29004 ;
  assign n29008 = n29005 | n29007 ;
  assign n29009 = n28982 | n29008 ;
  assign n29010 = n28982 & n29008 ;
  assign n36948 = ~n29010 ;
  assign n29011 = n29009 & n36948 ;
  assign n24199 = n895 & n35472 ;
  assign n23311 = n2849 & n35467 ;
  assign n23324 = n2861 & n35244 ;
  assign n29012 = n23311 | n23324 ;
  assign n29013 = n894 & n35465 ;
  assign n29014 = n29012 | n29013 ;
  assign n29015 = n24199 | n29014 ;
  assign n36949 = ~n29015 ;
  assign n29016 = x29 & n36949 ;
  assign n29017 = n30024 & n29015 ;
  assign n29018 = n29016 | n29017 ;
  assign n29019 = n29011 | n29018 ;
  assign n29020 = n29011 & n29018 ;
  assign n36950 = ~n29020 ;
  assign n29021 = n29019 & n36950 ;
  assign n36951 = ~n28900 ;
  assign n29022 = n28893 & n36951 ;
  assign n29023 = n28903 | n28905 ;
  assign n36952 = ~n29022 ;
  assign n29024 = n36952 & n29023 ;
  assign n29025 = n29021 & n29024 ;
  assign n29026 = n29021 | n29024 ;
  assign n36953 = ~n29025 ;
  assign n29027 = n36953 & n29026 ;
  assign n25297 = n3791 & n25288 ;
  assign n24075 = n3802 & n24057 ;
  assign n24098 = n209 & n24080 ;
  assign n29028 = n24075 | n24098 ;
  assign n29029 = n3818 & n24676 ;
  assign n29030 = n29028 | n29029 ;
  assign n29031 = n25297 | n29030 ;
  assign n36954 = ~n29031 ;
  assign n29032 = x26 & n36954 ;
  assign n29033 = n30019 & n29031 ;
  assign n29034 = n29032 | n29033 ;
  assign n29035 = n29027 | n29034 ;
  assign n29036 = n29027 & n29034 ;
  assign n36955 = ~n29036 ;
  assign n29037 = n29035 & n36955 ;
  assign n29038 = n28915 & n28917 ;
  assign n36956 = ~n28908 ;
  assign n29039 = n36956 & n28920 ;
  assign n29040 = n29038 | n29039 ;
  assign n36957 = ~n29040 ;
  assign n29041 = n29037 & n36957 ;
  assign n36958 = ~n29037 ;
  assign n29042 = n36958 & n29040 ;
  assign n29043 = n29041 | n29042 ;
  assign n25429 = n4135 & n35785 ;
  assign n24829 = n4148 & n24815 ;
  assign n24858 = n4185 & n35663 ;
  assign n29044 = n24829 | n24858 ;
  assign n29045 = n4165 & n35784 ;
  assign n29046 = n29044 | n29045 ;
  assign n29047 = n25429 | n29046 ;
  assign n36959 = ~n29047 ;
  assign n29048 = x23 & n36959 ;
  assign n29049 = n30030 & n29047 ;
  assign n29050 = n29048 | n29049 ;
  assign n29051 = n29043 | n29050 ;
  assign n29052 = n29043 & n29050 ;
  assign n36960 = ~n29052 ;
  assign n29053 = n29051 & n36960 ;
  assign n29054 = n28933 | n28934 ;
  assign n36961 = ~n28931 ;
  assign n29055 = n36961 & n29054 ;
  assign n29056 = n29053 & n29055 ;
  assign n29057 = n29053 | n29055 ;
  assign n36962 = ~n29056 ;
  assign n29058 = n36962 & n29057 ;
  assign n26286 = n4686 & n26284 ;
  assign n25812 = n4726 & n25796 ;
  assign n26054 = n4706 & n26039 ;
  assign n29059 = n25812 | n26054 ;
  assign n29060 = n4748 & n26278 ;
  assign n29061 = n29059 | n29060 ;
  assign n29062 = n26286 | n29061 ;
  assign n36963 = ~n29062 ;
  assign n29063 = x20 & n36963 ;
  assign n29064 = n30374 & n29062 ;
  assign n29065 = n29063 | n29064 ;
  assign n29066 = n29058 | n29065 ;
  assign n29067 = n29058 & n29065 ;
  assign n36964 = ~n29067 ;
  assign n29068 = n29066 & n36964 ;
  assign n29069 = n5164 | n26279 ;
  assign n29070 = n30580 & n29069 ;
  assign n29071 = x16 | n29069 ;
  assign n36965 = ~n29070 ;
  assign n29072 = n36965 & n29071 ;
  assign n29073 = n28947 | n28950 ;
  assign n36966 = ~n28945 ;
  assign n29074 = n36966 & n29073 ;
  assign n36967 = ~n29072 ;
  assign n29075 = n36967 & n29074 ;
  assign n36968 = ~n29074 ;
  assign n29076 = n29072 & n36968 ;
  assign n29077 = n29075 | n29076 ;
  assign n29078 = n29068 & n29077 ;
  assign n29080 = n29068 | n29077 ;
  assign n36969 = ~n29078 ;
  assign n29081 = n36969 & n29080 ;
  assign n36970 = ~n28953 ;
  assign n28966 = n36970 & n28964 ;
  assign n29082 = n28960 & n28961 ;
  assign n29083 = n28966 | n29082 ;
  assign n29084 = n29081 | n29083 ;
  assign n29085 = n29081 & n29083 ;
  assign n36971 = ~n29085 ;
  assign n29086 = n29084 & n36971 ;
  assign n29087 = n28856 | n28860 ;
  assign n29088 = n36937 & n29087 ;
  assign n29089 = n28972 | n29088 ;
  assign n36972 = ~n28971 ;
  assign n29090 = n36972 & n29089 ;
  assign n29091 = n29086 & n29090 ;
  assign n29092 = n29086 | n29090 ;
  assign n36973 = ~n29091 ;
  assign n29093 = n36973 & n29092 ;
  assign n36974 = ~n28981 ;
  assign n29094 = n36974 & n29093 ;
  assign n36975 = ~n29093 ;
  assign n29095 = n28981 & n36975 ;
  assign n29886 = n29094 | n29095 ;
  assign n29096 = n766 | n797 ;
  assign n29097 = n3967 | n29096 ;
  assign n29098 = n2709 | n29097 ;
  assign n29099 = n630 | n13738 ;
  assign n29100 = n28623 | n29099 ;
  assign n29101 = n29098 | n29100 ;
  assign n29102 = n239 | n668 ;
  assign n29103 = n416 | n475 ;
  assign n29104 = n29102 | n29103 ;
  assign n29105 = n2600 | n29104 ;
  assign n29106 = n4951 | n29105 ;
  assign n29107 = n29101 | n29106 ;
  assign n29108 = n14368 | n29107 ;
  assign n29109 = n389 | n3264 ;
  assign n29110 = n29108 | n29109 ;
  assign n36976 = ~n29110 ;
  assign n29111 = n28997 & n36976 ;
  assign n29112 = n36945 & n29110 ;
  assign n29113 = n29111 | n29112 ;
  assign n29006 = n28998 | n29004 ;
  assign n36977 = ~n28999 ;
  assign n29114 = n36977 & n29006 ;
  assign n29115 = n29113 & n29114 ;
  assign n29116 = n29113 | n29114 ;
  assign n36978 = ~n29115 ;
  assign n29117 = n36978 & n29116 ;
  assign n23406 = n889 & n35252 ;
  assign n22531 = n3311 & n35020 ;
  assign n23353 = n3329 & n23339 ;
  assign n29118 = n22531 | n23353 ;
  assign n29119 = n3343 & n35254 ;
  assign n29120 = n29118 | n29119 ;
  assign n29121 = n23406 | n29120 ;
  assign n29122 = n29117 | n29121 ;
  assign n29123 = n29117 & n29121 ;
  assign n36979 = ~n29123 ;
  assign n29124 = n29122 & n36979 ;
  assign n24178 = n895 & n24168 ;
  assign n23303 = n2861 & n35467 ;
  assign n24124 = n2849 & n35458 ;
  assign n29125 = n23303 | n24124 ;
  assign n29126 = n894 & n24080 ;
  assign n29127 = n29125 | n29126 ;
  assign n29128 = n24178 | n29127 ;
  assign n36980 = ~n29128 ;
  assign n29129 = x29 & n36980 ;
  assign n29130 = n30024 & n29128 ;
  assign n29131 = n29129 | n29130 ;
  assign n36981 = ~n29131 ;
  assign n29132 = n29124 & n36981 ;
  assign n36982 = ~n29124 ;
  assign n29133 = n36982 & n29131 ;
  assign n29134 = n29132 | n29133 ;
  assign n36983 = ~n28982 ;
  assign n29135 = n36983 & n29008 ;
  assign n36984 = ~n29135 ;
  assign n29136 = n29019 & n36984 ;
  assign n36985 = ~n29134 ;
  assign n29137 = n36985 & n29136 ;
  assign n36986 = ~n29136 ;
  assign n29138 = n29134 & n36986 ;
  assign n29139 = n29137 | n29138 ;
  assign n25329 = n3791 & n35670 ;
  assign n24076 = n209 & n24057 ;
  assign n24693 = n3802 & n24676 ;
  assign n29140 = n24076 | n24693 ;
  assign n29141 = n3818 & n35663 ;
  assign n29142 = n29140 | n29141 ;
  assign n29143 = n25329 | n29142 ;
  assign n36987 = ~n29143 ;
  assign n29144 = x26 & n36987 ;
  assign n29145 = n30019 & n29143 ;
  assign n29146 = n29144 | n29145 ;
  assign n36988 = ~n29146 ;
  assign n29147 = n29139 & n36988 ;
  assign n36989 = ~n29139 ;
  assign n29148 = n36989 & n29146 ;
  assign n29149 = n29147 | n29148 ;
  assign n36990 = ~n29024 ;
  assign n29150 = n29021 & n36990 ;
  assign n36991 = ~n29150 ;
  assign n29151 = n29035 & n36991 ;
  assign n36992 = ~n29149 ;
  assign n29152 = n36992 & n29151 ;
  assign n36993 = ~n29151 ;
  assign n29153 = n29149 & n36993 ;
  assign n29154 = n29152 | n29153 ;
  assign n25826 = n4135 & n35910 ;
  assign n24831 = n4185 & n24815 ;
  assign n25409 = n4148 & n35784 ;
  assign n29155 = n24831 | n25409 ;
  assign n29156 = n4165 & n25796 ;
  assign n29157 = n29155 | n29156 ;
  assign n29158 = n25826 | n29157 ;
  assign n36994 = ~n29158 ;
  assign n29159 = x23 & n36994 ;
  assign n29160 = n30030 & n29158 ;
  assign n29161 = n29159 | n29160 ;
  assign n36995 = ~n29161 ;
  assign n29162 = n29154 & n36995 ;
  assign n36996 = ~n29154 ;
  assign n29163 = n36996 & n29161 ;
  assign n29164 = n29162 | n29163 ;
  assign n26495 = n4686 & n36130 ;
  assign n26055 = n4726 & n26039 ;
  assign n26479 = n4706 & n26278 ;
  assign n29165 = n26055 | n26479 ;
  assign n29166 = n4748 & n36131 ;
  assign n29167 = n29165 | n29166 ;
  assign n29168 = n26495 | n29167 ;
  assign n29169 = x20 | n29168 ;
  assign n29170 = x20 & n29168 ;
  assign n36997 = ~n29170 ;
  assign n29171 = n29169 & n36997 ;
  assign n36998 = ~n29041 ;
  assign n29172 = n36998 & n29051 ;
  assign n29173 = n29171 & n29172 ;
  assign n29174 = n29171 | n29172 ;
  assign n36999 = ~n29173 ;
  assign n29175 = n36999 & n29174 ;
  assign n37000 = ~n29164 ;
  assign n29176 = n37000 & n29175 ;
  assign n37001 = ~n29175 ;
  assign n29177 = n29164 & n37001 ;
  assign n29178 = n29176 | n29177 ;
  assign n37002 = ~n29055 ;
  assign n29179 = n29053 & n37002 ;
  assign n37003 = ~n29179 ;
  assign n29180 = n29066 & n37003 ;
  assign n29181 = x17 & n29180 ;
  assign n29182 = x17 | n29180 ;
  assign n37004 = ~n29181 ;
  assign n29183 = n37004 & n29182 ;
  assign n37005 = ~n29178 ;
  assign n29184 = n37005 & n29183 ;
  assign n37006 = ~n29183 ;
  assign n29185 = n29178 & n37006 ;
  assign n29186 = n29184 | n29185 ;
  assign n37007 = ~n29068 ;
  assign n29079 = n37007 & n29077 ;
  assign n29187 = n29072 & n29074 ;
  assign n29188 = n29079 | n29187 ;
  assign n29189 = n29186 | n29188 ;
  assign n29190 = n29186 & n29188 ;
  assign n37008 = ~n29190 ;
  assign n29191 = n29189 & n37008 ;
  assign n37009 = ~n29083 ;
  assign n29192 = n29081 & n37009 ;
  assign n29193 = n36972 & n28978 ;
  assign n29194 = n29086 | n29193 ;
  assign n37010 = ~n29192 ;
  assign n29195 = n37010 & n29194 ;
  assign n37011 = ~n29191 ;
  assign n29196 = n37011 & n29195 ;
  assign n37012 = ~n29195 ;
  assign n29197 = n29191 & n37012 ;
  assign n29198 = n29196 | n29197 ;
  assign n29199 = n29095 | n29198 ;
  assign n29200 = n29095 & n29198 ;
  assign n37013 = ~n29200 ;
  assign n54 = n29199 & n37013 ;
  assign n1995 = n416 | n1994 ;
  assign n29201 = n126 | n412 ;
  assign n29202 = n1995 | n29201 ;
  assign n29203 = n3493 | n20725 ;
  assign n29204 = n29202 | n29203 ;
  assign n29205 = n948 | n2439 ;
  assign n29206 = n29204 | n29205 ;
  assign n29207 = n3670 | n23087 ;
  assign n29208 = n29206 | n29207 ;
  assign n29209 = n3957 | n29208 ;
  assign n29210 = n11255 | n29209 ;
  assign n29211 = n12348 | n29210 ;
  assign n29212 = n29110 | n29211 ;
  assign n29213 = n29110 & n29211 ;
  assign n37014 = ~n29213 ;
  assign n29214 = n29212 & n37014 ;
  assign n29215 = x17 & n29214 ;
  assign n29217 = x17 | n29214 ;
  assign n37015 = ~n29215 ;
  assign n29218 = n37015 & n29217 ;
  assign n23383 = n889 & n23372 ;
  assign n23337 = n3329 & n35244 ;
  assign n23351 = n3311 & n23339 ;
  assign n29219 = n23337 | n23351 ;
  assign n29220 = n3343 & n35246 ;
  assign n29221 = n29219 | n29220 ;
  assign n29222 = n23383 | n29221 ;
  assign n37016 = ~n29222 ;
  assign n29223 = n29218 & n37016 ;
  assign n37017 = ~n29218 ;
  assign n29224 = n37017 & n29222 ;
  assign n29225 = n29223 | n29224 ;
  assign n29226 = n28997 & n29110 ;
  assign n37018 = ~n29114 ;
  assign n29227 = n29113 & n37018 ;
  assign n29228 = n29226 | n29227 ;
  assign n29229 = n29225 | n29228 ;
  assign n29230 = n29225 & n29228 ;
  assign n37019 = ~n29230 ;
  assign n29231 = n29229 & n37019 ;
  assign n37020 = ~n29132 ;
  assign n29232 = n29122 & n37020 ;
  assign n37021 = ~n29231 ;
  assign n29233 = n37021 & n29232 ;
  assign n37022 = ~n29232 ;
  assign n29234 = n29231 & n37022 ;
  assign n29235 = n29233 | n29234 ;
  assign n24147 = n895 & n35457 ;
  assign n24088 = n2849 & n24080 ;
  assign n24113 = n2861 & n35458 ;
  assign n29236 = n24088 | n24113 ;
  assign n29237 = n894 & n24151 ;
  assign n29238 = n29236 | n29237 ;
  assign n29239 = n24147 | n29238 ;
  assign n37023 = ~n29239 ;
  assign n29240 = x29 & n37023 ;
  assign n29241 = n30024 & n29239 ;
  assign n29242 = n29240 | n29241 ;
  assign n37024 = ~n29242 ;
  assign n29243 = n29235 & n37024 ;
  assign n37025 = ~n29235 ;
  assign n29244 = n37025 & n29242 ;
  assign n29245 = n29243 | n29244 ;
  assign n24883 = n3791 & n35662 ;
  assign n24680 = n209 & n24676 ;
  assign n24851 = n3802 & n35663 ;
  assign n29246 = n24680 | n24851 ;
  assign n29247 = n3818 & n24815 ;
  assign n29248 = n29246 | n29247 ;
  assign n29249 = n24883 | n29248 ;
  assign n37026 = ~n29249 ;
  assign n29250 = x26 & n37026 ;
  assign n29251 = n30019 & n29249 ;
  assign n29252 = n29250 | n29251 ;
  assign n29253 = n29245 | n29252 ;
  assign n29254 = n29245 & n29252 ;
  assign n37027 = ~n29254 ;
  assign n29255 = n29253 & n37027 ;
  assign n29256 = n29134 | n29136 ;
  assign n37028 = ~n29147 ;
  assign n29257 = n37028 & n29256 ;
  assign n29258 = n29255 & n29257 ;
  assign n29259 = n29255 | n29257 ;
  assign n37029 = ~n29258 ;
  assign n29260 = n37029 & n29259 ;
  assign n26074 = n4135 & n26065 ;
  assign n25411 = n4185 & n35784 ;
  assign n25811 = n4148 & n25796 ;
  assign n29261 = n25411 | n25811 ;
  assign n29262 = n4165 & n26039 ;
  assign n29263 = n29261 | n29262 ;
  assign n29264 = n26074 | n29263 ;
  assign n37030 = ~n29264 ;
  assign n29265 = x23 & n37030 ;
  assign n29266 = n30030 & n29264 ;
  assign n29267 = n29265 | n29266 ;
  assign n29268 = n29260 | n29267 ;
  assign n29269 = n29260 & n29267 ;
  assign n37031 = ~n29269 ;
  assign n29270 = n29268 & n37031 ;
  assign n29271 = n29149 | n29151 ;
  assign n37032 = ~n29162 ;
  assign n29272 = n37032 & n29271 ;
  assign n29273 = n29270 & n29272 ;
  assign n29274 = n29270 | n29272 ;
  assign n37033 = ~n29273 ;
  assign n29275 = n37033 & n29274 ;
  assign n26704 = n4686 & n36192 ;
  assign n29276 = n4726 & n26278 ;
  assign n29277 = n4706 & n36131 ;
  assign n29278 = n29276 | n29277 ;
  assign n29279 = n26704 | n29278 ;
  assign n37034 = ~n29279 ;
  assign n29280 = x20 & n37034 ;
  assign n29281 = n30374 & n29279 ;
  assign n29282 = n29280 | n29281 ;
  assign n29283 = n29164 & n29175 ;
  assign n29284 = n29173 | n29283 ;
  assign n29285 = n29282 | n29284 ;
  assign n29286 = n29282 & n29284 ;
  assign n37035 = ~n29286 ;
  assign n29287 = n29285 & n37035 ;
  assign n37036 = ~n29275 ;
  assign n29288 = n37036 & n29287 ;
  assign n37037 = ~n29287 ;
  assign n29289 = n29275 & n37037 ;
  assign n29290 = n29288 | n29289 ;
  assign n37038 = ~n29184 ;
  assign n29291 = n29182 & n37038 ;
  assign n37039 = ~n29290 ;
  assign n29292 = n37039 & n29291 ;
  assign n37040 = ~n29291 ;
  assign n29293 = n29290 & n37040 ;
  assign n29294 = n29292 | n29293 ;
  assign n29295 = n29092 & n37010 ;
  assign n37041 = ~n29295 ;
  assign n29296 = n29191 & n37041 ;
  assign n37042 = ~n29296 ;
  assign n29297 = n29189 & n37042 ;
  assign n37043 = ~n29294 ;
  assign n29298 = n37043 & n29297 ;
  assign n37044 = ~n29297 ;
  assign n29299 = n29294 & n37044 ;
  assign n29300 = n29298 | n29299 ;
  assign n29301 = n29200 | n29300 ;
  assign n29302 = n29200 & n29300 ;
  assign n37045 = ~n29302 ;
  assign n55 = n29301 & n37045 ;
  assign n29216 = n30580 & n29214 ;
  assign n29303 = n29213 | n29216 ;
  assign n29304 = n811 | n814 ;
  assign n29305 = n1091 | n29304 ;
  assign n29306 = n185 | n292 ;
  assign n29307 = n29305 | n29306 ;
  assign n29308 = n1853 | n23897 ;
  assign n29309 = n29307 | n29308 ;
  assign n29310 = n1483 | n2288 ;
  assign n29311 = n2893 | n11246 ;
  assign n29312 = n29310 | n29311 ;
  assign n29313 = n2613 | n29312 ;
  assign n29314 = n29309 | n29313 ;
  assign n29315 = n2684 | n4594 ;
  assign n29316 = n29314 | n29315 ;
  assign n37046 = ~n29316 ;
  assign n29317 = n27904 & n37046 ;
  assign n29318 = n34916 & n29317 ;
  assign n37047 = ~n29303 ;
  assign n29319 = n37047 & n29318 ;
  assign n37048 = ~n29318 ;
  assign n29320 = n29303 & n37048 ;
  assign n29321 = n29319 | n29320 ;
  assign n24202 = n889 & n35472 ;
  assign n23298 = n3329 & n35467 ;
  assign n23325 = n3311 & n35244 ;
  assign n29322 = n23298 | n23325 ;
  assign n29323 = n3343 & n35465 ;
  assign n29324 = n29322 | n29323 ;
  assign n29325 = n24202 | n29324 ;
  assign n37049 = ~n29325 ;
  assign n29326 = n29321 & n37049 ;
  assign n37050 = ~n29321 ;
  assign n29327 = n37050 & n29325 ;
  assign n29328 = n29326 | n29327 ;
  assign n37051 = ~n29225 ;
  assign n29329 = n37051 & n29228 ;
  assign n29330 = n29223 | n29329 ;
  assign n37052 = ~n29330 ;
  assign n29331 = n29328 & n37052 ;
  assign n37053 = ~n29328 ;
  assign n29332 = n37053 & n29330 ;
  assign n29333 = n29331 | n29332 ;
  assign n25299 = n895 & n25288 ;
  assign n24059 = n2849 & n24057 ;
  assign n24099 = n2861 & n24080 ;
  assign n29334 = n24059 | n24099 ;
  assign n29335 = n894 & n24676 ;
  assign n29336 = n29334 | n29335 ;
  assign n29337 = n25299 | n29336 ;
  assign n37054 = ~n29337 ;
  assign n29338 = x29 & n37054 ;
  assign n29339 = n30024 & n29337 ;
  assign n29340 = n29338 | n29339 ;
  assign n29341 = n29333 | n29340 ;
  assign n29342 = n29333 & n29340 ;
  assign n37055 = ~n29342 ;
  assign n29343 = n29341 & n37055 ;
  assign n29344 = n29231 | n29232 ;
  assign n37056 = ~n29243 ;
  assign n29345 = n37056 & n29344 ;
  assign n29346 = n29343 & n29345 ;
  assign n29347 = n29343 | n29345 ;
  assign n37057 = ~n29346 ;
  assign n29348 = n37057 & n29347 ;
  assign n25430 = n3791 & n35785 ;
  assign n24830 = n3802 & n24815 ;
  assign n24855 = n209 & n35663 ;
  assign n29349 = n24830 | n24855 ;
  assign n29350 = n3818 & n35784 ;
  assign n29351 = n29349 | n29350 ;
  assign n29352 = n25430 | n29351 ;
  assign n37058 = ~n29352 ;
  assign n29353 = x26 & n37058 ;
  assign n29354 = n30019 & n29352 ;
  assign n29355 = n29353 | n29354 ;
  assign n29356 = n29348 | n29355 ;
  assign n29357 = n29348 & n29355 ;
  assign n37059 = ~n29357 ;
  assign n29358 = n29356 & n37059 ;
  assign n37060 = ~n29257 ;
  assign n29359 = n29255 & n37060 ;
  assign n37061 = ~n29359 ;
  assign n29360 = n29253 & n37061 ;
  assign n29361 = n29358 & n29360 ;
  assign n29362 = n29358 | n29360 ;
  assign n37062 = ~n29361 ;
  assign n29363 = n37062 & n29362 ;
  assign n26294 = n4135 & n26284 ;
  assign n25809 = n4185 & n25796 ;
  assign n26056 = n4148 & n26039 ;
  assign n29364 = n25809 | n26056 ;
  assign n29365 = n4165 & n26278 ;
  assign n29366 = n29364 | n29365 ;
  assign n29367 = n26294 | n29366 ;
  assign n37063 = ~n29367 ;
  assign n29368 = x23 & n37063 ;
  assign n29369 = n30030 & n29367 ;
  assign n29370 = n29368 | n29369 ;
  assign n29371 = n29363 | n29370 ;
  assign n29372 = n29363 & n29370 ;
  assign n37064 = ~n29372 ;
  assign n29373 = n29371 & n37064 ;
  assign n29374 = n4724 | n26279 ;
  assign n29375 = n30374 & n29374 ;
  assign n29376 = x19 | n29374 ;
  assign n37065 = ~n29375 ;
  assign n29377 = n37065 & n29376 ;
  assign n37066 = ~n29272 ;
  assign n29378 = n29270 & n37066 ;
  assign n37067 = ~n29378 ;
  assign n29379 = n29268 & n37067 ;
  assign n37068 = ~n29377 ;
  assign n29380 = n37068 & n29379 ;
  assign n37069 = ~n29379 ;
  assign n29381 = n29377 & n37069 ;
  assign n29382 = n29380 | n29381 ;
  assign n29383 = n29373 & n29382 ;
  assign n29385 = n29373 | n29382 ;
  assign n37070 = ~n29383 ;
  assign n29386 = n37070 & n29385 ;
  assign n37071 = ~n29288 ;
  assign n29387 = n29285 & n37071 ;
  assign n37072 = ~n29386 ;
  assign n29388 = n37072 & n29387 ;
  assign n37073 = ~n29387 ;
  assign n29389 = n29386 & n37073 ;
  assign n29390 = n29388 | n29389 ;
  assign n29391 = n29290 | n29291 ;
  assign n37074 = ~n29197 ;
  assign n29392 = n29189 & n37074 ;
  assign n37075 = ~n29392 ;
  assign n29393 = n29294 & n37075 ;
  assign n37076 = ~n29393 ;
  assign n29394 = n29391 & n37076 ;
  assign n29395 = n29390 & n29394 ;
  assign n29396 = n29390 | n29394 ;
  assign n37077 = ~n29395 ;
  assign n29397 = n37077 & n29396 ;
  assign n29398 = n37045 & n29397 ;
  assign n37078 = ~n29397 ;
  assign n29399 = n29302 & n37078 ;
  assign n29883 = n29398 | n29399 ;
  assign n29400 = n29303 & n29318 ;
  assign n29401 = n29321 & n29325 ;
  assign n29402 = n29400 | n29401 ;
  assign n29403 = n3906 | n21514 ;
  assign n29404 = n23110 | n29403 ;
  assign n29405 = n217 | n528 ;
  assign n29406 = n2244 | n29405 ;
  assign n29407 = n2396 | n29406 ;
  assign n29408 = n29099 | n29407 ;
  assign n29409 = n29404 | n29408 ;
  assign n29410 = n12340 | n27254 ;
  assign n29411 = n29409 | n29410 ;
  assign n37079 = ~n29411 ;
  assign n29412 = n11737 & n37079 ;
  assign n37080 = ~n5388 ;
  assign n29413 = n37080 & n29412 ;
  assign n37081 = ~n3978 ;
  assign n29414 = n37081 & n29413 ;
  assign n37082 = ~n29414 ;
  assign n29415 = n29318 & n37082 ;
  assign n29416 = n37048 & n29414 ;
  assign n29417 = n29415 | n29416 ;
  assign n24179 = n889 & n24168 ;
  assign n23312 = n3311 & n35467 ;
  assign n24125 = n3329 & n35458 ;
  assign n29418 = n23312 | n24125 ;
  assign n29419 = n3343 & n24080 ;
  assign n29420 = n29418 | n29419 ;
  assign n29421 = n24179 | n29420 ;
  assign n37083 = ~n29421 ;
  assign n29422 = n29417 & n37083 ;
  assign n37084 = ~n29417 ;
  assign n29424 = n37084 & n29421 ;
  assign n29425 = n29422 | n29424 ;
  assign n29426 = n29402 | n29425 ;
  assign n29427 = n29402 & n29425 ;
  assign n37085 = ~n29427 ;
  assign n29428 = n29426 & n37085 ;
  assign n37086 = ~n29332 ;
  assign n29429 = n37086 & n29341 ;
  assign n37087 = ~n29428 ;
  assign n29430 = n37087 & n29429 ;
  assign n37088 = ~n29429 ;
  assign n29431 = n29428 & n37088 ;
  assign n29432 = n29430 | n29431 ;
  assign n25322 = n895 & n35670 ;
  assign n24073 = n2861 & n24057 ;
  assign n24697 = n2849 & n24676 ;
  assign n29433 = n24073 | n24697 ;
  assign n29434 = n894 & n35663 ;
  assign n29435 = n29433 | n29434 ;
  assign n29436 = n25322 | n29435 ;
  assign n29437 = x29 | n29436 ;
  assign n29438 = x29 & n29436 ;
  assign n37089 = ~n29438 ;
  assign n29439 = n29437 & n37089 ;
  assign n29440 = n29432 & n29439 ;
  assign n29441 = n29432 | n29439 ;
  assign n37090 = ~n29440 ;
  assign n29442 = n37090 & n29441 ;
  assign n25834 = n3791 & n35910 ;
  assign n24832 = n209 & n24815 ;
  assign n25401 = n3802 & n35784 ;
  assign n29443 = n24832 | n25401 ;
  assign n29444 = n3818 & n25796 ;
  assign n29445 = n29443 | n29444 ;
  assign n29446 = n25834 | n29445 ;
  assign n37091 = ~n29446 ;
  assign n29447 = x26 & n37091 ;
  assign n29448 = n30019 & n29446 ;
  assign n29449 = n29447 | n29448 ;
  assign n29450 = n29442 | n29449 ;
  assign n29451 = n29442 & n29449 ;
  assign n37092 = ~n29451 ;
  assign n29452 = n29450 & n37092 ;
  assign n26496 = n4135 & n36130 ;
  assign n26047 = n4185 & n26039 ;
  assign n26480 = n4148 & n26278 ;
  assign n29453 = n26047 | n26480 ;
  assign n29454 = n4165 & n36131 ;
  assign n29455 = n29453 | n29454 ;
  assign n29456 = n26496 | n29455 ;
  assign n29457 = x23 | n29456 ;
  assign n29458 = x23 & n29456 ;
  assign n37093 = ~n29458 ;
  assign n29459 = n29457 & n37093 ;
  assign n37094 = ~n29345 ;
  assign n29460 = n29343 & n37094 ;
  assign n37095 = ~n29460 ;
  assign n29461 = n29356 & n37095 ;
  assign n29462 = n29459 & n29461 ;
  assign n29463 = n29459 | n29461 ;
  assign n37096 = ~n29462 ;
  assign n29464 = n37096 & n29463 ;
  assign n37097 = ~n29452 ;
  assign n29465 = n37097 & n29464 ;
  assign n37098 = ~n29464 ;
  assign n29467 = n29452 & n37098 ;
  assign n29468 = n29465 | n29467 ;
  assign n37099 = ~n29360 ;
  assign n29469 = n29358 & n37099 ;
  assign n37100 = ~n29469 ;
  assign n29470 = n29371 & n37100 ;
  assign n29471 = x20 & n29470 ;
  assign n29472 = x20 | n29470 ;
  assign n37101 = ~n29471 ;
  assign n29473 = n37101 & n29472 ;
  assign n29474 = n29468 & n29473 ;
  assign n29475 = n29468 | n29473 ;
  assign n37102 = ~n29474 ;
  assign n29476 = n37102 & n29475 ;
  assign n37103 = ~n29373 ;
  assign n29384 = n37103 & n29382 ;
  assign n29477 = n29377 & n29379 ;
  assign n29478 = n29384 | n29477 ;
  assign n29479 = n29476 | n29478 ;
  assign n29480 = n29476 & n29478 ;
  assign n37104 = ~n29480 ;
  assign n29481 = n29479 & n37104 ;
  assign n37105 = ~n29299 ;
  assign n29482 = n37105 & n29391 ;
  assign n29483 = n29390 | n29482 ;
  assign n37106 = ~n29389 ;
  assign n29484 = n37106 & n29483 ;
  assign n29485 = n29481 & n29484 ;
  assign n29486 = n29481 | n29484 ;
  assign n37107 = ~n29485 ;
  assign n29487 = n37107 & n29486 ;
  assign n37108 = ~n29399 ;
  assign n29488 = n37108 & n29487 ;
  assign n37109 = ~n29487 ;
  assign n29489 = n29399 & n37109 ;
  assign n29882 = n29488 | n29489 ;
  assign n37110 = ~n29402 ;
  assign n29490 = n37110 & n29425 ;
  assign n29491 = n29428 | n29429 ;
  assign n37111 = ~n29490 ;
  assign n29492 = n37111 & n29491 ;
  assign n29493 = n151 | n187 ;
  assign n29494 = n495 | n29493 ;
  assign n29495 = n2659 | n22226 ;
  assign n29496 = n29494 | n29495 ;
  assign n29497 = n1878 | n2503 ;
  assign n29498 = n29496 | n29497 ;
  assign n29499 = n2709 | n29498 ;
  assign n29500 = n2974 | n3197 ;
  assign n29501 = n3484 | n3997 ;
  assign n29502 = n29500 | n29501 ;
  assign n29503 = n754 | n29502 ;
  assign n37112 = ~n29503 ;
  assign n29504 = n13717 & n37112 ;
  assign n37113 = ~n29499 ;
  assign n29505 = n37113 & n29504 ;
  assign n37114 = ~n3733 ;
  assign n29506 = n37114 & n29505 ;
  assign n37115 = ~n11115 ;
  assign n29507 = n37115 & n29506 ;
  assign n29508 = n29318 & n29507 ;
  assign n29509 = n29318 | n29507 ;
  assign n37116 = ~n29508 ;
  assign n29510 = n37116 & n29509 ;
  assign n29511 = x20 & n29510 ;
  assign n29513 = x20 | n29510 ;
  assign n37117 = ~n29511 ;
  assign n29514 = n37117 & n29513 ;
  assign n29423 = n29415 | n29421 ;
  assign n37118 = ~n29416 ;
  assign n29515 = n37118 & n29423 ;
  assign n37119 = ~n29514 ;
  assign n29516 = n37119 & n29515 ;
  assign n37120 = ~n29515 ;
  assign n29517 = n29514 & n37120 ;
  assign n29518 = n29516 | n29517 ;
  assign n24141 = n889 & n35457 ;
  assign n24100 = n3329 & n24080 ;
  assign n24109 = n3311 & n35458 ;
  assign n29519 = n24100 | n24109 ;
  assign n29520 = n3343 & n24151 ;
  assign n29521 = n29519 | n29520 ;
  assign n29522 = n24141 | n29521 ;
  assign n29523 = n29518 | n29522 ;
  assign n29525 = n29518 & n29522 ;
  assign n37121 = ~n29525 ;
  assign n29526 = n29523 & n37121 ;
  assign n37122 = ~n29526 ;
  assign n29527 = n29492 & n37122 ;
  assign n37123 = ~n29492 ;
  assign n29528 = n37123 & n29526 ;
  assign n29529 = n29527 | n29528 ;
  assign n24878 = n895 & n35662 ;
  assign n24691 = n2861 & n24676 ;
  assign n24852 = n2849 & n35663 ;
  assign n29530 = n24691 | n24852 ;
  assign n29531 = n894 & n24815 ;
  assign n29532 = n29530 | n29531 ;
  assign n29533 = n24878 | n29532 ;
  assign n37124 = ~n29533 ;
  assign n29534 = x29 & n37124 ;
  assign n29535 = n30024 & n29533 ;
  assign n29536 = n29534 | n29535 ;
  assign n29537 = n29529 | n29536 ;
  assign n29538 = n29529 & n29536 ;
  assign n37125 = ~n29538 ;
  assign n29539 = n29537 & n37125 ;
  assign n26075 = n3791 & n26065 ;
  assign n25412 = n209 & n35784 ;
  assign n25813 = n3802 & n25796 ;
  assign n29540 = n25412 | n25813 ;
  assign n29541 = n3818 & n26039 ;
  assign n29542 = n29540 | n29541 ;
  assign n29543 = n26075 | n29542 ;
  assign n29544 = x26 | n29543 ;
  assign n29545 = x26 & n29543 ;
  assign n37126 = ~n29545 ;
  assign n29546 = n29544 & n37126 ;
  assign n37127 = ~n29432 ;
  assign n29547 = n37127 & n29439 ;
  assign n37128 = ~n29442 ;
  assign n29548 = n37128 & n29449 ;
  assign n29549 = n29547 | n29548 ;
  assign n37129 = ~n29549 ;
  assign n29550 = n29546 & n37129 ;
  assign n37130 = ~n29546 ;
  assign n29551 = n37130 & n29549 ;
  assign n29552 = n29550 | n29551 ;
  assign n37131 = ~n29539 ;
  assign n29553 = n37131 & n29552 ;
  assign n37132 = ~n29552 ;
  assign n29555 = n29539 & n37132 ;
  assign n29556 = n29553 | n29555 ;
  assign n26701 = n4135 & n36192 ;
  assign n29557 = n4185 & n26278 ;
  assign n29558 = n4148 & n36131 ;
  assign n29559 = n29557 | n29558 ;
  assign n29560 = n26701 | n29559 ;
  assign n37133 = ~n29560 ;
  assign n29561 = x23 & n37133 ;
  assign n29562 = n30030 & n29560 ;
  assign n29563 = n29561 | n29562 ;
  assign n37134 = ~n29563 ;
  assign n29564 = n29556 & n37134 ;
  assign n37135 = ~n29556 ;
  assign n29565 = n37135 & n29563 ;
  assign n29566 = n29564 | n29565 ;
  assign n29466 = n29452 & n29464 ;
  assign n37136 = ~n29466 ;
  assign n29567 = n29463 & n37136 ;
  assign n37137 = ~n29566 ;
  assign n29568 = n37137 & n29567 ;
  assign n37138 = ~n29567 ;
  assign n29569 = n29566 & n37138 ;
  assign n29570 = n29568 | n29569 ;
  assign n37139 = ~n29468 ;
  assign n29571 = n37139 & n29473 ;
  assign n29572 = n29471 | n29571 ;
  assign n37140 = ~n29572 ;
  assign n29573 = n29570 & n37140 ;
  assign n37141 = ~n29570 ;
  assign n29574 = n37141 & n29572 ;
  assign n29575 = n29573 | n29574 ;
  assign n37142 = ~n29478 ;
  assign n29576 = n29476 & n37142 ;
  assign n29577 = n37106 & n29396 ;
  assign n29578 = n29481 | n29577 ;
  assign n37143 = ~n29576 ;
  assign n29579 = n37143 & n29578 ;
  assign n29580 = n29575 & n29579 ;
  assign n29581 = n29575 | n29579 ;
  assign n37144 = ~n29580 ;
  assign n29582 = n37144 & n29581 ;
  assign n37145 = ~n29489 ;
  assign n29583 = n37145 & n29582 ;
  assign n37146 = ~n29582 ;
  assign n29584 = n29489 & n37146 ;
  assign n29881 = n29583 | n29584 ;
  assign n29512 = n30374 & n29510 ;
  assign n37147 = ~n29512 ;
  assign n29585 = n29509 & n37147 ;
  assign n29586 = n474 | n1537 ;
  assign n29587 = n1625 | n29586 ;
  assign n29588 = n4294 | n13506 ;
  assign n29589 = n29587 | n29588 ;
  assign n29590 = n1759 | n23176 ;
  assign n29591 = n29589 | n29590 ;
  assign n29592 = n1481 | n13565 ;
  assign n29593 = n29591 | n29592 ;
  assign n29594 = n578 | n1579 ;
  assign n29595 = n12821 | n29594 ;
  assign n29596 = n29593 | n29595 ;
  assign n29597 = n12348 | n29596 ;
  assign n29598 = n29585 & n29597 ;
  assign n29599 = n29585 | n29597 ;
  assign n37148 = ~n29598 ;
  assign n29600 = n37148 & n29599 ;
  assign n25298 = n889 & n25288 ;
  assign n24077 = n3329 & n24057 ;
  assign n24101 = n3311 & n24080 ;
  assign n29601 = n24077 | n24101 ;
  assign n29602 = n3343 & n24676 ;
  assign n29603 = n29601 | n29602 ;
  assign n29604 = n25298 | n29603 ;
  assign n37149 = ~n29604 ;
  assign n29605 = n29600 & n37149 ;
  assign n37150 = ~n29600 ;
  assign n29606 = n37150 & n29604 ;
  assign n29607 = n29605 | n29606 ;
  assign n29524 = n29516 | n29522 ;
  assign n37151 = ~n29517 ;
  assign n29608 = n37151 & n29524 ;
  assign n29609 = n29607 & n29608 ;
  assign n29610 = n29607 | n29608 ;
  assign n37152 = ~n29609 ;
  assign n29611 = n37152 & n29610 ;
  assign n25431 = n895 & n35785 ;
  assign n24833 = n2849 & n24815 ;
  assign n24857 = n2861 & n35663 ;
  assign n29612 = n24833 | n24857 ;
  assign n29613 = n894 & n35784 ;
  assign n29614 = n29612 | n29613 ;
  assign n29615 = n25431 | n29614 ;
  assign n37153 = ~n29615 ;
  assign n29616 = x29 & n37153 ;
  assign n29617 = n30024 & n29615 ;
  assign n29618 = n29616 | n29617 ;
  assign n37154 = ~n29618 ;
  assign n29619 = n29611 & n37154 ;
  assign n37155 = ~n29611 ;
  assign n29620 = n37155 & n29618 ;
  assign n29621 = n29619 | n29620 ;
  assign n37156 = ~n29529 ;
  assign n29622 = n37156 & n29536 ;
  assign n29623 = n29527 | n29622 ;
  assign n29624 = n29621 | n29623 ;
  assign n29625 = n29621 & n29623 ;
  assign n37157 = ~n29625 ;
  assign n29626 = n29624 & n37157 ;
  assign n26293 = n3791 & n26284 ;
  assign n25815 = n209 & n25796 ;
  assign n26050 = n3802 & n26039 ;
  assign n29627 = n25815 | n26050 ;
  assign n29628 = n3818 & n26278 ;
  assign n29629 = n29627 | n29628 ;
  assign n29630 = n26293 | n29629 ;
  assign n37158 = ~n29630 ;
  assign n29631 = x26 & n37158 ;
  assign n29632 = n30019 & n29630 ;
  assign n29633 = n29631 | n29632 ;
  assign n37159 = ~n29633 ;
  assign n29634 = n29626 & n37159 ;
  assign n37160 = ~n29626 ;
  assign n29635 = n37160 & n29633 ;
  assign n29636 = n29634 | n29635 ;
  assign n29637 = n4183 | n26279 ;
  assign n29638 = n30030 & n29637 ;
  assign n29639 = x22 | n29637 ;
  assign n37161 = ~n29638 ;
  assign n29640 = n37161 & n29639 ;
  assign n29554 = n29539 & n29552 ;
  assign n29641 = n29546 | n29549 ;
  assign n37162 = ~n29554 ;
  assign n29642 = n37162 & n29641 ;
  assign n37163 = ~n29640 ;
  assign n29643 = n37163 & n29642 ;
  assign n37164 = ~n29642 ;
  assign n29644 = n29640 & n37164 ;
  assign n29645 = n29643 | n29644 ;
  assign n37165 = ~n29636 ;
  assign n29646 = n37165 & n29645 ;
  assign n37166 = ~n29645 ;
  assign n29647 = n29636 & n37166 ;
  assign n29648 = n29646 | n29647 ;
  assign n29649 = n29566 | n29567 ;
  assign n37167 = ~n29564 ;
  assign n29650 = n37167 & n29649 ;
  assign n29651 = n29648 & n29650 ;
  assign n29652 = n29648 | n29650 ;
  assign n37168 = ~n29651 ;
  assign n29653 = n37168 & n29652 ;
  assign n29654 = n29486 & n37143 ;
  assign n29655 = n29575 | n29654 ;
  assign n37169 = ~n29573 ;
  assign n29656 = n37169 & n29655 ;
  assign n37170 = ~n29653 ;
  assign n29657 = n37170 & n29656 ;
  assign n37171 = ~n29656 ;
  assign n29658 = n29653 & n37171 ;
  assign n29659 = n29657 | n29658 ;
  assign n29660 = n29584 | n29659 ;
  assign n29661 = n29584 & n29659 ;
  assign n37172 = ~n29661 ;
  assign n59 = n29660 & n37172 ;
  assign n37173 = ~n29634 ;
  assign n29662 = n29624 & n37173 ;
  assign n29663 = x23 & n29662 ;
  assign n29664 = x23 | n29662 ;
  assign n37174 = ~n29663 ;
  assign n29665 = n37174 & n29664 ;
  assign n29666 = n486 | n827 ;
  assign n29667 = n233 | n29666 ;
  assign n29668 = n514 | n29667 ;
  assign n29669 = n1126 | n23896 ;
  assign n29670 = n29668 | n29669 ;
  assign n29671 = n237 | n347 ;
  assign n29672 = n751 | n4652 ;
  assign n29673 = n29671 | n29672 ;
  assign n29674 = n13435 | n29673 ;
  assign n29675 = n29670 | n29674 ;
  assign n29676 = n24703 | n27917 ;
  assign n29677 = n29675 | n29676 ;
  assign n37175 = ~n29677 ;
  assign n29678 = n20247 & n37175 ;
  assign n29679 = n32659 & n29678 ;
  assign n29681 = n29597 | n29679 ;
  assign n29682 = n29597 & n29679 ;
  assign n37176 = ~n29682 ;
  assign n29683 = n29681 & n37176 ;
  assign n29684 = n29600 & n29604 ;
  assign n37177 = ~n29684 ;
  assign n29685 = n29599 & n37177 ;
  assign n29686 = n29683 & n29685 ;
  assign n29687 = n29683 | n29685 ;
  assign n37178 = ~n29686 ;
  assign n29688 = n37178 & n29687 ;
  assign n25328 = n889 & n35670 ;
  assign n24078 = n3311 & n24057 ;
  assign n24681 = n3329 & n24676 ;
  assign n29689 = n24078 | n24681 ;
  assign n29690 = n3343 & n35663 ;
  assign n29691 = n29689 | n29690 ;
  assign n29692 = n25328 | n29691 ;
  assign n29693 = n29688 | n29692 ;
  assign n29694 = n29688 & n29692 ;
  assign n37179 = ~n29694 ;
  assign n29695 = n29693 & n37179 ;
  assign n37180 = ~n29619 ;
  assign n29696 = n29610 & n37180 ;
  assign n37181 = ~n29695 ;
  assign n29697 = n37181 & n29696 ;
  assign n37182 = ~n29696 ;
  assign n29698 = n29695 & n37182 ;
  assign n29699 = n29697 | n29698 ;
  assign n25832 = n895 & n35910 ;
  assign n24835 = n2861 & n24815 ;
  assign n25407 = n2849 & n35784 ;
  assign n29700 = n24835 | n25407 ;
  assign n29701 = n894 & n25796 ;
  assign n29702 = n29700 | n29701 ;
  assign n29703 = n25832 | n29702 ;
  assign n29704 = x29 | n29703 ;
  assign n29705 = x29 & n29703 ;
  assign n37183 = ~n29705 ;
  assign n29706 = n29704 & n37183 ;
  assign n29707 = n29699 & n29706 ;
  assign n29708 = n29699 | n29706 ;
  assign n37184 = ~n29707 ;
  assign n29709 = n37184 & n29708 ;
  assign n26488 = n3791 & n36130 ;
  assign n26057 = n209 & n26039 ;
  assign n26481 = n3802 & n26278 ;
  assign n29710 = n26057 | n26481 ;
  assign n29711 = n3818 & n36131 ;
  assign n29712 = n29710 | n29711 ;
  assign n29713 = n26488 | n29712 ;
  assign n37185 = ~n29713 ;
  assign n29714 = x26 & n37185 ;
  assign n29715 = n30019 & n29713 ;
  assign n29716 = n29714 | n29715 ;
  assign n29717 = n29709 | n29716 ;
  assign n29718 = n29709 & n29716 ;
  assign n37186 = ~n29718 ;
  assign n29719 = n29717 & n37186 ;
  assign n29720 = n29665 & n29719 ;
  assign n29721 = n29665 | n29719 ;
  assign n37187 = ~n29720 ;
  assign n29722 = n37187 & n29721 ;
  assign n29723 = n29640 & n29642 ;
  assign n29724 = n29636 & n29645 ;
  assign n29725 = n29723 | n29724 ;
  assign n29726 = n29722 | n29725 ;
  assign n29727 = n29722 & n29725 ;
  assign n37188 = ~n29727 ;
  assign n29728 = n29726 & n37188 ;
  assign n29729 = n37169 & n29581 ;
  assign n29730 = n29651 | n29729 ;
  assign n29731 = n29652 & n29730 ;
  assign n29732 = n29728 & n29731 ;
  assign n29733 = n29728 | n29731 ;
  assign n37189 = ~n29732 ;
  assign n29734 = n37189 & n29733 ;
  assign n29735 = n37172 & n29734 ;
  assign n37190 = ~n29734 ;
  assign n29736 = n29661 & n37190 ;
  assign n29879 = n29735 | n29736 ;
  assign n29680 = x23 & n29679 ;
  assign n29737 = x23 | n29679 ;
  assign n37191 = ~n29680 ;
  assign n29738 = n37191 & n29737 ;
  assign n29739 = n1435 | n3022 ;
  assign n29740 = n4918 | n29739 ;
  assign n29741 = n276 | n380 ;
  assign n29742 = n930 | n29741 ;
  assign n29743 = n5901 | n29742 ;
  assign n29744 = n29740 | n29743 ;
  assign n29745 = n1366 | n11214 ;
  assign n29746 = n13415 | n29745 ;
  assign n29747 = n29744 | n29746 ;
  assign n37192 = ~n29747 ;
  assign n29748 = n5814 & n37192 ;
  assign n37193 = ~n14993 ;
  assign n29749 = n37193 & n29748 ;
  assign n29750 = n29738 & n29749 ;
  assign n29751 = n29738 | n29749 ;
  assign n37194 = ~n29750 ;
  assign n29752 = n37194 & n29751 ;
  assign n37195 = ~n29685 ;
  assign n29753 = n29681 & n37195 ;
  assign n29754 = n29682 | n29753 ;
  assign n37196 = ~n29752 ;
  assign n29755 = n37196 & n29754 ;
  assign n37197 = ~n29754 ;
  assign n29756 = n29752 & n37197 ;
  assign n29757 = n29755 | n29756 ;
  assign n24884 = n889 & n35662 ;
  assign n24698 = n3311 & n24676 ;
  assign n24842 = n3329 & n35663 ;
  assign n29758 = n24698 | n24842 ;
  assign n29759 = n3343 & n24815 ;
  assign n29760 = n29758 | n29759 ;
  assign n29761 = n24884 | n29760 ;
  assign n29762 = n29757 | n29761 ;
  assign n29763 = n29757 & n29761 ;
  assign n37198 = ~n29763 ;
  assign n29764 = n29762 & n37198 ;
  assign n26076 = n895 & n26065 ;
  assign n25397 = n2861 & n35784 ;
  assign n25816 = n2849 & n25796 ;
  assign n29765 = n25397 | n25816 ;
  assign n29766 = n894 & n26039 ;
  assign n29767 = n29765 | n29766 ;
  assign n29768 = n26076 | n29767 ;
  assign n37199 = ~n29768 ;
  assign n29769 = x29 & n37199 ;
  assign n29770 = n30024 & n29768 ;
  assign n29771 = n29769 | n29770 ;
  assign n37200 = ~n29771 ;
  assign n29772 = n29764 & n37200 ;
  assign n37201 = ~n29764 ;
  assign n29773 = n37201 & n29771 ;
  assign n29774 = n29772 | n29773 ;
  assign n37202 = ~n29692 ;
  assign n29775 = n29688 & n37202 ;
  assign n29776 = n29695 | n29696 ;
  assign n37203 = ~n29775 ;
  assign n29777 = n37203 & n29776 ;
  assign n37204 = ~n29774 ;
  assign n29778 = n37204 & n29777 ;
  assign n37205 = ~n29777 ;
  assign n29779 = n29774 & n37205 ;
  assign n29780 = n29778 | n29779 ;
  assign n26702 = n3791 & n36192 ;
  assign n29781 = n209 & n26278 ;
  assign n29782 = n3802 & n36131 ;
  assign n29783 = n29781 | n29782 ;
  assign n29784 = n26702 | n29783 ;
  assign n29785 = x26 | n29784 ;
  assign n29786 = x26 & n29784 ;
  assign n37206 = ~n29786 ;
  assign n29787 = n29785 & n37206 ;
  assign n37207 = ~n29706 ;
  assign n29788 = n29699 & n37207 ;
  assign n37208 = ~n29788 ;
  assign n29789 = n29717 & n37208 ;
  assign n29790 = n29787 & n29789 ;
  assign n29791 = n29787 | n29789 ;
  assign n37209 = ~n29790 ;
  assign n29792 = n37209 & n29791 ;
  assign n37210 = ~n29780 ;
  assign n29793 = n37210 & n29792 ;
  assign n37211 = ~n29792 ;
  assign n29794 = n29780 & n37211 ;
  assign n29795 = n29793 | n29794 ;
  assign n37212 = ~n29719 ;
  assign n29796 = n29665 & n37212 ;
  assign n29797 = n29663 | n29796 ;
  assign n37213 = ~n29795 ;
  assign n29798 = n37213 & n29797 ;
  assign n37214 = ~n29797 ;
  assign n29799 = n29795 & n37214 ;
  assign n29800 = n29798 | n29799 ;
  assign n37215 = ~n29725 ;
  assign n29801 = n29722 & n37215 ;
  assign n29802 = n29651 | n29656 ;
  assign n29803 = n29652 & n29802 ;
  assign n29804 = n29728 | n29803 ;
  assign n37216 = ~n29801 ;
  assign n29805 = n37216 & n29804 ;
  assign n29806 = n29800 & n29805 ;
  assign n29807 = n29800 | n29805 ;
  assign n37217 = ~n29806 ;
  assign n29808 = n37217 & n29807 ;
  assign n37218 = ~n29736 ;
  assign n29809 = n37218 & n29808 ;
  assign n37219 = ~n29808 ;
  assign n29810 = n29736 & n37219 ;
  assign n29878 = n29809 | n29810 ;
  assign n37220 = ~n29756 ;
  assign n29811 = n37220 & n29762 ;
  assign n29812 = n912 | n1712 ;
  assign n29813 = n2954 | n29812 ;
  assign n29814 = n171 | n187 ;
  assign n29815 = n332 | n29814 ;
  assign n29816 = n250 | n594 ;
  assign n29817 = n29815 | n29816 ;
  assign n29818 = n29813 | n29817 ;
  assign n29819 = n686 | n5438 ;
  assign n29820 = n29818 | n29819 ;
  assign n29821 = n785 | n1067 ;
  assign n29822 = n2524 | n29821 ;
  assign n29823 = n5804 | n29822 ;
  assign n29824 = n29820 | n29823 ;
  assign n29825 = n4903 | n29824 ;
  assign n29826 = n13426 | n29825 ;
  assign n29827 = n25349 | n29826 ;
  assign n37221 = ~n29749 ;
  assign n29828 = n29738 & n37221 ;
  assign n37222 = ~n29828 ;
  assign n29829 = n29737 & n37222 ;
  assign n29830 = n29827 & n29829 ;
  assign n29831 = n29827 | n29829 ;
  assign n37223 = ~n29830 ;
  assign n29832 = n37223 & n29831 ;
  assign n25432 = n889 & n35785 ;
  assign n24834 = n3329 & n24815 ;
  assign n24859 = n3311 & n35663 ;
  assign n29833 = n24834 | n24859 ;
  assign n29834 = n3343 & n35784 ;
  assign n29835 = n29833 | n29834 ;
  assign n29836 = n25432 | n29835 ;
  assign n29837 = n29832 | n29836 ;
  assign n29839 = n29832 & n29836 ;
  assign n37224 = ~n29839 ;
  assign n29840 = n29837 & n37224 ;
  assign n29841 = n29811 & n29840 ;
  assign n29842 = n29811 | n29840 ;
  assign n37225 = ~n29841 ;
  assign n29843 = n37225 & n29842 ;
  assign n26291 = n895 & n26284 ;
  assign n25817 = n2861 & n25796 ;
  assign n26058 = n2849 & n26039 ;
  assign n29844 = n25817 | n26058 ;
  assign n29845 = n894 & n26278 ;
  assign n29846 = n29844 | n29845 ;
  assign n29847 = n26291 | n29846 ;
  assign n37226 = ~n29847 ;
  assign n29848 = x29 & n37226 ;
  assign n29849 = n30024 & n29847 ;
  assign n29850 = n29848 | n29849 ;
  assign n37227 = ~n29850 ;
  assign n29851 = n29843 & n37227 ;
  assign n37228 = ~n29843 ;
  assign n29852 = n37228 & n29850 ;
  assign n29853 = n29851 | n29852 ;
  assign n29854 = n209 & n36131 ;
  assign n29855 = x26 & n29854 ;
  assign n29856 = x26 | n29854 ;
  assign n37229 = ~n29855 ;
  assign n29857 = n37229 & n29856 ;
  assign n29858 = n29774 | n29777 ;
  assign n37230 = ~n29772 ;
  assign n29859 = n37230 & n29858 ;
  assign n29860 = n29857 & n29859 ;
  assign n29861 = n29857 | n29859 ;
  assign n37231 = ~n29860 ;
  assign n29862 = n37231 & n29861 ;
  assign n37232 = ~n29853 ;
  assign n29863 = n37232 & n29862 ;
  assign n37233 = ~n29862 ;
  assign n29864 = n29853 & n37233 ;
  assign n29865 = n29863 | n29864 ;
  assign n29866 = n29790 | n29793 ;
  assign n37234 = ~n29866 ;
  assign n29867 = n29865 & n37234 ;
  assign n37235 = ~n29865 ;
  assign n29868 = n37235 & n29866 ;
  assign n29869 = n29867 | n29868 ;
  assign n29870 = n29798 | n29805 ;
  assign n37236 = ~n29799 ;
  assign n29871 = n37236 & n29870 ;
  assign n37237 = ~n29871 ;
  assign n29872 = n29869 & n37237 ;
  assign n37238 = ~n29869 ;
  assign n29873 = n37238 & n29871 ;
  assign n29874 = n29872 | n29873 ;
  assign n37239 = ~n29874 ;
  assign n29875 = n29810 & n37239 ;
  assign n37240 = ~n29810 ;
  assign n29876 = n37240 & n29874 ;
  assign n62 = n29875 | n29876 ;
  assign n29987 = n29853 & n29862 ;
  assign n29988 = n29860 | n29987 ;
  assign n26494 = n895 & n36130 ;
  assign n26044 = n2861 & n26039 ;
  assign n26483 = n2849 & n26278 ;
  assign n29943 = n26044 | n26483 ;
  assign n29944 = n894 & n36131 ;
  assign n29945 = n29943 | n29944 ;
  assign n29946 = n26494 | n29945 ;
  assign n29947 = x29 | n29946 ;
  assign n29948 = x29 & n29946 ;
  assign n37241 = ~n29948 ;
  assign n29949 = n29947 & n37241 ;
  assign n29951 = n30019 & n29949 ;
  assign n37242 = ~n29949 ;
  assign n29952 = x26 & n37242 ;
  assign n29953 = n29951 | n29952 ;
  assign n37243 = ~n15209 ;
  assign n29912 = n5767 & n37243 ;
  assign n37244 = ~n2166 ;
  assign n29913 = n37244 & n29912 ;
  assign n29914 = n5820 | n5894 ;
  assign n37245 = ~n29914 ;
  assign n29915 = n29913 & n37245 ;
  assign n37246 = ~n5835 ;
  assign n29916 = n37246 & n29915 ;
  assign n29917 = n29827 | n29916 ;
  assign n29918 = n29826 & n29916 ;
  assign n37247 = ~n29918 ;
  assign n29919 = n29917 & n37247 ;
  assign n37248 = ~n29836 ;
  assign n29838 = n29831 & n37248 ;
  assign n29920 = n29830 | n29838 ;
  assign n37249 = ~n29920 ;
  assign n29921 = n29919 & n37249 ;
  assign n37250 = ~n29919 ;
  assign n29923 = n37250 & n29920 ;
  assign n29924 = n29921 | n29923 ;
  assign n25835 = n889 & n35910 ;
  assign n24836 = n3311 & n24815 ;
  assign n25414 = n3329 & n35784 ;
  assign n29925 = n24836 | n25414 ;
  assign n29926 = n3343 & n25796 ;
  assign n29927 = n29925 | n29926 ;
  assign n29928 = n25835 | n29927 ;
  assign n37251 = ~n29928 ;
  assign n29929 = n29924 & n37251 ;
  assign n37252 = ~n29924 ;
  assign n29930 = n37252 & n29928 ;
  assign n29931 = n29929 | n29930 ;
  assign n37253 = ~n29851 ;
  assign n29932 = n29842 & n37253 ;
  assign n37254 = ~n29931 ;
  assign n29933 = n37254 & n29932 ;
  assign n37255 = ~n29932 ;
  assign n29954 = n29931 & n37255 ;
  assign n29955 = n29933 | n29954 ;
  assign n29956 = n29953 | n29955 ;
  assign n29989 = n29953 & n29955 ;
  assign n37256 = ~n29989 ;
  assign n29990 = n29956 & n37256 ;
  assign n37257 = ~n29990 ;
  assign n29991 = n29988 & n37257 ;
  assign n37258 = ~n29988 ;
  assign n29994 = n37258 & n29990 ;
  assign n30003 = n29991 | n29994 ;
  assign n29981 = n29810 & n29874 ;
  assign n29982 = n29865 & n29866 ;
  assign n37259 = ~n29982 ;
  assign n29983 = n29981 & n37259 ;
  assign n29985 = n29869 & n29871 ;
  assign n29986 = n29982 | n29985 ;
  assign n37260 = ~n29981 ;
  assign n30008 = n37260 & n29986 ;
  assign n30009 = n29983 | n30008 ;
  assign n37261 = ~n30003 ;
  assign n30010 = n37261 & n30009 ;
  assign n37262 = ~n30009 ;
  assign n30011 = n30003 & n37262 ;
  assign n30012 = n30010 | n30011 ;
  assign n29993 = n29981 | n29986 ;
  assign n37263 = ~n29994 ;
  assign n29995 = n29993 & n37263 ;
  assign n29984 = n29981 & n29982 ;
  assign n29934 = n29930 | n29933 ;
  assign n26482 = n2861 & n26278 ;
  assign n26705 = n895 & n36192 ;
  assign n29935 = n26482 | n26705 ;
  assign n29922 = n29918 | n29920 ;
  assign n29936 = n29917 & n29922 ;
  assign n37264 = ~n29935 ;
  assign n29937 = n37264 & n29936 ;
  assign n37265 = ~n29936 ;
  assign n29938 = n29935 & n37265 ;
  assign n29939 = n29937 | n29938 ;
  assign n37266 = ~n29934 ;
  assign n29940 = n37266 & n29939 ;
  assign n37267 = ~n29939 ;
  assign n29941 = n29934 & n37267 ;
  assign n29942 = n29940 | n29941 ;
  assign n29950 = x26 & n29949 ;
  assign n37268 = ~n29955 ;
  assign n29957 = n29953 & n37268 ;
  assign n29958 = n29950 | n29957 ;
  assign n29959 = n5788 | n5909 ;
  assign n37293 = x26 & x29 ;
  assign n29960 = x26 | x29 ;
  assign n37269 = ~n37293 ;
  assign n29961 = n37269 & n29960 ;
  assign n29962 = n29827 & n29961 ;
  assign n29963 = n29827 | n29961 ;
  assign n37270 = ~n29962 ;
  assign n29964 = n37270 & n29963 ;
  assign n29965 = n29959 & n29964 ;
  assign n29966 = n29959 | n29964 ;
  assign n37271 = ~n29965 ;
  assign n29967 = n37271 & n29966 ;
  assign n26069 = n889 & n26065 ;
  assign n25413 = n3311 & n35784 ;
  assign n25814 = n3329 & n25796 ;
  assign n29968 = n25413 | n25814 ;
  assign n29969 = n3343 & n26039 ;
  assign n29970 = n29968 | n29969 ;
  assign n29971 = n26069 | n29970 ;
  assign n37272 = ~n29971 ;
  assign n29972 = n29967 & n37272 ;
  assign n37273 = ~n29967 ;
  assign n29973 = n37273 & n29971 ;
  assign n29974 = n29972 | n29973 ;
  assign n37274 = ~n29974 ;
  assign n29975 = n29958 & n37274 ;
  assign n37275 = ~n29958 ;
  assign n29976 = n37275 & n29974 ;
  assign n29977 = n29975 | n29976 ;
  assign n37276 = ~n29977 ;
  assign n29978 = n29942 & n37276 ;
  assign n37277 = ~n29942 ;
  assign n29979 = n37277 & n29977 ;
  assign n29980 = n29978 | n29979 ;
  assign n37278 = ~n29991 ;
  assign n29996 = n29980 & n37278 ;
  assign n37279 = ~n29984 ;
  assign n29997 = n37279 & n29996 ;
  assign n37280 = ~n29995 ;
  assign n29998 = n37280 & n29997 ;
  assign n37281 = ~n29980 ;
  assign n29992 = n37281 & n29991 ;
  assign n29999 = n29992 | n29996 ;
  assign n37282 = ~n29999 ;
  assign n30000 = n29984 & n37282 ;
  assign n30001 = n29998 | n30000 ;
  assign n30002 = n37279 & n29991 ;
  assign n30004 = n29993 & n37261 ;
  assign n30005 = n30002 | n30004 ;
  assign n30006 = n37281 & n30005 ;
  assign n64 = n30001 | n30006 ;
  assign n35 = ~n29909 ;
  assign n36 = ~n29908 ;
  assign n37 = ~n29907 ;
  assign n38 = ~n29905 ;
  assign n39 = ~n29904 ;
  assign n40 = ~n29902 ;
  assign n45 = ~n29895 ;
  assign n46 = ~n29894 ;
  assign n47 = ~n29893 ;
  assign n49 = ~n29891 ;
  assign n51 = ~n29889 ;
  assign n52 = ~n29887 ;
  assign n53 = ~n29886 ;
  assign n56 = ~n29883 ;
  assign n57 = ~n29882 ;
  assign n58 = ~n29881 ;
  assign n60 = ~n29879 ;
  assign n61 = ~n29878 ;
  assign n63 = ~n30012 ;
  assign y0 = n33 ;
  assign y1 = n34 ;
  assign y2 = n35 ;
  assign y3 = n36 ;
  assign y4 = n37 ;
  assign y5 = n38 ;
  assign y6 = n39 ;
  assign y7 = n40 ;
  assign y8 = n41 ;
  assign y9 = n42 ;
  assign y10 = n43 ;
  assign y11 = n44 ;
  assign y12 = n45 ;
  assign y13 = n46 ;
  assign y14 = n47 ;
  assign y15 = n48 ;
  assign y16 = n49 ;
  assign y17 = n50 ;
  assign y18 = n51 ;
  assign y19 = n52 ;
  assign y20 = n53 ;
  assign y21 = n54 ;
  assign y22 = n55 ;
  assign y23 = n56 ;
  assign y24 = n57 ;
  assign y25 = n58 ;
  assign y26 = n59 ;
  assign y27 = n60 ;
  assign y28 = n61 ;
  assign y29 = n62 ;
  assign y30 = n63 ;
  assign y31 = n64 ;
endmodule
