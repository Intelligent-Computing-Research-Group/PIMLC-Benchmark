module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 ;
  assign n16 = x27 & x28 ;
  assign n106 = x29 & n16 ;
  assign n165 = x23 & x24 ;
  assign n175 = x25 & n165 ;
  assign n107 = x21 | x22 ;
  assign n108 = x16 | x18 ;
  assign n109 = x12 | x13 ;
  assign n110 = n108 | n109 ;
  assign n111 = x9 | x10 ;
  assign n112 = x11 & n111 ;
  assign n113 = n110 | n112 ;
  assign n175 = x14 & x15 ;
  assign n114 = n175 | n108 ;
  assign n18 = x19 & x20 ;
  assign n115 = x17 | x18 ;
  assign n116 = n18 & n115 ;
  assign n117 = n114 & n116 ;
  assign n118 = n113 & n117 ;
  assign n119 = n107 | n118 ;
  assign n120 = n175 & n119 ;
  assign n121 = x26 | n120 ;
  assign n122 = n106 & n121 ;
  assign n123 = x3 | x4 ;
  assign n124 = x5 | x6 ;
  assign n125 = n123 | n124 ;
  assign n126 = x1 | x2 ;
  assign n127 = n107 | n126 ;
  assign n128 = n125 | n127 ;
  assign n129 = x7 | x8 ;
  assign n130 = x10 | x26 ;
  assign n131 = n129 | n130 ;
  assign n132 = n110 | n131 ;
  assign n133 = n128 | n132 ;
  assign n134 = n122 & n133 ;
  assign n174 = x0 & x1 ;
  assign n20 = x2 & x3 ;
  assign n135 = n174 & n20 ;
  assign n136 = n175 & n18 ;
  assign n137 = n135 & n136 ;
  assign n175 = x8 & x11 ;
  assign n138 = x17 & n175 ;
  assign n22 = x4 & x5 ;
  assign n175 = x6 & x7 ;
  assign n139 = n22 & n175 ;
  assign n140 = n138 & n139 ;
  assign n141 = n175 & n106 ;
  assign n142 = n140 & n141 ;
  assign n143 = n137 & n142 ;
  assign n145 = n122 | n143 ;
  assign n170 = ~n134 ;
  assign n146 = n170 & n145 ;
  assign n175 = x49 & x50 ;
  assign n175 = x44 & x45 ;
  assign n175 = x46 | n175 ;
  assign n26 = x47 & n175 ;
  assign n175 = x48 | n26 ;
  assign n28 = n175 & n175 ;
  assign n12 = x33 & x34 ;
  assign n175 = x35 & x36 ;
  assign n97 = n12 & n175 ;
  assign n14 = x31 & x32 ;
  assign n171 = ~x0 ;
  assign n98 = n171 & x30 ;
  assign n99 = n14 & n98 ;
  assign n100 = n97 & n99 ;
  assign n175 = x57 & x58 ;
  assign n175 = x59 & n175 ;
  assign n90 = x37 & x38 ;
  assign n175 = x41 & n90 ;
  assign n10 = x53 & x54 ;
  assign n175 = x55 & n10 ;
  assign n101 = n175 & n175 ;
  assign n102 = n175 & n101 ;
  assign n103 = n100 & n102 ;
  assign n104 = n28 & n103 ;
  assign n30 = x56 | n175 ;
  assign n32 = n30 & n175 ;
  assign n149 = x51 | x52 ;
  assign n150 = x56 | n149 ;
  assign n152 = x39 | x40 ;
  assign n153 = x41 & n152 ;
  assign n24 = x46 | x48 ;
  assign n154 = x42 | x43 ;
  assign n155 = n24 | n154 ;
  assign n156 = n153 | n155 ;
  assign n157 = n28 & n156 ;
  assign n158 = n150 | n157 ;
  assign n159 = n32 & n158 ;
  assign n160 = n104 | n159 ;
  assign n105 = x0 | x30 ;
  assign n175 = x31 | x32 ;
  assign n91 = x33 | x34 ;
  assign n92 = x35 | x36 ;
  assign n93 = n91 | n92 ;
  assign n94 = n175 | n93 ;
  assign n95 = x37 | x38 ;
  assign n96 = x40 | n95 ;
  assign n151 = n96 | n150 ;
  assign n161 = n151 | n155 ;
  assign n162 = n94 | n161 ;
  assign n166 = n105 | n162 ;
  assign n167 = n145 & n166 ;
  assign n168 = n160 & n167 ;
  assign n169 = n134 | n168 ;
  assign n172 = ~n122 ;
  assign n144 = n172 & n143 ;
  assign n173 = ~n133 ;
  assign n147 = n122 & n173 ;
  assign n148 = n144 | n147 ;
  assign n8 = x0 & x30 ;
  assign n163 = n8 | n162 ;
  assign n164 = n159 & n163 ;
  assign n63 = n148 & n164 ;
  assign n61 = ~n146 ;
  assign n62 = ~n169 ;
  assign y0 = n61 ;
  assign y1 = n62 ;
  assign y2 = n63 ;
endmodule
