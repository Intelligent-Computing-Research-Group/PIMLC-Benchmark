module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 ;
  assign n305 = x0 & x32 ;
  assign n200 = x0 | x32 ;
  assign n314 = ~n305 ;
  assign n65 = n314 & n200 ;
  assign n309 = x1 & x33 ;
  assign n126 = x1 | x33 ;
  assign n315 = ~n309 ;
  assign n202 = n315 & n126 ;
  assign n203 = n314 & n202 ;
  assign n316 = ~n202 ;
  assign n204 = n305 & n316 ;
  assign n66 = n203 | n204 ;
  assign n127 = n305 | n309 ;
  assign n128 = n126 & n127 ;
  assign n241 = x2 & x34 ;
  assign n125 = x2 | x34 ;
  assign n317 = ~n241 ;
  assign n206 = n317 & n125 ;
  assign n207 = n128 & n206 ;
  assign n208 = n128 | n206 ;
  assign n318 = ~n207 ;
  assign n67 = n318 & n208 ;
  assign n129 = n125 & n128 ;
  assign n130 = n241 | n129 ;
  assign n301 = x3 & x35 ;
  assign n124 = x3 | x35 ;
  assign n319 = ~n301 ;
  assign n210 = n319 & n124 ;
  assign n211 = n130 | n210 ;
  assign n212 = n130 & n210 ;
  assign n320 = ~n212 ;
  assign n68 = n211 & n320 ;
  assign n131 = n301 | n130 ;
  assign n132 = n124 & n131 ;
  assign n237 = x4 & x36 ;
  assign n123 = x4 | x36 ;
  assign n321 = ~n237 ;
  assign n214 = n321 & n123 ;
  assign n215 = n132 & n214 ;
  assign n216 = n132 | n214 ;
  assign n322 = ~n215 ;
  assign n69 = n322 & n216 ;
  assign n133 = n123 & n132 ;
  assign n134 = n237 | n133 ;
  assign n297 = x5 & x37 ;
  assign n122 = x5 | x37 ;
  assign n323 = ~n297 ;
  assign n218 = n323 & n122 ;
  assign n324 = ~n134 ;
  assign n219 = n324 & n218 ;
  assign n325 = ~n218 ;
  assign n220 = n134 & n325 ;
  assign n70 = n219 | n220 ;
  assign n135 = n122 & n134 ;
  assign n136 = n297 | n135 ;
  assign n233 = x6 & x38 ;
  assign n121 = x6 | x38 ;
  assign n326 = ~n233 ;
  assign n222 = n326 & n121 ;
  assign n223 = n136 & n222 ;
  assign n224 = n136 | n222 ;
  assign n327 = ~n223 ;
  assign n71 = n327 & n224 ;
  assign n137 = n121 & n136 ;
  assign n138 = n233 | n137 ;
  assign n293 = x7 & x39 ;
  assign n120 = x7 | x39 ;
  assign n328 = ~n293 ;
  assign n226 = n328 & n120 ;
  assign n227 = n138 | n226 ;
  assign n228 = n138 & n226 ;
  assign n329 = ~n228 ;
  assign n72 = n227 & n329 ;
  assign n139 = n120 & n138 ;
  assign n140 = n293 | n139 ;
  assign n229 = x8 & x40 ;
  assign n119 = x8 | x40 ;
  assign n330 = ~n229 ;
  assign n230 = n330 & n119 ;
  assign n231 = n140 & n230 ;
  assign n232 = n140 | n230 ;
  assign n331 = ~n231 ;
  assign n73 = n331 & n232 ;
  assign n141 = n119 & n140 ;
  assign n142 = n229 | n141 ;
  assign n289 = x9 & x41 ;
  assign n118 = x9 | x41 ;
  assign n332 = ~n289 ;
  assign n234 = n332 & n118 ;
  assign n333 = ~n142 ;
  assign n235 = n333 & n234 ;
  assign n334 = ~n234 ;
  assign n236 = n142 & n334 ;
  assign n74 = n235 | n236 ;
  assign n143 = n118 & n142 ;
  assign n144 = n289 | n143 ;
  assign n225 = x10 & x42 ;
  assign n117 = x10 | x42 ;
  assign n335 = ~n225 ;
  assign n238 = n335 & n117 ;
  assign n239 = n144 & n238 ;
  assign n240 = n144 | n238 ;
  assign n336 = ~n239 ;
  assign n75 = n336 & n240 ;
  assign n145 = n117 & n144 ;
  assign n146 = n225 | n145 ;
  assign n285 = x11 & x43 ;
  assign n116 = x11 | x43 ;
  assign n337 = ~n285 ;
  assign n242 = n337 & n116 ;
  assign n243 = n146 | n242 ;
  assign n244 = n146 & n242 ;
  assign n338 = ~n244 ;
  assign n76 = n243 & n338 ;
  assign n147 = n116 & n146 ;
  assign n148 = n285 | n147 ;
  assign n221 = x12 & x44 ;
  assign n115 = x12 | x44 ;
  assign n339 = ~n221 ;
  assign n246 = n339 & n115 ;
  assign n247 = n148 & n246 ;
  assign n248 = n148 | n246 ;
  assign n340 = ~n247 ;
  assign n77 = n340 & n248 ;
  assign n149 = n115 & n148 ;
  assign n150 = n221 | n149 ;
  assign n281 = x13 & x45 ;
  assign n114 = x13 | x45 ;
  assign n341 = ~n281 ;
  assign n250 = n341 & n114 ;
  assign n342 = ~n150 ;
  assign n251 = n342 & n250 ;
  assign n343 = ~n250 ;
  assign n252 = n150 & n343 ;
  assign n78 = n251 | n252 ;
  assign n151 = n114 & n150 ;
  assign n152 = n281 | n151 ;
  assign n217 = x14 & x46 ;
  assign n113 = x14 | x46 ;
  assign n344 = ~n217 ;
  assign n254 = n344 & n113 ;
  assign n255 = n152 & n254 ;
  assign n256 = n152 | n254 ;
  assign n345 = ~n255 ;
  assign n79 = n345 & n256 ;
  assign n153 = n113 & n152 ;
  assign n154 = n217 | n153 ;
  assign n277 = x15 & x47 ;
  assign n112 = x15 | x47 ;
  assign n346 = ~n277 ;
  assign n258 = n346 & n112 ;
  assign n259 = n154 | n258 ;
  assign n260 = n154 & n258 ;
  assign n347 = ~n260 ;
  assign n80 = n259 & n347 ;
  assign n155 = n112 & n154 ;
  assign n156 = n277 | n155 ;
  assign n213 = x16 & x48 ;
  assign n111 = x16 | x48 ;
  assign n348 = ~n213 ;
  assign n262 = n348 & n111 ;
  assign n263 = n156 & n262 ;
  assign n264 = n156 | n262 ;
  assign n349 = ~n263 ;
  assign n81 = n349 & n264 ;
  assign n157 = n111 & n156 ;
  assign n158 = n213 | n157 ;
  assign n273 = x17 & x49 ;
  assign n110 = x17 | x49 ;
  assign n350 = ~n273 ;
  assign n266 = n350 & n110 ;
  assign n351 = ~n158 ;
  assign n267 = n351 & n266 ;
  assign n352 = ~n266 ;
  assign n268 = n158 & n352 ;
  assign n82 = n267 | n268 ;
  assign n159 = n110 & n158 ;
  assign n160 = n273 | n159 ;
  assign n209 = x18 & x50 ;
  assign n109 = x18 | x50 ;
  assign n353 = ~n209 ;
  assign n270 = n353 & n109 ;
  assign n271 = n160 & n270 ;
  assign n272 = n160 | n270 ;
  assign n354 = ~n271 ;
  assign n83 = n354 & n272 ;
  assign n161 = n109 & n160 ;
  assign n162 = n209 | n161 ;
  assign n269 = x19 & x51 ;
  assign n108 = x19 | x51 ;
  assign n355 = ~n269 ;
  assign n274 = n355 & n108 ;
  assign n275 = n162 | n274 ;
  assign n276 = n162 & n274 ;
  assign n356 = ~n276 ;
  assign n84 = n275 & n356 ;
  assign n163 = n108 & n162 ;
  assign n164 = n269 | n163 ;
  assign n205 = x20 & x52 ;
  assign n107 = x20 | x52 ;
  assign n357 = ~n205 ;
  assign n278 = n357 & n107 ;
  assign n279 = n164 & n278 ;
  assign n280 = n164 | n278 ;
  assign n358 = ~n279 ;
  assign n85 = n358 & n280 ;
  assign n165 = n107 & n164 ;
  assign n166 = n205 | n165 ;
  assign n265 = x21 & x53 ;
  assign n106 = x21 | x53 ;
  assign n359 = ~n265 ;
  assign n282 = n359 & n106 ;
  assign n360 = ~n166 ;
  assign n283 = n360 & n282 ;
  assign n361 = ~n282 ;
  assign n284 = n166 & n361 ;
  assign n86 = n283 | n284 ;
  assign n167 = n106 & n166 ;
  assign n168 = n265 | n167 ;
  assign n201 = x22 & x54 ;
  assign n105 = x22 | x54 ;
  assign n362 = ~n201 ;
  assign n286 = n362 & n105 ;
  assign n287 = n168 & n286 ;
  assign n288 = n168 | n286 ;
  assign n363 = ~n287 ;
  assign n87 = n363 & n288 ;
  assign n169 = n105 & n168 ;
  assign n170 = n201 | n169 ;
  assign n261 = x23 & x55 ;
  assign n104 = x23 | x55 ;
  assign n364 = ~n261 ;
  assign n290 = n364 & n104 ;
  assign n291 = n170 | n290 ;
  assign n292 = n170 & n290 ;
  assign n365 = ~n292 ;
  assign n88 = n291 & n365 ;
  assign n171 = n104 & n170 ;
  assign n172 = n261 | n171 ;
  assign n199 = x24 & x56 ;
  assign n103 = x24 | x56 ;
  assign n366 = ~n199 ;
  assign n294 = n366 & n103 ;
  assign n295 = n172 & n294 ;
  assign n296 = n172 | n294 ;
  assign n367 = ~n295 ;
  assign n89 = n367 & n296 ;
  assign n173 = n103 & n172 ;
  assign n174 = n199 | n173 ;
  assign n257 = x25 & x57 ;
  assign n102 = x25 | x57 ;
  assign n368 = ~n257 ;
  assign n298 = n368 & n102 ;
  assign n369 = ~n174 ;
  assign n299 = n369 & n298 ;
  assign n370 = ~n298 ;
  assign n300 = n174 & n370 ;
  assign n90 = n299 | n300 ;
  assign n175 = n102 & n174 ;
  assign n176 = n257 | n175 ;
  assign n192 = x26 & x58 ;
  assign n101 = x26 | x58 ;
  assign n371 = ~n192 ;
  assign n302 = n371 & n101 ;
  assign n372 = ~n302 ;
  assign n303 = n176 & n372 ;
  assign n373 = ~n176 ;
  assign n304 = n373 & n302 ;
  assign n91 = n303 | n304 ;
  assign n177 = n101 & n176 ;
  assign n178 = n192 | n177 ;
  assign n253 = x27 & x59 ;
  assign n100 = x27 | x59 ;
  assign n374 = ~n253 ;
  assign n306 = n374 & n100 ;
  assign n307 = n178 | n306 ;
  assign n308 = n178 & n306 ;
  assign n375 = ~n308 ;
  assign n92 = n307 & n375 ;
  assign n179 = n100 & n178 ;
  assign n180 = n253 | n179 ;
  assign n186 = x28 & x60 ;
  assign n99 = x28 | x60 ;
  assign n376 = ~n186 ;
  assign n310 = n376 & n99 ;
  assign n311 = n180 & n310 ;
  assign n312 = n180 | n310 ;
  assign n377 = ~n311 ;
  assign n93 = n377 & n312 ;
  assign n249 = x29 & x61 ;
  assign n97 = x29 | x61 ;
  assign n378 = ~n249 ;
  assign n98 = n378 & n97 ;
  assign n181 = n99 & n180 ;
  assign n182 = n186 | n181 ;
  assign n183 = n98 | n182 ;
  assign n185 = n98 & n182 ;
  assign n379 = ~n185 ;
  assign n94 = n183 & n379 ;
  assign n245 = x30 & x62 ;
  assign n187 = x30 | x62 ;
  assign n380 = ~n245 ;
  assign n188 = n380 & n187 ;
  assign n184 = n249 | n182 ;
  assign n189 = n97 & n184 ;
  assign n190 = n188 & n189 ;
  assign n191 = n188 | n189 ;
  assign n381 = ~n190 ;
  assign n95 = n381 & n191 ;
  assign n193 = n245 | n189 ;
  assign n194 = n187 & n193 ;
  assign n313 = x31 & x63 ;
  assign n195 = x31 | x63 ;
  assign n382 = ~n313 ;
  assign n196 = n382 & n195 ;
  assign n197 = n194 | n196 ;
  assign n198 = n194 & n196 ;
  assign n383 = ~n198 ;
  assign n96 = n197 & n383 ;
  assign y0 = n65 ;
  assign y1 = n66 ;
  assign y2 = n67 ;
  assign y3 = n68 ;
  assign y4 = n69 ;
  assign y5 = n70 ;
  assign y6 = n71 ;
  assign y7 = n72 ;
  assign y8 = n73 ;
  assign y9 = n74 ;
  assign y10 = n75 ;
  assign y11 = n76 ;
  assign y12 = n77 ;
  assign y13 = n78 ;
  assign y14 = n79 ;
  assign y15 = n80 ;
  assign y16 = n81 ;
  assign y17 = n82 ;
  assign y18 = n83 ;
  assign y19 = n84 ;
  assign y20 = n85 ;
  assign y21 = n86 ;
  assign y22 = n87 ;
  assign y23 = n88 ;
  assign y24 = n89 ;
  assign y25 = n90 ;
  assign y26 = n91 ;
  assign y27 = n92 ;
  assign y28 = n93 ;
  assign y29 = n94 ;
  assign y30 = n95 ;
  assign y31 = n96 ;
endmodule
