module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 ;
  assign n57 = x0 & x8 ;
  assign n25 = x0 | x8 ;
  assign n74 = ~n57 ;
  assign n17 = n74 & n25 ;
  assign n69 = x1 & x9 ;
  assign n32 = x1 | x9 ;
  assign n75 = ~n69 ;
  assign n70 = n75 & n32 ;
  assign n71 = n57 | n70 ;
  assign n72 = n57 & n70 ;
  assign n76 = ~n72 ;
  assign n18 = n71 & n76 ;
  assign n33 = n57 | n69 ;
  assign n34 = n32 & n33 ;
  assign n53 = x2 & x10 ;
  assign n31 = x2 | x10 ;
  assign n77 = ~n53 ;
  assign n66 = n77 & n31 ;
  assign n67 = n34 & n66 ;
  assign n68 = n34 | n66 ;
  assign n78 = ~n67 ;
  assign n19 = n78 & n68 ;
  assign n35 = n53 | n34 ;
  assign n36 = n31 & n35 ;
  assign n65 = x3 & x11 ;
  assign n30 = x3 | x11 ;
  assign n79 = ~n65 ;
  assign n62 = n79 & n30 ;
  assign n63 = n36 | n62 ;
  assign n64 = n36 & n62 ;
  assign n80 = ~n64 ;
  assign n20 = n63 & n80 ;
  assign n37 = n65 | n36 ;
  assign n38 = n30 & n37 ;
  assign n49 = x4 & x12 ;
  assign n29 = x4 | x12 ;
  assign n81 = ~n49 ;
  assign n58 = n81 & n29 ;
  assign n59 = n38 & n58 ;
  assign n60 = n38 | n58 ;
  assign n82 = ~n59 ;
  assign n21 = n82 & n60 ;
  assign n39 = n49 | n38 ;
  assign n40 = n29 & n39 ;
  assign n61 = x5 & x13 ;
  assign n28 = x5 | x13 ;
  assign n83 = ~n61 ;
  assign n54 = n83 & n28 ;
  assign n55 = n40 | n54 ;
  assign n56 = n40 & n54 ;
  assign n84 = ~n56 ;
  assign n22 = n55 & n84 ;
  assign n41 = n61 | n40 ;
  assign n42 = n28 & n41 ;
  assign n26 = x6 & x14 ;
  assign n27 = x6 | x14 ;
  assign n85 = ~n26 ;
  assign n50 = n85 & n27 ;
  assign n51 = n42 & n50 ;
  assign n52 = n42 | n50 ;
  assign n86 = ~n51 ;
  assign n23 = n86 & n52 ;
  assign n43 = n26 | n42 ;
  assign n44 = n27 & n43 ;
  assign n73 = x7 & x15 ;
  assign n45 = x7 | x15 ;
  assign n87 = ~n73 ;
  assign n46 = n87 & n45 ;
  assign n47 = n44 | n46 ;
  assign n48 = n44 & n46 ;
  assign n88 = ~n48 ;
  assign n24 = n47 & n88 ;
  assign y0 = n17 ;
  assign y1 = n18 ;
  assign y2 = n19 ;
  assign y3 = n20 ;
  assign y4 = n21 ;
  assign y5 = n22 ;
  assign y6 = n23 ;
  assign y7 = n24 ;
endmodule
