module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 ;
  assign n18268 = x126 | x127 ;
  assign n18273 = x125 | n18268 ;
  assign n18278 = x124 | n18273 ;
  assign n18283 = x123 | n18278 ;
  assign n18288 = x122 | n18283 ;
  assign n18293 = x121 | n18288 ;
  assign n18298 = x120 | n18293 ;
  assign n18303 = x119 | n18298 ;
  assign n18308 = x118 | n18303 ;
  assign n18313 = x117 | n18308 ;
  assign n18318 = x116 | n18313 ;
  assign n18323 = x115 | n18318 ;
  assign n18328 = x114 | n18323 ;
  assign n18333 = x113 | n18328 ;
  assign n18338 = x112 | n18333 ;
  assign n18343 = x111 | n18338 ;
  assign n18348 = x110 | n18343 ;
  assign n18353 = x109 | n18348 ;
  assign n18357 = x108 | n18353 ;
  assign n18363 = x107 | n18357 ;
  assign n18368 = x106 | n18363 ;
  assign n18373 = x105 | n18368 ;
  assign n18378 = x104 | n18373 ;
  assign n18383 = x103 | n18378 ;
  assign n18388 = x102 | n18383 ;
  assign n18393 = x101 | n18388 ;
  assign n18398 = x100 | n18393 ;
  assign n18403 = x99 | n18398 ;
  assign n18408 = x98 | n18403 ;
  assign n18413 = x97 | n18408 ;
  assign n18418 = x96 | n18413 ;
  assign n18423 = x95 | n18418 ;
  assign n18428 = x94 | n18423 ;
  assign n18433 = x93 | n18428 ;
  assign n18438 = x92 | n18433 ;
  assign n18443 = x91 | n18438 ;
  assign n18448 = x90 | n18443 ;
  assign n18453 = x89 | n18448 ;
  assign n18458 = x88 | n18453 ;
  assign n18463 = x87 | n18458 ;
  assign n18468 = x86 | n18463 ;
  assign n18473 = x85 | n18468 ;
  assign n18478 = x84 | n18473 ;
  assign n18483 = x83 | n18478 ;
  assign n18488 = x82 | n18483 ;
  assign n18493 = x81 | n18488 ;
  assign n18498 = x80 | n18493 ;
  assign n18503 = x79 | n18498 ;
  assign n18508 = x78 | n18503 ;
  assign n18513 = x77 | n18508 ;
  assign n18518 = x76 | n18513 ;
  assign n18523 = x75 | n18518 ;
  assign n18528 = x74 | n18523 ;
  assign n18533 = x73 | n18528 ;
  assign n18538 = x72 | n18533 ;
  assign n18543 = x71 | n18538 ;
  assign n18548 = x70 | n18543 ;
  assign n18553 = x69 | n18548 ;
  assign n18558 = x68 | n18553 ;
  assign n18563 = x67 | n18558 ;
  assign n18579 = ~x62 ;
  assign n18568 = n18579 & x64 ;
  assign n18573 = x65 & n18568 ;
  assign n18263 = x64 | x65 ;
  assign n18580 = ~x66 ;
  assign n18578 = n18580 & n18263 ;
  assign n18581 = ~n18573 ;
  assign n18586 = n18581 & n18578 ;
  assign n18582 = ~n18563 ;
  assign n18594 = n18582 & n18586 ;
  assign n18583 = ~n18594 ;
  assign n18608 = x63 & n18583 ;
  assign n18584 = ~x61 ;
  assign n18772 = n18584 & x64 ;
  assign n18814 = x65 | n18772 ;
  assign n18585 = ~x63 ;
  assign n18622 = n18585 & x65 ;
  assign n18639 = x66 | n18622 ;
  assign n18661 = n18568 | n18639 ;
  assign n18685 = n18563 | n18661 ;
  assign n191 = ~n18685 ;
  assign n18706 = x64 & n191 ;
  assign n18587 = ~n18706 ;
  assign n18736 = x62 & n18587 ;
  assign n18852 = x65 & n18772 ;
  assign n18588 = ~n18852 ;
  assign n18887 = n18736 & n18588 ;
  assign n18589 = ~n18887 ;
  assign n18942 = n18814 & n18589 ;
  assign n18983 = x66 | n18942 ;
  assign n19032 = x66 & n18942 ;
  assign n19096 = n18563 | n19032 ;
  assign n18590 = ~n19096 ;
  assign n19211 = n18983 & n18590 ;
  assign n18591 = ~n19211 ;
  assign n19275 = n18608 & n18591 ;
  assign n18592 = ~x60 ;
  assign n19464 = n18592 & x64 ;
  assign n19614 = x65 | n19464 ;
  assign n19537 = x65 & n19464 ;
  assign n18593 = ~n18608 ;
  assign n19139 = n18593 & n18983 ;
  assign n19696 = n19096 | n19139 ;
  assign n190 = ~n19696 ;
  assign n19773 = x64 & n190 ;
  assign n19882 = x61 & n19773 ;
  assign n19954 = x61 | n19773 ;
  assign n18595 = ~n19882 ;
  assign n20045 = n18595 & n19954 ;
  assign n18596 = ~n19537 ;
  assign n20168 = n18596 & n20045 ;
  assign n18597 = ~n20168 ;
  assign n20260 = n19614 & n18597 ;
  assign n20581 = x66 | n20260 ;
  assign n20388 = x66 & n20260 ;
  assign n20689 = n18814 & n18588 ;
  assign n20799 = n190 & n20689 ;
  assign n18598 = ~n18736 ;
  assign n20950 = n18598 & n20799 ;
  assign n18599 = ~n20799 ;
  assign n21057 = n18736 & n18599 ;
  assign n21217 = n20950 | n21057 ;
  assign n18600 = ~n20388 ;
  assign n21326 = n18600 & n21217 ;
  assign n18601 = ~n21326 ;
  assign n21454 = n20581 & n18601 ;
  assign n18602 = ~n21454 ;
  assign n21583 = n19275 & n18602 ;
  assign n21884 = n18582 & n21583 ;
  assign n18603 = ~x4 ;
  assign n5497 = n18603 & x64 ;
  assign n5498 = x65 | n5497 ;
  assign n18604 = ~x6 ;
  assign n5499 = n18604 & x64 ;
  assign n5501 = x65 | n5499 ;
  assign n5500 = x65 & n5499 ;
  assign n18605 = ~n21583 ;
  assign n21755 = x67 & n18605 ;
  assign n22024 = n18558 | n21755 ;
  assign n18606 = ~n19275 ;
  assign n22164 = n18606 & n21454 ;
  assign n22312 = n22024 | n22164 ;
  assign n20473 = n18580 & n20260 ;
  assign n18607 = ~n20260 ;
  assign n22509 = x66 & n18607 ;
  assign n22639 = n20473 | n22509 ;
  assign n189 = ~n22312 ;
  assign n22843 = n189 & n22639 ;
  assign n18609 = ~n21217 ;
  assign n23035 = n18609 & n22843 ;
  assign n18610 = ~n22843 ;
  assign n23179 = n21217 & n18610 ;
  assign n23395 = n23035 | n23179 ;
  assign n19339 = x68 & n18606 ;
  assign n271 = n18553 | n19339 ;
  assign n18611 = ~x59 ;
  assign n23603 = n18611 & x64 ;
  assign n23991 = x65 | n23603 ;
  assign n23765 = x65 & n23603 ;
  assign n24198 = x64 & n189 ;
  assign n24362 = x60 & n24198 ;
  assign n24600 = x60 | n24198 ;
  assign n18612 = ~n24362 ;
  assign n24822 = n18612 & n24600 ;
  assign n18613 = ~n23765 ;
  assign n24989 = n18613 & n24822 ;
  assign n18614 = ~n24989 ;
  assign n25240 = n23991 & n18614 ;
  assign n257 = x66 | n25240 ;
  assign n25304 = x66 & n25240 ;
  assign n258 = n18596 & n19614 ;
  assign n259 = n189 & n258 ;
  assign n260 = n20045 & n259 ;
  assign n261 = n20045 | n259 ;
  assign n18615 = ~n260 ;
  assign n262 = n18615 & n261 ;
  assign n18616 = ~n25304 ;
  assign n263 = n18616 & n262 ;
  assign n18617 = ~n263 ;
  assign n264 = n257 & n18617 ;
  assign n265 = x67 & n264 ;
  assign n18618 = ~n265 ;
  assign n266 = n23395 & n18618 ;
  assign n267 = n19275 & n22024 ;
  assign n18619 = ~x68 ;
  assign n268 = n18619 & n267 ;
  assign n269 = x67 | n264 ;
  assign n18620 = ~n268 ;
  assign n270 = n18620 & n269 ;
  assign n18621 = ~n266 ;
  assign n272 = n18621 & n270 ;
  assign n273 = n271 | n272 ;
  assign n274 = n18618 & n269 ;
  assign n188 = ~n273 ;
  assign n275 = n188 & n274 ;
  assign n18623 = ~n23395 ;
  assign n276 = n18623 & n275 ;
  assign n18624 = ~n275 ;
  assign n277 = n23395 & n18624 ;
  assign n278 = n276 | n277 ;
  assign n18625 = ~n18553 ;
  assign n279 = n18625 & n267 ;
  assign n280 = n272 & n279 ;
  assign n18626 = ~x58 ;
  assign n281 = n18626 & x64 ;
  assign n282 = x65 | n281 ;
  assign n283 = x65 & n281 ;
  assign n284 = x64 & n188 ;
  assign n285 = x59 & n284 ;
  assign n286 = x59 | n284 ;
  assign n18627 = ~n285 ;
  assign n287 = n18627 & n286 ;
  assign n18628 = ~n283 ;
  assign n288 = n18628 & n287 ;
  assign n18629 = ~n288 ;
  assign n289 = n282 & n18629 ;
  assign n291 = x66 | n289 ;
  assign n290 = x66 & n289 ;
  assign n292 = n18613 & n23991 ;
  assign n293 = n188 & n292 ;
  assign n294 = n24822 & n293 ;
  assign n295 = n24822 | n293 ;
  assign n18630 = ~n294 ;
  assign n296 = n18630 & n295 ;
  assign n18631 = ~n290 ;
  assign n297 = n18631 & n296 ;
  assign n18632 = ~n297 ;
  assign n298 = n291 & n18632 ;
  assign n299 = x67 & n298 ;
  assign n300 = n18616 & n257 ;
  assign n301 = n188 & n300 ;
  assign n302 = n262 & n301 ;
  assign n303 = n262 | n301 ;
  assign n18633 = ~n302 ;
  assign n304 = n18633 & n303 ;
  assign n305 = x67 | n298 ;
  assign n18634 = ~n304 ;
  assign n306 = n18634 & n305 ;
  assign n307 = n299 | n306 ;
  assign n309 = x68 | n307 ;
  assign n18635 = ~n278 ;
  assign n310 = n18635 & n309 ;
  assign n308 = x68 & n307 ;
  assign n18636 = ~n267 ;
  assign n311 = x69 & n18636 ;
  assign n312 = n18548 | n311 ;
  assign n313 = n308 | n312 ;
  assign n314 = n310 | n313 ;
  assign n18637 = ~n280 ;
  assign n315 = n18637 & n314 ;
  assign n18638 = ~n308 ;
  assign n316 = n18638 & n309 ;
  assign n187 = ~n315 ;
  assign n317 = n187 & n316 ;
  assign n318 = n18635 & n317 ;
  assign n18640 = ~n317 ;
  assign n319 = n278 & n18640 ;
  assign n320 = n318 | n319 ;
  assign n18641 = ~x57 ;
  assign n324 = n18641 & x64 ;
  assign n325 = x65 | n324 ;
  assign n326 = x64 & n187 ;
  assign n18642 = ~n326 ;
  assign n327 = x58 & n18642 ;
  assign n328 = n281 & n187 ;
  assign n329 = n327 | n328 ;
  assign n330 = x65 & n324 ;
  assign n18643 = ~n330 ;
  assign n331 = n329 & n18643 ;
  assign n18644 = ~n331 ;
  assign n332 = n325 & n18644 ;
  assign n333 = x66 | n332 ;
  assign n334 = x66 & n332 ;
  assign n335 = n282 & n18628 ;
  assign n336 = n187 & n335 ;
  assign n18645 = ~n336 ;
  assign n337 = n287 & n18645 ;
  assign n18646 = ~n287 ;
  assign n338 = n18646 & n336 ;
  assign n339 = n337 | n338 ;
  assign n18647 = ~n334 ;
  assign n340 = n18647 & n339 ;
  assign n18648 = ~n340 ;
  assign n341 = n333 & n18648 ;
  assign n342 = x67 & n341 ;
  assign n343 = x67 | n341 ;
  assign n344 = n291 & n187 ;
  assign n345 = n297 & n344 ;
  assign n346 = n18631 & n344 ;
  assign n347 = n296 | n346 ;
  assign n18649 = ~n345 ;
  assign n348 = n18649 & n347 ;
  assign n18650 = ~n348 ;
  assign n349 = n343 & n18650 ;
  assign n350 = n342 | n349 ;
  assign n351 = x68 & n350 ;
  assign n352 = x68 | n350 ;
  assign n18651 = ~n299 ;
  assign n353 = n18651 & n305 ;
  assign n354 = n187 & n353 ;
  assign n355 = n304 & n354 ;
  assign n356 = n304 | n354 ;
  assign n18652 = ~n355 ;
  assign n357 = n18652 & n356 ;
  assign n18653 = ~n357 ;
  assign n358 = n352 & n18653 ;
  assign n359 = n351 | n358 ;
  assign n362 = x69 & n359 ;
  assign n18654 = ~n362 ;
  assign n363 = n320 & n18654 ;
  assign n19409 = n18553 & n19275 ;
  assign n321 = n19409 & n314 ;
  assign n322 = n21884 | n321 ;
  assign n18655 = ~x70 ;
  assign n323 = n18655 & n322 ;
  assign n360 = x69 | n359 ;
  assign n18656 = ~n323 ;
  assign n364 = n18656 & n360 ;
  assign n18657 = ~n363 ;
  assign n365 = n18657 & n364 ;
  assign n366 = n18543 | n365 ;
  assign n18658 = ~n322 ;
  assign n367 = x70 & n18658 ;
  assign n368 = n366 | n367 ;
  assign n18659 = ~n359 ;
  assign n361 = x69 & n18659 ;
  assign n18660 = ~x69 ;
  assign n369 = n18660 & n359 ;
  assign n370 = n361 | n369 ;
  assign n186 = ~n368 ;
  assign n371 = n186 & n370 ;
  assign n372 = n320 & n371 ;
  assign n373 = n320 | n371 ;
  assign n18662 = ~n372 ;
  assign n374 = n18662 & n373 ;
  assign n18663 = ~x56 ;
  assign n375 = n18663 & x64 ;
  assign n377 = x65 | n375 ;
  assign n376 = x65 & n375 ;
  assign n378 = x64 & n186 ;
  assign n379 = x57 & n378 ;
  assign n380 = x57 | n378 ;
  assign n18664 = ~n379 ;
  assign n381 = n18664 & n380 ;
  assign n18665 = ~n376 ;
  assign n382 = n18665 & n381 ;
  assign n18666 = ~n382 ;
  assign n383 = n377 & n18666 ;
  assign n384 = x66 & n383 ;
  assign n385 = x66 | n383 ;
  assign n386 = n325 & n186 ;
  assign n388 = n331 & n386 ;
  assign n387 = n18643 & n386 ;
  assign n389 = n329 | n387 ;
  assign n18667 = ~n388 ;
  assign n390 = n18667 & n389 ;
  assign n18668 = ~n390 ;
  assign n391 = n385 & n18668 ;
  assign n392 = n384 | n391 ;
  assign n393 = x67 & n392 ;
  assign n394 = x67 | n392 ;
  assign n395 = n333 & n186 ;
  assign n396 = n340 & n395 ;
  assign n397 = n18647 & n395 ;
  assign n398 = n339 | n397 ;
  assign n18669 = ~n396 ;
  assign n399 = n18669 & n398 ;
  assign n18670 = ~n399 ;
  assign n400 = n394 & n18670 ;
  assign n401 = n393 | n400 ;
  assign n403 = x68 | n401 ;
  assign n402 = x68 & n401 ;
  assign n404 = n342 | n368 ;
  assign n18671 = ~n404 ;
  assign n405 = n343 & n18671 ;
  assign n18672 = ~n405 ;
  assign n406 = n348 & n18672 ;
  assign n407 = n349 & n18671 ;
  assign n408 = n406 | n407 ;
  assign n18673 = ~n402 ;
  assign n409 = n18673 & n408 ;
  assign n18674 = ~n409 ;
  assign n410 = n403 & n18674 ;
  assign n411 = x69 | n410 ;
  assign n412 = x69 & n410 ;
  assign n18675 = ~n351 ;
  assign n413 = n18675 & n352 ;
  assign n414 = n186 & n413 ;
  assign n415 = n18653 & n414 ;
  assign n18676 = ~n414 ;
  assign n416 = n357 & n18676 ;
  assign n417 = n415 | n416 ;
  assign n18677 = ~n412 ;
  assign n418 = n18677 & n417 ;
  assign n18678 = ~n418 ;
  assign n419 = n411 & n18678 ;
  assign n420 = x70 | n419 ;
  assign n421 = x70 & n419 ;
  assign n18679 = ~n421 ;
  assign n422 = n374 & n18679 ;
  assign n18680 = ~n422 ;
  assign n423 = n420 & n18680 ;
  assign n18681 = ~n18538 ;
  assign n424 = n18681 & n322 ;
  assign n18682 = ~n423 ;
  assign n425 = n18682 & n424 ;
  assign n18683 = ~n425 ;
  assign n428 = n18543 & n18683 ;
  assign n426 = n322 & n366 ;
  assign n18684 = ~n426 ;
  assign n429 = n423 & n18684 ;
  assign n430 = n428 | n429 ;
  assign n431 = n420 & n18679 ;
  assign n185 = ~n430 ;
  assign n432 = n185 & n431 ;
  assign n433 = n374 & n432 ;
  assign n434 = n374 | n432 ;
  assign n18686 = ~n433 ;
  assign n435 = n18686 & n434 ;
  assign n18687 = ~x55 ;
  assign n436 = n18687 & x64 ;
  assign n438 = x65 | n436 ;
  assign n437 = x65 & n436 ;
  assign n439 = x64 & n185 ;
  assign n440 = x56 & n439 ;
  assign n441 = x56 | n439 ;
  assign n18688 = ~n440 ;
  assign n442 = n18688 & n441 ;
  assign n18689 = ~n437 ;
  assign n443 = n18689 & n442 ;
  assign n18690 = ~n443 ;
  assign n444 = n438 & n18690 ;
  assign n445 = x66 & n444 ;
  assign n446 = x66 | n444 ;
  assign n447 = n18665 & n377 ;
  assign n448 = n185 & n447 ;
  assign n449 = n381 & n448 ;
  assign n450 = n381 | n448 ;
  assign n18691 = ~n449 ;
  assign n451 = n18691 & n450 ;
  assign n18692 = ~n451 ;
  assign n452 = n446 & n18692 ;
  assign n453 = n445 | n452 ;
  assign n454 = x67 & n453 ;
  assign n455 = x67 | n453 ;
  assign n18693 = ~n384 ;
  assign n456 = n18693 & n385 ;
  assign n457 = n185 & n456 ;
  assign n458 = n390 & n457 ;
  assign n459 = n390 | n457 ;
  assign n18694 = ~n458 ;
  assign n460 = n18694 & n459 ;
  assign n18695 = ~n460 ;
  assign n461 = n455 & n18695 ;
  assign n462 = n454 | n461 ;
  assign n463 = x68 & n462 ;
  assign n464 = x68 | n462 ;
  assign n18696 = ~n393 ;
  assign n465 = n18696 & n394 ;
  assign n466 = n185 & n465 ;
  assign n467 = n18670 & n466 ;
  assign n18697 = ~n466 ;
  assign n468 = n399 & n18697 ;
  assign n469 = n467 | n468 ;
  assign n18698 = ~n469 ;
  assign n470 = n464 & n18698 ;
  assign n471 = n463 | n470 ;
  assign n472 = x69 & n471 ;
  assign n473 = x69 | n471 ;
  assign n474 = n18673 & n403 ;
  assign n475 = n185 & n474 ;
  assign n476 = n408 | n475 ;
  assign n477 = n408 & n475 ;
  assign n18699 = ~n477 ;
  assign n478 = n476 & n18699 ;
  assign n18700 = ~n478 ;
  assign n479 = n473 & n18700 ;
  assign n480 = n472 | n479 ;
  assign n481 = x70 & n480 ;
  assign n482 = x70 | n480 ;
  assign n483 = n411 & n18677 ;
  assign n484 = n185 & n483 ;
  assign n485 = n417 & n484 ;
  assign n486 = n417 | n484 ;
  assign n18701 = ~n485 ;
  assign n487 = n18701 & n486 ;
  assign n18702 = ~n487 ;
  assign n488 = n482 & n18702 ;
  assign n489 = n481 | n488 ;
  assign n491 = x71 | n489 ;
  assign n18703 = ~n435 ;
  assign n492 = n18703 & n491 ;
  assign n490 = x71 & n489 ;
  assign n427 = x72 & n18684 ;
  assign n493 = n18533 | n427 ;
  assign n494 = n490 | n493 ;
  assign n495 = n492 | n494 ;
  assign n496 = n322 & n428 ;
  assign n497 = n18681 & n496 ;
  assign n18704 = ~n497 ;
  assign n498 = n495 & n18704 ;
  assign n18705 = ~n490 ;
  assign n499 = n18705 & n491 ;
  assign n184 = ~n498 ;
  assign n500 = n184 & n499 ;
  assign n501 = n435 & n500 ;
  assign n502 = n435 | n500 ;
  assign n18707 = ~n501 ;
  assign n503 = n18707 & n502 ;
  assign n504 = n496 & n498 ;
  assign n18708 = ~n504 ;
  assign n508 = x73 & n18708 ;
  assign n18709 = ~x54 ;
  assign n509 = n18709 & x64 ;
  assign n510 = x65 | n509 ;
  assign n511 = x64 & n184 ;
  assign n18710 = ~n511 ;
  assign n512 = x55 & n18710 ;
  assign n513 = n436 & n184 ;
  assign n514 = n512 | n513 ;
  assign n515 = x65 & n509 ;
  assign n18711 = ~n515 ;
  assign n516 = n514 & n18711 ;
  assign n18712 = ~n516 ;
  assign n517 = n510 & n18712 ;
  assign n518 = x66 & n517 ;
  assign n519 = n18689 & n438 ;
  assign n520 = n184 & n519 ;
  assign n521 = n442 & n520 ;
  assign n522 = n442 | n520 ;
  assign n18713 = ~n521 ;
  assign n523 = n18713 & n522 ;
  assign n524 = x66 | n517 ;
  assign n18714 = ~n523 ;
  assign n525 = n18714 & n524 ;
  assign n526 = n518 | n525 ;
  assign n527 = x67 & n526 ;
  assign n528 = x67 | n526 ;
  assign n18715 = ~n445 ;
  assign n529 = n18715 & n446 ;
  assign n530 = n184 & n529 ;
  assign n531 = n451 & n530 ;
  assign n532 = n451 | n530 ;
  assign n18716 = ~n531 ;
  assign n533 = n18716 & n532 ;
  assign n18717 = ~n533 ;
  assign n534 = n528 & n18717 ;
  assign n535 = n527 | n534 ;
  assign n536 = x68 & n535 ;
  assign n537 = x68 | n535 ;
  assign n18718 = ~n454 ;
  assign n538 = n18718 & n455 ;
  assign n539 = n184 & n538 ;
  assign n540 = n460 & n539 ;
  assign n541 = n460 | n539 ;
  assign n18719 = ~n540 ;
  assign n542 = n18719 & n541 ;
  assign n18720 = ~n542 ;
  assign n543 = n537 & n18720 ;
  assign n544 = n536 | n543 ;
  assign n545 = x69 & n544 ;
  assign n546 = x69 | n544 ;
  assign n18721 = ~n463 ;
  assign n547 = n18721 & n464 ;
  assign n548 = n184 & n547 ;
  assign n549 = n18698 & n548 ;
  assign n18722 = ~n548 ;
  assign n550 = n469 & n18722 ;
  assign n551 = n549 | n550 ;
  assign n18723 = ~n551 ;
  assign n552 = n546 & n18723 ;
  assign n553 = n545 | n552 ;
  assign n554 = x70 & n553 ;
  assign n555 = x70 | n553 ;
  assign n18724 = ~n472 ;
  assign n556 = n18724 & n473 ;
  assign n557 = n184 & n556 ;
  assign n558 = n478 & n557 ;
  assign n559 = n478 | n557 ;
  assign n18725 = ~n558 ;
  assign n560 = n18725 & n559 ;
  assign n18726 = ~n560 ;
  assign n561 = n555 & n18726 ;
  assign n562 = n554 | n561 ;
  assign n563 = x71 & n562 ;
  assign n564 = x71 | n562 ;
  assign n18727 = ~n481 ;
  assign n565 = n18727 & n482 ;
  assign n566 = n184 & n565 ;
  assign n567 = n487 & n566 ;
  assign n568 = n487 | n566 ;
  assign n18728 = ~n567 ;
  assign n569 = n18728 & n568 ;
  assign n18729 = ~n569 ;
  assign n570 = n564 & n18729 ;
  assign n571 = n563 | n570 ;
  assign n574 = x72 & n571 ;
  assign n18730 = ~n574 ;
  assign n575 = n503 & n18730 ;
  assign n18731 = ~x73 ;
  assign n507 = n18731 & n504 ;
  assign n572 = x72 | n571 ;
  assign n18732 = ~n507 ;
  assign n576 = n18732 & n572 ;
  assign n18733 = ~n575 ;
  assign n577 = n18733 & n576 ;
  assign n578 = n18528 | n577 ;
  assign n579 = n508 | n578 ;
  assign n18734 = ~n571 ;
  assign n573 = x72 & n18734 ;
  assign n18735 = ~x72 ;
  assign n580 = n18735 & n571 ;
  assign n581 = n573 | n580 ;
  assign n183 = ~n579 ;
  assign n582 = n183 & n581 ;
  assign n583 = n503 & n582 ;
  assign n584 = n503 | n582 ;
  assign n18737 = ~n583 ;
  assign n585 = n18737 & n584 ;
  assign n586 = n504 & n578 ;
  assign n18738 = ~n18528 ;
  assign n587 = n18738 & n586 ;
  assign n18739 = ~x53 ;
  assign n588 = n18739 & x64 ;
  assign n590 = x65 | n588 ;
  assign n589 = x65 & n588 ;
  assign n591 = x64 & n183 ;
  assign n592 = x54 & n591 ;
  assign n593 = x54 | n591 ;
  assign n18740 = ~n592 ;
  assign n594 = n18740 & n593 ;
  assign n18741 = ~n589 ;
  assign n595 = n18741 & n594 ;
  assign n18742 = ~n595 ;
  assign n596 = n590 & n18742 ;
  assign n597 = x66 & n596 ;
  assign n598 = x66 | n596 ;
  assign n599 = n510 & n183 ;
  assign n600 = n516 & n599 ;
  assign n601 = n18711 & n599 ;
  assign n602 = n514 | n601 ;
  assign n18743 = ~n600 ;
  assign n603 = n18743 & n602 ;
  assign n18744 = ~n603 ;
  assign n604 = n598 & n18744 ;
  assign n605 = n597 | n604 ;
  assign n607 = x67 | n605 ;
  assign n606 = x67 & n605 ;
  assign n18745 = ~n518 ;
  assign n608 = n18745 & n524 ;
  assign n609 = n183 & n608 ;
  assign n610 = n523 & n609 ;
  assign n611 = n523 | n609 ;
  assign n18746 = ~n610 ;
  assign n612 = n18746 & n611 ;
  assign n18747 = ~n606 ;
  assign n613 = n18747 & n612 ;
  assign n18748 = ~n613 ;
  assign n614 = n607 & n18748 ;
  assign n615 = x68 | n614 ;
  assign n616 = x68 & n614 ;
  assign n18749 = ~n527 ;
  assign n617 = n18749 & n528 ;
  assign n618 = n183 & n617 ;
  assign n619 = n533 & n618 ;
  assign n620 = n533 | n618 ;
  assign n18750 = ~n619 ;
  assign n621 = n18750 & n620 ;
  assign n18751 = ~n616 ;
  assign n622 = n18751 & n621 ;
  assign n18752 = ~n622 ;
  assign n623 = n615 & n18752 ;
  assign n624 = x69 | n623 ;
  assign n625 = x69 & n623 ;
  assign n18753 = ~n536 ;
  assign n626 = n18753 & n537 ;
  assign n627 = n183 & n626 ;
  assign n628 = n18720 & n627 ;
  assign n18754 = ~n627 ;
  assign n629 = n542 & n18754 ;
  assign n630 = n628 | n629 ;
  assign n18755 = ~n625 ;
  assign n631 = n18755 & n630 ;
  assign n18756 = ~n631 ;
  assign n632 = n624 & n18756 ;
  assign n633 = x70 | n632 ;
  assign n634 = x70 & n632 ;
  assign n18757 = ~n545 ;
  assign n635 = n18757 & n546 ;
  assign n636 = n183 & n635 ;
  assign n637 = n18723 & n636 ;
  assign n18758 = ~n636 ;
  assign n638 = n551 & n18758 ;
  assign n639 = n637 | n638 ;
  assign n18759 = ~n634 ;
  assign n640 = n18759 & n639 ;
  assign n18760 = ~n640 ;
  assign n641 = n633 & n18760 ;
  assign n642 = x71 | n641 ;
  assign n643 = x71 & n641 ;
  assign n18761 = ~n554 ;
  assign n644 = n18761 & n555 ;
  assign n645 = n183 & n644 ;
  assign n646 = n560 & n645 ;
  assign n647 = n560 | n645 ;
  assign n18762 = ~n646 ;
  assign n648 = n18762 & n647 ;
  assign n18763 = ~n643 ;
  assign n649 = n18763 & n648 ;
  assign n18764 = ~n649 ;
  assign n650 = n642 & n18764 ;
  assign n651 = x72 | n650 ;
  assign n652 = x72 & n650 ;
  assign n18765 = ~n563 ;
  assign n653 = n18765 & n564 ;
  assign n654 = n183 & n653 ;
  assign n655 = n569 & n654 ;
  assign n656 = n569 | n654 ;
  assign n18766 = ~n655 ;
  assign n657 = n18766 & n656 ;
  assign n18767 = ~n652 ;
  assign n658 = n18767 & n657 ;
  assign n18768 = ~n658 ;
  assign n659 = n651 & n18768 ;
  assign n661 = x73 | n659 ;
  assign n18769 = ~n585 ;
  assign n662 = n18769 & n661 ;
  assign n660 = x73 & n659 ;
  assign n505 = x74 & n18708 ;
  assign n663 = n18523 | n505 ;
  assign n664 = n660 | n663 ;
  assign n665 = n662 | n664 ;
  assign n18770 = ~n587 ;
  assign n666 = n18770 & n665 ;
  assign n18771 = ~n660 ;
  assign n667 = n18771 & n661 ;
  assign n182 = ~n666 ;
  assign n668 = n182 & n667 ;
  assign n669 = n18769 & n668 ;
  assign n18773 = ~n668 ;
  assign n670 = n585 & n18773 ;
  assign n671 = n669 | n670 ;
  assign n18774 = ~x52 ;
  assign n672 = n18774 & x64 ;
  assign n673 = x65 | n672 ;
  assign n674 = x65 & n672 ;
  assign n675 = x64 & n182 ;
  assign n676 = x53 & n675 ;
  assign n677 = x53 | n675 ;
  assign n18775 = ~n676 ;
  assign n678 = n18775 & n677 ;
  assign n18776 = ~n674 ;
  assign n679 = n18776 & n678 ;
  assign n18777 = ~n679 ;
  assign n680 = n673 & n18777 ;
  assign n682 = x66 | n680 ;
  assign n681 = x66 & n680 ;
  assign n683 = n18741 & n590 ;
  assign n684 = n182 & n683 ;
  assign n685 = n594 & n684 ;
  assign n686 = n594 | n684 ;
  assign n18778 = ~n685 ;
  assign n687 = n18778 & n686 ;
  assign n18779 = ~n681 ;
  assign n688 = n18779 & n687 ;
  assign n18780 = ~n688 ;
  assign n689 = n682 & n18780 ;
  assign n690 = x67 | n689 ;
  assign n691 = x67 & n689 ;
  assign n18781 = ~n597 ;
  assign n692 = n18781 & n598 ;
  assign n693 = n182 & n692 ;
  assign n18782 = ~n693 ;
  assign n694 = n603 & n18782 ;
  assign n695 = n18744 & n693 ;
  assign n696 = n694 | n695 ;
  assign n18783 = ~n691 ;
  assign n697 = n18783 & n696 ;
  assign n18784 = ~n697 ;
  assign n698 = n690 & n18784 ;
  assign n699 = x68 | n698 ;
  assign n700 = x68 & n698 ;
  assign n701 = n18747 & n607 ;
  assign n702 = n182 & n701 ;
  assign n18785 = ~n612 ;
  assign n703 = n18785 & n702 ;
  assign n18786 = ~n702 ;
  assign n704 = n612 & n18786 ;
  assign n705 = n703 | n704 ;
  assign n18787 = ~n700 ;
  assign n706 = n18787 & n705 ;
  assign n18788 = ~n706 ;
  assign n707 = n699 & n18788 ;
  assign n708 = x69 | n707 ;
  assign n709 = x69 & n707 ;
  assign n710 = n615 & n18751 ;
  assign n711 = n182 & n710 ;
  assign n18789 = ~n621 ;
  assign n712 = n18789 & n711 ;
  assign n18790 = ~n711 ;
  assign n713 = n621 & n18790 ;
  assign n714 = n712 | n713 ;
  assign n18791 = ~n709 ;
  assign n715 = n18791 & n714 ;
  assign n18792 = ~n715 ;
  assign n716 = n708 & n18792 ;
  assign n717 = x70 | n716 ;
  assign n718 = x70 & n716 ;
  assign n719 = n624 & n18755 ;
  assign n720 = n182 & n719 ;
  assign n18793 = ~n630 ;
  assign n721 = n18793 & n720 ;
  assign n18794 = ~n720 ;
  assign n722 = n630 & n18794 ;
  assign n723 = n721 | n722 ;
  assign n18795 = ~n718 ;
  assign n724 = n18795 & n723 ;
  assign n18796 = ~n724 ;
  assign n725 = n717 & n18796 ;
  assign n726 = x71 | n725 ;
  assign n727 = x71 & n725 ;
  assign n728 = n633 & n18759 ;
  assign n729 = n182 & n728 ;
  assign n18797 = ~n639 ;
  assign n730 = n18797 & n729 ;
  assign n18798 = ~n729 ;
  assign n731 = n639 & n18798 ;
  assign n732 = n730 | n731 ;
  assign n18799 = ~n727 ;
  assign n733 = n18799 & n732 ;
  assign n18800 = ~n733 ;
  assign n734 = n726 & n18800 ;
  assign n735 = x72 | n734 ;
  assign n736 = x72 & n734 ;
  assign n737 = n642 & n18763 ;
  assign n738 = n182 & n737 ;
  assign n739 = n648 & n738 ;
  assign n740 = n648 | n738 ;
  assign n18801 = ~n739 ;
  assign n741 = n18801 & n740 ;
  assign n18802 = ~n736 ;
  assign n742 = n18802 & n741 ;
  assign n18803 = ~n742 ;
  assign n743 = n735 & n18803 ;
  assign n744 = x73 | n743 ;
  assign n745 = x73 & n743 ;
  assign n746 = n651 & n18767 ;
  assign n747 = n182 & n746 ;
  assign n748 = n657 & n747 ;
  assign n749 = n657 | n747 ;
  assign n18804 = ~n748 ;
  assign n750 = n18804 & n749 ;
  assign n18805 = ~n745 ;
  assign n751 = n18805 & n750 ;
  assign n18806 = ~n751 ;
  assign n752 = n744 & n18806 ;
  assign n755 = x74 & n752 ;
  assign n18807 = ~n755 ;
  assign n756 = n671 & n18807 ;
  assign n753 = x74 | n752 ;
  assign n506 = n18528 & n504 ;
  assign n757 = n506 & n665 ;
  assign n18808 = ~x75 ;
  assign n758 = n18808 & n757 ;
  assign n18809 = ~n758 ;
  assign n759 = n753 & n18809 ;
  assign n18810 = ~n756 ;
  assign n760 = n18810 & n759 ;
  assign n761 = n18518 | n760 ;
  assign n18811 = ~n586 ;
  assign n762 = x75 & n18811 ;
  assign n763 = n761 | n762 ;
  assign n18812 = ~n752 ;
  assign n754 = x74 & n18812 ;
  assign n18813 = ~x74 ;
  assign n764 = n18813 & n752 ;
  assign n765 = n754 | n764 ;
  assign n181 = ~n763 ;
  assign n766 = n181 & n765 ;
  assign n18815 = ~n671 ;
  assign n767 = n18815 & n766 ;
  assign n18816 = ~n766 ;
  assign n768 = n671 & n18816 ;
  assign n769 = n767 | n768 ;
  assign n18817 = ~x51 ;
  assign n773 = n18817 & x64 ;
  assign n774 = x65 | n773 ;
  assign n775 = x65 & n773 ;
  assign n776 = x64 & n181 ;
  assign n777 = x52 & n776 ;
  assign n778 = x52 | n776 ;
  assign n18818 = ~n777 ;
  assign n779 = n18818 & n778 ;
  assign n18819 = ~n775 ;
  assign n780 = n18819 & n779 ;
  assign n18820 = ~n780 ;
  assign n781 = n774 & n18820 ;
  assign n783 = x66 | n781 ;
  assign n782 = x66 & n781 ;
  assign n784 = n673 & n18776 ;
  assign n785 = n181 & n784 ;
  assign n786 = n678 & n785 ;
  assign n787 = n678 | n785 ;
  assign n18821 = ~n786 ;
  assign n788 = n18821 & n787 ;
  assign n18822 = ~n782 ;
  assign n789 = n18822 & n788 ;
  assign n18823 = ~n789 ;
  assign n790 = n783 & n18823 ;
  assign n791 = x67 & n790 ;
  assign n792 = x67 | n790 ;
  assign n793 = n682 & n181 ;
  assign n794 = n688 & n793 ;
  assign n795 = n18779 & n793 ;
  assign n796 = n687 | n795 ;
  assign n18824 = ~n794 ;
  assign n797 = n18824 & n796 ;
  assign n18825 = ~n797 ;
  assign n798 = n792 & n18825 ;
  assign n799 = n791 | n798 ;
  assign n800 = x68 & n799 ;
  assign n801 = x68 | n799 ;
  assign n802 = n690 & n181 ;
  assign n803 = n697 & n802 ;
  assign n804 = n18783 & n802 ;
  assign n805 = n696 | n804 ;
  assign n18826 = ~n803 ;
  assign n806 = n18826 & n805 ;
  assign n18827 = ~n806 ;
  assign n807 = n801 & n18827 ;
  assign n808 = n800 | n807 ;
  assign n810 = x69 | n808 ;
  assign n809 = x69 & n808 ;
  assign n811 = n699 & n18787 ;
  assign n812 = n181 & n811 ;
  assign n18828 = ~n705 ;
  assign n813 = n18828 & n812 ;
  assign n18829 = ~n812 ;
  assign n814 = n705 & n18829 ;
  assign n815 = n813 | n814 ;
  assign n18830 = ~n809 ;
  assign n816 = n18830 & n815 ;
  assign n18831 = ~n816 ;
  assign n817 = n810 & n18831 ;
  assign n818 = x70 | n817 ;
  assign n819 = x70 & n817 ;
  assign n820 = n708 & n18791 ;
  assign n821 = n181 & n820 ;
  assign n822 = n714 & n821 ;
  assign n823 = n714 | n821 ;
  assign n18832 = ~n822 ;
  assign n824 = n18832 & n823 ;
  assign n18833 = ~n819 ;
  assign n825 = n18833 & n824 ;
  assign n18834 = ~n825 ;
  assign n826 = n818 & n18834 ;
  assign n827 = x71 | n826 ;
  assign n828 = x71 & n826 ;
  assign n829 = n717 & n18795 ;
  assign n830 = n181 & n829 ;
  assign n831 = n723 & n830 ;
  assign n832 = n723 | n830 ;
  assign n18835 = ~n831 ;
  assign n833 = n18835 & n832 ;
  assign n18836 = ~n828 ;
  assign n834 = n18836 & n833 ;
  assign n18837 = ~n834 ;
  assign n835 = n827 & n18837 ;
  assign n836 = x72 | n835 ;
  assign n837 = x72 & n835 ;
  assign n838 = n726 & n18799 ;
  assign n839 = n181 & n838 ;
  assign n840 = n732 & n839 ;
  assign n841 = n732 | n839 ;
  assign n18838 = ~n840 ;
  assign n842 = n18838 & n841 ;
  assign n18839 = ~n837 ;
  assign n843 = n18839 & n842 ;
  assign n18840 = ~n843 ;
  assign n844 = n836 & n18840 ;
  assign n845 = x73 | n844 ;
  assign n846 = x73 & n844 ;
  assign n847 = n735 & n18802 ;
  assign n848 = n181 & n847 ;
  assign n849 = n741 & n848 ;
  assign n850 = n741 | n848 ;
  assign n18841 = ~n849 ;
  assign n851 = n18841 & n850 ;
  assign n18842 = ~n846 ;
  assign n852 = n18842 & n851 ;
  assign n18843 = ~n852 ;
  assign n853 = n845 & n18843 ;
  assign n854 = x74 | n853 ;
  assign n855 = x74 & n853 ;
  assign n856 = n744 & n18805 ;
  assign n857 = n181 & n856 ;
  assign n858 = n750 & n857 ;
  assign n859 = n750 | n857 ;
  assign n18844 = ~n858 ;
  assign n860 = n18844 & n859 ;
  assign n18845 = ~n855 ;
  assign n861 = n18845 & n860 ;
  assign n18846 = ~n861 ;
  assign n862 = n854 & n18846 ;
  assign n864 = x75 & n862 ;
  assign n18847 = ~n864 ;
  assign n865 = n769 & n18847 ;
  assign n770 = n757 & n761 ;
  assign n771 = n21884 | n770 ;
  assign n18848 = ~x76 ;
  assign n772 = n18848 & n771 ;
  assign n863 = x75 | n862 ;
  assign n18849 = ~n772 ;
  assign n866 = n18849 & n863 ;
  assign n18850 = ~n865 ;
  assign n867 = n18850 & n866 ;
  assign n868 = n18513 | n867 ;
  assign n18851 = ~n771 ;
  assign n870 = x76 & n18851 ;
  assign n871 = n868 | n870 ;
  assign n872 = n863 & n18847 ;
  assign n180 = ~n871 ;
  assign n873 = n180 & n872 ;
  assign n18853 = ~n769 ;
  assign n874 = n18853 & n873 ;
  assign n18854 = ~n873 ;
  assign n875 = n769 & n18854 ;
  assign n876 = n874 | n875 ;
  assign n869 = n21884 | n868 ;
  assign n877 = n771 & n869 ;
  assign n18855 = ~n877 ;
  assign n878 = x77 & n18855 ;
  assign n879 = n18508 | n878 ;
  assign n18856 = ~x50 ;
  assign n880 = n18856 & x64 ;
  assign n882 = x65 | n880 ;
  assign n881 = x65 & n880 ;
  assign n883 = x64 & n180 ;
  assign n884 = x51 & n883 ;
  assign n885 = x51 | n883 ;
  assign n18857 = ~n884 ;
  assign n886 = n18857 & n885 ;
  assign n18858 = ~n881 ;
  assign n887 = n18858 & n886 ;
  assign n18859 = ~n887 ;
  assign n888 = n882 & n18859 ;
  assign n889 = x66 & n888 ;
  assign n890 = x66 | n888 ;
  assign n891 = n774 & n18819 ;
  assign n892 = n180 & n891 ;
  assign n893 = n779 & n892 ;
  assign n894 = n779 | n892 ;
  assign n18860 = ~n893 ;
  assign n895 = n18860 & n894 ;
  assign n18861 = ~n895 ;
  assign n896 = n890 & n18861 ;
  assign n897 = n889 | n896 ;
  assign n898 = x67 & n897 ;
  assign n899 = x67 | n897 ;
  assign n900 = n783 & n180 ;
  assign n901 = n789 & n900 ;
  assign n902 = n18822 & n900 ;
  assign n903 = n788 | n902 ;
  assign n18862 = ~n901 ;
  assign n904 = n18862 & n903 ;
  assign n18863 = ~n904 ;
  assign n905 = n899 & n18863 ;
  assign n906 = n898 | n905 ;
  assign n907 = x68 & n906 ;
  assign n908 = x68 | n906 ;
  assign n18864 = ~n791 ;
  assign n909 = n18864 & n792 ;
  assign n910 = n180 & n909 ;
  assign n911 = n797 & n910 ;
  assign n912 = n797 | n910 ;
  assign n18865 = ~n911 ;
  assign n913 = n18865 & n912 ;
  assign n18866 = ~n913 ;
  assign n914 = n908 & n18866 ;
  assign n915 = n907 | n914 ;
  assign n916 = x69 & n915 ;
  assign n917 = x69 | n915 ;
  assign n18867 = ~n800 ;
  assign n918 = n18867 & n801 ;
  assign n919 = n180 & n918 ;
  assign n920 = n806 & n919 ;
  assign n921 = n806 | n919 ;
  assign n18868 = ~n920 ;
  assign n922 = n18868 & n921 ;
  assign n18869 = ~n922 ;
  assign n923 = n917 & n18869 ;
  assign n924 = n916 | n923 ;
  assign n925 = x70 & n924 ;
  assign n926 = x70 | n924 ;
  assign n927 = n18830 & n810 ;
  assign n928 = n180 & n927 ;
  assign n18870 = ~n815 ;
  assign n929 = n18870 & n928 ;
  assign n18871 = ~n928 ;
  assign n930 = n815 & n18871 ;
  assign n931 = n929 | n930 ;
  assign n18872 = ~n931 ;
  assign n932 = n926 & n18872 ;
  assign n933 = n925 | n932 ;
  assign n934 = x71 & n933 ;
  assign n935 = x71 | n933 ;
  assign n936 = n818 & n18833 ;
  assign n937 = n180 & n936 ;
  assign n938 = n824 & n937 ;
  assign n939 = n824 | n937 ;
  assign n18873 = ~n938 ;
  assign n940 = n18873 & n939 ;
  assign n18874 = ~n940 ;
  assign n941 = n935 & n18874 ;
  assign n942 = n934 | n941 ;
  assign n943 = x72 & n942 ;
  assign n944 = x72 | n942 ;
  assign n945 = n827 & n18836 ;
  assign n946 = n180 & n945 ;
  assign n947 = n833 & n946 ;
  assign n948 = n833 | n946 ;
  assign n18875 = ~n947 ;
  assign n949 = n18875 & n948 ;
  assign n18876 = ~n949 ;
  assign n950 = n944 & n18876 ;
  assign n951 = n943 | n950 ;
  assign n952 = x73 & n951 ;
  assign n953 = x73 | n951 ;
  assign n954 = n836 & n18839 ;
  assign n955 = n180 & n954 ;
  assign n956 = n842 & n955 ;
  assign n957 = n842 | n955 ;
  assign n18877 = ~n956 ;
  assign n958 = n18877 & n957 ;
  assign n18878 = ~n958 ;
  assign n959 = n953 & n18878 ;
  assign n960 = n952 | n959 ;
  assign n961 = x74 & n960 ;
  assign n962 = x74 | n960 ;
  assign n963 = n845 & n18842 ;
  assign n964 = n180 & n963 ;
  assign n965 = n851 & n964 ;
  assign n966 = n851 | n964 ;
  assign n18879 = ~n965 ;
  assign n967 = n18879 & n966 ;
  assign n18880 = ~n967 ;
  assign n968 = n962 & n18880 ;
  assign n969 = n961 | n968 ;
  assign n970 = x75 & n969 ;
  assign n971 = x75 | n969 ;
  assign n972 = n854 & n18845 ;
  assign n973 = n180 & n972 ;
  assign n974 = n860 & n973 ;
  assign n975 = n860 | n973 ;
  assign n18881 = ~n974 ;
  assign n976 = n18881 & n975 ;
  assign n18882 = ~n976 ;
  assign n977 = n971 & n18882 ;
  assign n978 = n970 | n977 ;
  assign n979 = x76 & n978 ;
  assign n18883 = ~n979 ;
  assign n980 = n876 & n18883 ;
  assign n18884 = ~x77 ;
  assign n981 = n18884 & n877 ;
  assign n982 = x76 | n978 ;
  assign n18885 = ~n981 ;
  assign n983 = n18885 & n982 ;
  assign n18886 = ~n980 ;
  assign n984 = n18886 & n983 ;
  assign n985 = n879 | n984 ;
  assign n987 = n18883 & n982 ;
  assign n179 = ~n985 ;
  assign n988 = n179 & n987 ;
  assign n18888 = ~n876 ;
  assign n989 = n18888 & n988 ;
  assign n18889 = ~n988 ;
  assign n990 = n876 & n18889 ;
  assign n991 = n989 | n990 ;
  assign n986 = n21884 | n985 ;
  assign n992 = n877 & n986 ;
  assign n18890 = ~n18508 ;
  assign n994 = n18890 & n992 ;
  assign n18891 = ~x49 ;
  assign n995 = n18891 & x64 ;
  assign n996 = x65 | n995 ;
  assign n997 = x65 & n995 ;
  assign n998 = x64 & n179 ;
  assign n999 = x50 & n998 ;
  assign n1000 = x50 | n998 ;
  assign n18892 = ~n999 ;
  assign n1001 = n18892 & n1000 ;
  assign n18893 = ~n997 ;
  assign n1002 = n18893 & n1001 ;
  assign n18894 = ~n1002 ;
  assign n1003 = n996 & n18894 ;
  assign n1005 = x66 | n1003 ;
  assign n1004 = x66 & n1003 ;
  assign n1006 = n18858 & n882 ;
  assign n1007 = n179 & n1006 ;
  assign n1008 = n886 & n1007 ;
  assign n1009 = n886 | n1007 ;
  assign n18895 = ~n1008 ;
  assign n1010 = n18895 & n1009 ;
  assign n18896 = ~n1004 ;
  assign n1011 = n18896 & n1010 ;
  assign n18897 = ~n1011 ;
  assign n1012 = n1005 & n18897 ;
  assign n1013 = x67 | n1012 ;
  assign n1014 = x67 & n1012 ;
  assign n18898 = ~n889 ;
  assign n1015 = n18898 & n890 ;
  assign n1016 = n179 & n1015 ;
  assign n1017 = n895 & n1016 ;
  assign n1018 = n895 | n1016 ;
  assign n18899 = ~n1017 ;
  assign n1019 = n18899 & n1018 ;
  assign n18900 = ~n1014 ;
  assign n1020 = n18900 & n1019 ;
  assign n18901 = ~n1020 ;
  assign n1021 = n1013 & n18901 ;
  assign n1022 = x68 | n1021 ;
  assign n1023 = x68 & n1021 ;
  assign n18902 = ~n898 ;
  assign n1024 = n18902 & n899 ;
  assign n1025 = n179 & n1024 ;
  assign n1026 = n904 & n1025 ;
  assign n1027 = n904 | n1025 ;
  assign n18903 = ~n1026 ;
  assign n1028 = n18903 & n1027 ;
  assign n18904 = ~n1023 ;
  assign n1029 = n18904 & n1028 ;
  assign n18905 = ~n1029 ;
  assign n1030 = n1022 & n18905 ;
  assign n1031 = x69 | n1030 ;
  assign n1032 = x69 & n1030 ;
  assign n18906 = ~n907 ;
  assign n1033 = n18906 & n908 ;
  assign n1034 = n179 & n1033 ;
  assign n1035 = n18866 & n1034 ;
  assign n18907 = ~n1034 ;
  assign n1036 = n913 & n18907 ;
  assign n1037 = n1035 | n1036 ;
  assign n18908 = ~n1032 ;
  assign n1038 = n18908 & n1037 ;
  assign n18909 = ~n1038 ;
  assign n1039 = n1031 & n18909 ;
  assign n1040 = x70 | n1039 ;
  assign n1041 = x70 & n1039 ;
  assign n18910 = ~n916 ;
  assign n1042 = n18910 & n917 ;
  assign n1043 = n179 & n1042 ;
  assign n1044 = n18869 & n1043 ;
  assign n18911 = ~n1043 ;
  assign n1045 = n922 & n18911 ;
  assign n1046 = n1044 | n1045 ;
  assign n18912 = ~n1041 ;
  assign n1047 = n18912 & n1046 ;
  assign n18913 = ~n1047 ;
  assign n1048 = n1040 & n18913 ;
  assign n1049 = x71 | n1048 ;
  assign n1050 = x71 & n1048 ;
  assign n18914 = ~n925 ;
  assign n1051 = n18914 & n926 ;
  assign n1052 = n179 & n1051 ;
  assign n1053 = n931 & n1052 ;
  assign n1054 = n931 | n1052 ;
  assign n18915 = ~n1053 ;
  assign n1055 = n18915 & n1054 ;
  assign n18916 = ~n1050 ;
  assign n1056 = n18916 & n1055 ;
  assign n18917 = ~n1056 ;
  assign n1057 = n1049 & n18917 ;
  assign n1058 = x72 | n1057 ;
  assign n1059 = x72 & n1057 ;
  assign n18918 = ~n934 ;
  assign n1060 = n18918 & n935 ;
  assign n1061 = n179 & n1060 ;
  assign n1062 = n940 & n1061 ;
  assign n1063 = n940 | n1061 ;
  assign n18919 = ~n1062 ;
  assign n1064 = n18919 & n1063 ;
  assign n18920 = ~n1059 ;
  assign n1065 = n18920 & n1064 ;
  assign n18921 = ~n1065 ;
  assign n1066 = n1058 & n18921 ;
  assign n1067 = x73 | n1066 ;
  assign n1068 = x73 & n1066 ;
  assign n18922 = ~n943 ;
  assign n1069 = n18922 & n944 ;
  assign n1070 = n179 & n1069 ;
  assign n1071 = n949 & n1070 ;
  assign n1072 = n949 | n1070 ;
  assign n18923 = ~n1071 ;
  assign n1073 = n18923 & n1072 ;
  assign n18924 = ~n1068 ;
  assign n1074 = n18924 & n1073 ;
  assign n18925 = ~n1074 ;
  assign n1075 = n1067 & n18925 ;
  assign n1076 = x74 | n1075 ;
  assign n1077 = x74 & n1075 ;
  assign n18926 = ~n952 ;
  assign n1078 = n18926 & n953 ;
  assign n1079 = n179 & n1078 ;
  assign n1080 = n958 & n1079 ;
  assign n1081 = n958 | n1079 ;
  assign n18927 = ~n1080 ;
  assign n1082 = n18927 & n1081 ;
  assign n18928 = ~n1077 ;
  assign n1083 = n18928 & n1082 ;
  assign n18929 = ~n1083 ;
  assign n1084 = n1076 & n18929 ;
  assign n1085 = x75 | n1084 ;
  assign n1086 = x75 & n1084 ;
  assign n18930 = ~n961 ;
  assign n1087 = n18930 & n962 ;
  assign n1088 = n179 & n1087 ;
  assign n1089 = n967 & n1088 ;
  assign n1090 = n967 | n1088 ;
  assign n18931 = ~n1089 ;
  assign n1091 = n18931 & n1090 ;
  assign n18932 = ~n1086 ;
  assign n1092 = n18932 & n1091 ;
  assign n18933 = ~n1092 ;
  assign n1093 = n1085 & n18933 ;
  assign n1094 = x76 | n1093 ;
  assign n1095 = x76 & n1093 ;
  assign n18934 = ~n970 ;
  assign n1096 = n18934 & n971 ;
  assign n1097 = n179 & n1096 ;
  assign n1098 = n976 & n1097 ;
  assign n1099 = n976 | n1097 ;
  assign n18935 = ~n1098 ;
  assign n1100 = n18935 & n1099 ;
  assign n18936 = ~n1095 ;
  assign n1101 = n18936 & n1100 ;
  assign n18937 = ~n1101 ;
  assign n1102 = n1094 & n18937 ;
  assign n1104 = x77 | n1102 ;
  assign n18938 = ~n991 ;
  assign n1105 = n18938 & n1104 ;
  assign n1103 = x77 & n1102 ;
  assign n1106 = n18503 | n994 ;
  assign n18939 = ~n992 ;
  assign n1107 = x78 & n18939 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = n1103 | n1108 ;
  assign n1110 = n1105 | n1109 ;
  assign n18940 = ~n994 ;
  assign n1111 = n18940 & n1110 ;
  assign n18941 = ~n1103 ;
  assign n1112 = n18941 & n1104 ;
  assign n178 = ~n1111 ;
  assign n1113 = n178 & n1112 ;
  assign n1114 = n18938 & n1113 ;
  assign n18943 = ~n1113 ;
  assign n1115 = n991 & n18943 ;
  assign n1116 = n1114 | n1115 ;
  assign n18944 = ~x48 ;
  assign n1117 = n18944 & x64 ;
  assign n1119 = x65 | n1117 ;
  assign n1118 = x65 & n1117 ;
  assign n1120 = x64 & n178 ;
  assign n1121 = x49 & n1120 ;
  assign n1122 = x49 | n1120 ;
  assign n18945 = ~n1121 ;
  assign n1123 = n18945 & n1122 ;
  assign n18946 = ~n1118 ;
  assign n1124 = n18946 & n1123 ;
  assign n18947 = ~n1124 ;
  assign n1125 = n1119 & n18947 ;
  assign n1126 = x66 & n1125 ;
  assign n1127 = x66 | n1125 ;
  assign n1128 = n996 & n18893 ;
  assign n1129 = n178 & n1128 ;
  assign n1130 = n1001 & n1129 ;
  assign n1131 = n1001 | n1129 ;
  assign n18948 = ~n1130 ;
  assign n1132 = n18948 & n1131 ;
  assign n18949 = ~n1132 ;
  assign n1133 = n1127 & n18949 ;
  assign n1134 = n1126 | n1133 ;
  assign n1135 = x67 & n1134 ;
  assign n1136 = x67 | n1134 ;
  assign n1137 = n1005 & n178 ;
  assign n1138 = n1011 & n1137 ;
  assign n1139 = n18896 & n1137 ;
  assign n1140 = n1010 | n1139 ;
  assign n18950 = ~n1138 ;
  assign n1141 = n18950 & n1140 ;
  assign n18951 = ~n1141 ;
  assign n1142 = n1136 & n18951 ;
  assign n1143 = n1135 | n1142 ;
  assign n1144 = x68 & n1143 ;
  assign n1145 = x68 | n1143 ;
  assign n1146 = n1013 & n18900 ;
  assign n1147 = n178 & n1146 ;
  assign n18952 = ~n1019 ;
  assign n1148 = n18952 & n1147 ;
  assign n18953 = ~n1147 ;
  assign n1149 = n1019 & n18953 ;
  assign n1150 = n1148 | n1149 ;
  assign n18954 = ~n1150 ;
  assign n1151 = n1145 & n18954 ;
  assign n1152 = n1144 | n1151 ;
  assign n1153 = x69 & n1152 ;
  assign n1154 = x69 | n1152 ;
  assign n1155 = n1022 & n18904 ;
  assign n1156 = n178 & n1155 ;
  assign n18955 = ~n1028 ;
  assign n1157 = n18955 & n1156 ;
  assign n18956 = ~n1156 ;
  assign n1158 = n1028 & n18956 ;
  assign n1159 = n1157 | n1158 ;
  assign n18957 = ~n1159 ;
  assign n1160 = n1154 & n18957 ;
  assign n1161 = n1153 | n1160 ;
  assign n1162 = x70 & n1161 ;
  assign n1163 = x70 | n1161 ;
  assign n1164 = n1031 & n18908 ;
  assign n1165 = n178 & n1164 ;
  assign n18958 = ~n1037 ;
  assign n1166 = n18958 & n1165 ;
  assign n18959 = ~n1165 ;
  assign n1167 = n1037 & n18959 ;
  assign n1168 = n1166 | n1167 ;
  assign n18960 = ~n1168 ;
  assign n1169 = n1163 & n18960 ;
  assign n1170 = n1162 | n1169 ;
  assign n1171 = x71 & n1170 ;
  assign n1172 = x71 | n1170 ;
  assign n1173 = n1040 & n18912 ;
  assign n1174 = n178 & n1173 ;
  assign n18961 = ~n1046 ;
  assign n1175 = n18961 & n1174 ;
  assign n18962 = ~n1174 ;
  assign n1176 = n1046 & n18962 ;
  assign n1177 = n1175 | n1176 ;
  assign n18963 = ~n1177 ;
  assign n1178 = n1172 & n18963 ;
  assign n1179 = n1171 | n1178 ;
  assign n1180 = x72 & n1179 ;
  assign n1181 = x72 | n1179 ;
  assign n1182 = n1049 & n18916 ;
  assign n1183 = n178 & n1182 ;
  assign n1184 = n1055 & n1183 ;
  assign n1185 = n1055 | n1183 ;
  assign n18964 = ~n1184 ;
  assign n1186 = n18964 & n1185 ;
  assign n18965 = ~n1186 ;
  assign n1187 = n1181 & n18965 ;
  assign n1188 = n1180 | n1187 ;
  assign n1189 = x73 & n1188 ;
  assign n1190 = x73 | n1188 ;
  assign n1191 = n1058 & n18920 ;
  assign n1192 = n178 & n1191 ;
  assign n1193 = n1064 & n1192 ;
  assign n1194 = n1064 | n1192 ;
  assign n18966 = ~n1193 ;
  assign n1195 = n18966 & n1194 ;
  assign n18967 = ~n1195 ;
  assign n1196 = n1190 & n18967 ;
  assign n1197 = n1189 | n1196 ;
  assign n1198 = x74 & n1197 ;
  assign n1199 = x74 | n1197 ;
  assign n1200 = n1067 & n18924 ;
  assign n1201 = n178 & n1200 ;
  assign n1202 = n1073 & n1201 ;
  assign n1203 = n1073 | n1201 ;
  assign n18968 = ~n1202 ;
  assign n1204 = n18968 & n1203 ;
  assign n18969 = ~n1204 ;
  assign n1205 = n1199 & n18969 ;
  assign n1206 = n1198 | n1205 ;
  assign n1207 = x75 & n1206 ;
  assign n1208 = x75 | n1206 ;
  assign n1209 = n1076 & n18928 ;
  assign n1210 = n178 & n1209 ;
  assign n1211 = n1082 & n1210 ;
  assign n1212 = n1082 | n1210 ;
  assign n18970 = ~n1211 ;
  assign n1213 = n18970 & n1212 ;
  assign n18971 = ~n1213 ;
  assign n1214 = n1208 & n18971 ;
  assign n1215 = n1207 | n1214 ;
  assign n1216 = x76 & n1215 ;
  assign n1217 = x76 | n1215 ;
  assign n1218 = n1085 & n18932 ;
  assign n1219 = n178 & n1218 ;
  assign n1220 = n1091 & n1219 ;
  assign n1221 = n1091 | n1219 ;
  assign n18972 = ~n1220 ;
  assign n1222 = n18972 & n1221 ;
  assign n18973 = ~n1222 ;
  assign n1223 = n1217 & n18973 ;
  assign n1224 = n1216 | n1223 ;
  assign n1225 = x77 & n1224 ;
  assign n1226 = x77 | n1224 ;
  assign n1227 = n1094 & n18936 ;
  assign n1228 = n178 & n1227 ;
  assign n1229 = n1100 & n1228 ;
  assign n1230 = n1100 | n1228 ;
  assign n18974 = ~n1229 ;
  assign n1231 = n18974 & n1230 ;
  assign n18975 = ~n1231 ;
  assign n1232 = n1226 & n18975 ;
  assign n1233 = n1225 | n1232 ;
  assign n1236 = x78 & n1233 ;
  assign n18976 = ~n1236 ;
  assign n1237 = n1116 & n18976 ;
  assign n1234 = x78 | n1233 ;
  assign n993 = n18508 & n992 ;
  assign n1238 = n993 & n1110 ;
  assign n1239 = n21884 | n1238 ;
  assign n18977 = ~x79 ;
  assign n1240 = n18977 & n1239 ;
  assign n18978 = ~n1240 ;
  assign n1241 = n1234 & n18978 ;
  assign n18979 = ~n1237 ;
  assign n1242 = n18979 & n1241 ;
  assign n1243 = n18498 | n1242 ;
  assign n18980 = ~n1239 ;
  assign n1244 = x79 & n18980 ;
  assign n1245 = n1243 | n1244 ;
  assign n18981 = ~n1233 ;
  assign n1235 = x78 & n18981 ;
  assign n18982 = ~x78 ;
  assign n1246 = n18982 & n1233 ;
  assign n1247 = n1235 | n1246 ;
  assign n177 = ~n1245 ;
  assign n1248 = n177 & n1247 ;
  assign n1249 = n1116 & n1248 ;
  assign n1250 = n1116 | n1248 ;
  assign n18984 = ~n1249 ;
  assign n1251 = n18984 & n1250 ;
  assign n18985 = ~x47 ;
  assign n1255 = n18985 & x64 ;
  assign n1257 = x65 | n1255 ;
  assign n1256 = x65 & n1255 ;
  assign n1258 = x64 & n177 ;
  assign n1259 = x48 & n1258 ;
  assign n1260 = x48 | n1258 ;
  assign n18986 = ~n1259 ;
  assign n1261 = n18986 & n1260 ;
  assign n18987 = ~n1256 ;
  assign n1262 = n18987 & n1261 ;
  assign n18988 = ~n1262 ;
  assign n1263 = n1257 & n18988 ;
  assign n1264 = x66 & n1263 ;
  assign n1265 = x66 | n1263 ;
  assign n1266 = n18946 & n1119 ;
  assign n1267 = n177 & n1266 ;
  assign n1268 = n1123 & n1267 ;
  assign n1269 = n1123 | n1267 ;
  assign n18989 = ~n1268 ;
  assign n1270 = n18989 & n1269 ;
  assign n18990 = ~n1270 ;
  assign n1271 = n1265 & n18990 ;
  assign n1272 = n1264 | n1271 ;
  assign n1273 = x67 & n1272 ;
  assign n1274 = x67 | n1272 ;
  assign n18991 = ~n1126 ;
  assign n1275 = n18991 & n1127 ;
  assign n1276 = n177 & n1275 ;
  assign n1277 = n1132 & n1276 ;
  assign n1278 = n1132 | n1276 ;
  assign n18992 = ~n1277 ;
  assign n1279 = n18992 & n1278 ;
  assign n18993 = ~n1279 ;
  assign n1280 = n1274 & n18993 ;
  assign n1281 = n1273 | n1280 ;
  assign n1282 = x68 & n1281 ;
  assign n1283 = x68 | n1281 ;
  assign n18994 = ~n1135 ;
  assign n1284 = n18994 & n1136 ;
  assign n1285 = n177 & n1284 ;
  assign n1286 = n1141 & n1285 ;
  assign n1287 = n1141 | n1285 ;
  assign n18995 = ~n1286 ;
  assign n1288 = n18995 & n1287 ;
  assign n18996 = ~n1288 ;
  assign n1289 = n1283 & n18996 ;
  assign n1290 = n1282 | n1289 ;
  assign n1291 = x69 & n1290 ;
  assign n1292 = x69 | n1290 ;
  assign n18997 = ~n1144 ;
  assign n1293 = n18997 & n1145 ;
  assign n1294 = n177 & n1293 ;
  assign n1295 = n1150 & n1294 ;
  assign n1296 = n1150 | n1294 ;
  assign n18998 = ~n1295 ;
  assign n1297 = n18998 & n1296 ;
  assign n18999 = ~n1297 ;
  assign n1298 = n1292 & n18999 ;
  assign n1299 = n1291 | n1298 ;
  assign n1300 = x70 & n1299 ;
  assign n1301 = x70 | n1299 ;
  assign n19000 = ~n1153 ;
  assign n1302 = n19000 & n1154 ;
  assign n1303 = n177 & n1302 ;
  assign n1304 = n18957 & n1303 ;
  assign n19001 = ~n1303 ;
  assign n1305 = n1159 & n19001 ;
  assign n1306 = n1304 | n1305 ;
  assign n19002 = ~n1306 ;
  assign n1307 = n1301 & n19002 ;
  assign n1308 = n1300 | n1307 ;
  assign n1309 = x71 & n1308 ;
  assign n1310 = x71 | n1308 ;
  assign n19003 = ~n1162 ;
  assign n1311 = n19003 & n1163 ;
  assign n1312 = n177 & n1311 ;
  assign n1313 = n1168 & n1312 ;
  assign n1314 = n1168 | n1312 ;
  assign n19004 = ~n1313 ;
  assign n1315 = n19004 & n1314 ;
  assign n19005 = ~n1315 ;
  assign n1316 = n1310 & n19005 ;
  assign n1317 = n1309 | n1316 ;
  assign n1318 = x72 & n1317 ;
  assign n1319 = x72 | n1317 ;
  assign n19006 = ~n1171 ;
  assign n1320 = n19006 & n1172 ;
  assign n1321 = n177 & n1320 ;
  assign n1322 = n1177 & n1321 ;
  assign n1323 = n1177 | n1321 ;
  assign n19007 = ~n1322 ;
  assign n1324 = n19007 & n1323 ;
  assign n19008 = ~n1324 ;
  assign n1325 = n1319 & n19008 ;
  assign n1326 = n1318 | n1325 ;
  assign n1327 = x73 & n1326 ;
  assign n1328 = x73 | n1326 ;
  assign n19009 = ~n1180 ;
  assign n1329 = n19009 & n1181 ;
  assign n1330 = n177 & n1329 ;
  assign n1331 = n1186 & n1330 ;
  assign n1332 = n1186 | n1330 ;
  assign n19010 = ~n1331 ;
  assign n1333 = n19010 & n1332 ;
  assign n19011 = ~n1333 ;
  assign n1334 = n1328 & n19011 ;
  assign n1335 = n1327 | n1334 ;
  assign n1336 = x74 & n1335 ;
  assign n1337 = x74 | n1335 ;
  assign n19012 = ~n1189 ;
  assign n1338 = n19012 & n1190 ;
  assign n1339 = n177 & n1338 ;
  assign n1340 = n1195 & n1339 ;
  assign n1341 = n1195 | n1339 ;
  assign n19013 = ~n1340 ;
  assign n1342 = n19013 & n1341 ;
  assign n19014 = ~n1342 ;
  assign n1343 = n1337 & n19014 ;
  assign n1344 = n1336 | n1343 ;
  assign n1345 = x75 & n1344 ;
  assign n1346 = x75 | n1344 ;
  assign n19015 = ~n1198 ;
  assign n1347 = n19015 & n1199 ;
  assign n1348 = n177 & n1347 ;
  assign n1349 = n1204 & n1348 ;
  assign n1350 = n1204 | n1348 ;
  assign n19016 = ~n1349 ;
  assign n1351 = n19016 & n1350 ;
  assign n19017 = ~n1351 ;
  assign n1352 = n1346 & n19017 ;
  assign n1353 = n1345 | n1352 ;
  assign n1354 = x76 & n1353 ;
  assign n1355 = x76 | n1353 ;
  assign n19018 = ~n1207 ;
  assign n1356 = n19018 & n1208 ;
  assign n1357 = n177 & n1356 ;
  assign n1358 = n1213 & n1357 ;
  assign n1359 = n1213 | n1357 ;
  assign n19019 = ~n1358 ;
  assign n1360 = n19019 & n1359 ;
  assign n19020 = ~n1360 ;
  assign n1361 = n1355 & n19020 ;
  assign n1362 = n1354 | n1361 ;
  assign n1363 = x77 & n1362 ;
  assign n1364 = x77 | n1362 ;
  assign n19021 = ~n1216 ;
  assign n1365 = n19021 & n1217 ;
  assign n1366 = n177 & n1365 ;
  assign n1367 = n1222 & n1366 ;
  assign n1368 = n1222 | n1366 ;
  assign n19022 = ~n1367 ;
  assign n1369 = n19022 & n1368 ;
  assign n19023 = ~n1369 ;
  assign n1370 = n1364 & n19023 ;
  assign n1371 = n1363 | n1370 ;
  assign n1372 = x78 & n1371 ;
  assign n1373 = x78 | n1371 ;
  assign n19024 = ~n1225 ;
  assign n1374 = n19024 & n1226 ;
  assign n1375 = n177 & n1374 ;
  assign n1376 = n1231 & n1375 ;
  assign n1377 = n1231 | n1375 ;
  assign n19025 = ~n1376 ;
  assign n1378 = n19025 & n1377 ;
  assign n19026 = ~n1378 ;
  assign n1379 = n1373 & n19026 ;
  assign n1380 = n1372 | n1379 ;
  assign n1382 = x79 & n1380 ;
  assign n19027 = ~n1382 ;
  assign n1383 = n1251 & n19027 ;
  assign n1252 = n1238 & n1243 ;
  assign n1253 = n21884 | n1252 ;
  assign n19028 = ~x80 ;
  assign n1254 = n19028 & n1253 ;
  assign n1381 = x79 | n1380 ;
  assign n19029 = ~n1254 ;
  assign n1384 = n19029 & n1381 ;
  assign n19030 = ~n1383 ;
  assign n1385 = n19030 & n1384 ;
  assign n1386 = n18493 | n1385 ;
  assign n19031 = ~n1253 ;
  assign n1387 = x80 & n19031 ;
  assign n1388 = n1386 | n1387 ;
  assign n1389 = n1381 & n19027 ;
  assign n176 = ~n1388 ;
  assign n1390 = n176 & n1389 ;
  assign n1391 = n1251 & n1390 ;
  assign n1392 = n1251 | n1390 ;
  assign n19033 = ~n1391 ;
  assign n1393 = n19033 & n1392 ;
  assign n19034 = ~x46 ;
  assign n1394 = n19034 & x64 ;
  assign n1395 = x65 | n1394 ;
  assign n1396 = x65 & n1394 ;
  assign n1397 = x64 & n176 ;
  assign n1398 = x47 & n1397 ;
  assign n1399 = x47 | n1397 ;
  assign n19035 = ~n1398 ;
  assign n1400 = n19035 & n1399 ;
  assign n19036 = ~n1396 ;
  assign n1401 = n19036 & n1400 ;
  assign n19037 = ~n1401 ;
  assign n1402 = n1395 & n19037 ;
  assign n1404 = x66 | n1402 ;
  assign n1403 = x66 & n1402 ;
  assign n1405 = n18987 & n1257 ;
  assign n1406 = n176 & n1405 ;
  assign n1407 = n1261 & n1406 ;
  assign n1408 = n1261 | n1406 ;
  assign n19038 = ~n1407 ;
  assign n1409 = n19038 & n1408 ;
  assign n19039 = ~n1403 ;
  assign n1410 = n19039 & n1409 ;
  assign n19040 = ~n1410 ;
  assign n1411 = n1404 & n19040 ;
  assign n1412 = x67 | n1411 ;
  assign n1413 = x67 & n1411 ;
  assign n19041 = ~n1264 ;
  assign n1414 = n19041 & n1265 ;
  assign n1415 = n176 & n1414 ;
  assign n1416 = n1270 & n1415 ;
  assign n1417 = n1270 | n1415 ;
  assign n19042 = ~n1416 ;
  assign n1418 = n19042 & n1417 ;
  assign n19043 = ~n1413 ;
  assign n1419 = n19043 & n1418 ;
  assign n19044 = ~n1419 ;
  assign n1420 = n1412 & n19044 ;
  assign n1421 = x68 | n1420 ;
  assign n1422 = x68 & n1420 ;
  assign n19045 = ~n1273 ;
  assign n1423 = n19045 & n1274 ;
  assign n1424 = n176 & n1423 ;
  assign n1425 = n1279 & n1424 ;
  assign n1426 = n1279 | n1424 ;
  assign n19046 = ~n1425 ;
  assign n1427 = n19046 & n1426 ;
  assign n19047 = ~n1422 ;
  assign n1428 = n19047 & n1427 ;
  assign n19048 = ~n1428 ;
  assign n1429 = n1421 & n19048 ;
  assign n1430 = x69 | n1429 ;
  assign n1431 = x69 & n1429 ;
  assign n19049 = ~n1282 ;
  assign n1432 = n19049 & n1283 ;
  assign n1433 = n176 & n1432 ;
  assign n1434 = n18996 & n1433 ;
  assign n19050 = ~n1433 ;
  assign n1435 = n1288 & n19050 ;
  assign n1436 = n1434 | n1435 ;
  assign n19051 = ~n1431 ;
  assign n1437 = n19051 & n1436 ;
  assign n19052 = ~n1437 ;
  assign n1438 = n1430 & n19052 ;
  assign n1439 = x70 | n1438 ;
  assign n1440 = x70 & n1438 ;
  assign n19053 = ~n1291 ;
  assign n1441 = n19053 & n1292 ;
  assign n1442 = n176 & n1441 ;
  assign n1443 = n1297 & n1442 ;
  assign n1444 = n1297 | n1442 ;
  assign n19054 = ~n1443 ;
  assign n1445 = n19054 & n1444 ;
  assign n19055 = ~n1440 ;
  assign n1446 = n19055 & n1445 ;
  assign n19056 = ~n1446 ;
  assign n1447 = n1439 & n19056 ;
  assign n1448 = x71 | n1447 ;
  assign n1449 = x71 & n1447 ;
  assign n19057 = ~n1300 ;
  assign n1450 = n19057 & n1301 ;
  assign n1451 = n176 & n1450 ;
  assign n1452 = n1306 & n1451 ;
  assign n1453 = n1306 | n1451 ;
  assign n19058 = ~n1452 ;
  assign n1454 = n19058 & n1453 ;
  assign n19059 = ~n1449 ;
  assign n1455 = n19059 & n1454 ;
  assign n19060 = ~n1455 ;
  assign n1456 = n1448 & n19060 ;
  assign n1457 = x72 | n1456 ;
  assign n1458 = x72 & n1456 ;
  assign n19061 = ~n1309 ;
  assign n1459 = n19061 & n1310 ;
  assign n1460 = n176 & n1459 ;
  assign n1461 = n1315 & n1460 ;
  assign n1462 = n1315 | n1460 ;
  assign n19062 = ~n1461 ;
  assign n1463 = n19062 & n1462 ;
  assign n19063 = ~n1458 ;
  assign n1464 = n19063 & n1463 ;
  assign n19064 = ~n1464 ;
  assign n1465 = n1457 & n19064 ;
  assign n1466 = x73 | n1465 ;
  assign n1467 = x73 & n1465 ;
  assign n19065 = ~n1318 ;
  assign n1468 = n19065 & n1319 ;
  assign n1469 = n176 & n1468 ;
  assign n1470 = n1324 & n1469 ;
  assign n1471 = n1324 | n1469 ;
  assign n19066 = ~n1470 ;
  assign n1472 = n19066 & n1471 ;
  assign n19067 = ~n1467 ;
  assign n1473 = n19067 & n1472 ;
  assign n19068 = ~n1473 ;
  assign n1474 = n1466 & n19068 ;
  assign n1475 = x74 | n1474 ;
  assign n1476 = x74 & n1474 ;
  assign n19069 = ~n1327 ;
  assign n1477 = n19069 & n1328 ;
  assign n1478 = n176 & n1477 ;
  assign n1479 = n1333 & n1478 ;
  assign n1480 = n1333 | n1478 ;
  assign n19070 = ~n1479 ;
  assign n1481 = n19070 & n1480 ;
  assign n19071 = ~n1476 ;
  assign n1482 = n19071 & n1481 ;
  assign n19072 = ~n1482 ;
  assign n1483 = n1475 & n19072 ;
  assign n1484 = x75 | n1483 ;
  assign n1485 = x75 & n1483 ;
  assign n19073 = ~n1336 ;
  assign n1486 = n19073 & n1337 ;
  assign n1487 = n176 & n1486 ;
  assign n1488 = n1342 & n1487 ;
  assign n1489 = n1342 | n1487 ;
  assign n19074 = ~n1488 ;
  assign n1490 = n19074 & n1489 ;
  assign n19075 = ~n1485 ;
  assign n1491 = n19075 & n1490 ;
  assign n19076 = ~n1491 ;
  assign n1492 = n1484 & n19076 ;
  assign n1493 = x76 | n1492 ;
  assign n1494 = x76 & n1492 ;
  assign n19077 = ~n1345 ;
  assign n1495 = n19077 & n1346 ;
  assign n1496 = n176 & n1495 ;
  assign n1497 = n1351 & n1496 ;
  assign n1498 = n1351 | n1496 ;
  assign n19078 = ~n1497 ;
  assign n1499 = n19078 & n1498 ;
  assign n19079 = ~n1494 ;
  assign n1500 = n19079 & n1499 ;
  assign n19080 = ~n1500 ;
  assign n1501 = n1493 & n19080 ;
  assign n1502 = x77 | n1501 ;
  assign n1503 = x77 & n1501 ;
  assign n19081 = ~n1354 ;
  assign n1504 = n19081 & n1355 ;
  assign n1505 = n176 & n1504 ;
  assign n1506 = n1360 & n1505 ;
  assign n1507 = n1360 | n1505 ;
  assign n19082 = ~n1506 ;
  assign n1508 = n19082 & n1507 ;
  assign n19083 = ~n1503 ;
  assign n1509 = n19083 & n1508 ;
  assign n19084 = ~n1509 ;
  assign n1510 = n1502 & n19084 ;
  assign n1511 = x78 | n1510 ;
  assign n1512 = x78 & n1510 ;
  assign n19085 = ~n1363 ;
  assign n1513 = n19085 & n1364 ;
  assign n1514 = n176 & n1513 ;
  assign n1515 = n1369 & n1514 ;
  assign n1516 = n1369 | n1514 ;
  assign n19086 = ~n1515 ;
  assign n1517 = n19086 & n1516 ;
  assign n19087 = ~n1512 ;
  assign n1518 = n19087 & n1517 ;
  assign n19088 = ~n1518 ;
  assign n1519 = n1511 & n19088 ;
  assign n1520 = x79 | n1519 ;
  assign n1521 = x79 & n1519 ;
  assign n19089 = ~n1372 ;
  assign n1522 = n19089 & n1373 ;
  assign n1523 = n176 & n1522 ;
  assign n1524 = n1378 & n1523 ;
  assign n1525 = n1378 | n1523 ;
  assign n19090 = ~n1524 ;
  assign n1526 = n19090 & n1525 ;
  assign n19091 = ~n1521 ;
  assign n1527 = n19091 & n1526 ;
  assign n19092 = ~n1527 ;
  assign n1528 = n1520 & n19092 ;
  assign n1529 = x80 | n1528 ;
  assign n1530 = x80 & n1528 ;
  assign n19093 = ~n1530 ;
  assign n1531 = n1393 & n19093 ;
  assign n19094 = ~n1531 ;
  assign n1532 = n1529 & n19094 ;
  assign n1534 = x81 & n1532 ;
  assign n1535 = n18488 | n1534 ;
  assign n1533 = x81 | n1532 ;
  assign n1536 = n1252 & n1386 ;
  assign n1537 = n21884 | n1536 ;
  assign n19095 = ~n1537 ;
  assign n1539 = n1533 & n19095 ;
  assign n1540 = n1535 | n1539 ;
  assign n1541 = n1529 & n19093 ;
  assign n175 = ~n1540 ;
  assign n1542 = n175 & n1541 ;
  assign n1543 = n1393 & n1542 ;
  assign n1544 = n1393 | n1542 ;
  assign n19097 = ~n1543 ;
  assign n1545 = n19097 & n1544 ;
  assign n1538 = x82 & n19095 ;
  assign n1697 = n18483 | n1538 ;
  assign n19098 = ~x45 ;
  assign n1546 = n19098 & x64 ;
  assign n1547 = x65 | n1546 ;
  assign n1548 = x65 & n1546 ;
  assign n1549 = x64 & n175 ;
  assign n1550 = x46 & n1549 ;
  assign n1551 = x46 | n1549 ;
  assign n19099 = ~n1550 ;
  assign n1552 = n19099 & n1551 ;
  assign n19100 = ~n1548 ;
  assign n1553 = n19100 & n1552 ;
  assign n19101 = ~n1553 ;
  assign n1554 = n1547 & n19101 ;
  assign n1556 = x66 | n1554 ;
  assign n1555 = x66 & n1554 ;
  assign n1557 = n1395 & n19036 ;
  assign n1558 = n175 & n1557 ;
  assign n1559 = n1400 & n1558 ;
  assign n1560 = n1400 | n1558 ;
  assign n19102 = ~n1559 ;
  assign n1561 = n19102 & n1560 ;
  assign n19103 = ~n1555 ;
  assign n1562 = n19103 & n1561 ;
  assign n19104 = ~n1562 ;
  assign n1563 = n1556 & n19104 ;
  assign n1564 = x67 & n1563 ;
  assign n1565 = x67 | n1563 ;
  assign n1566 = n1404 & n175 ;
  assign n1567 = n1410 & n1566 ;
  assign n1568 = n19039 & n1566 ;
  assign n1569 = n1409 | n1568 ;
  assign n19105 = ~n1567 ;
  assign n1570 = n19105 & n1569 ;
  assign n19106 = ~n1570 ;
  assign n1571 = n1565 & n19106 ;
  assign n1572 = n1564 | n1571 ;
  assign n1573 = x68 & n1572 ;
  assign n1574 = x68 | n1572 ;
  assign n1575 = n1412 & n175 ;
  assign n1576 = n1419 & n1575 ;
  assign n1577 = n19043 & n1575 ;
  assign n1578 = n1418 | n1577 ;
  assign n19107 = ~n1576 ;
  assign n1579 = n19107 & n1578 ;
  assign n19108 = ~n1579 ;
  assign n1580 = n1574 & n19108 ;
  assign n1581 = n1573 | n1580 ;
  assign n1582 = x69 & n1581 ;
  assign n1583 = x69 | n1581 ;
  assign n1584 = n1421 & n19047 ;
  assign n1585 = n175 & n1584 ;
  assign n19109 = ~n1427 ;
  assign n1586 = n19109 & n1585 ;
  assign n19110 = ~n1585 ;
  assign n1587 = n1427 & n19110 ;
  assign n1588 = n1586 | n1587 ;
  assign n19111 = ~n1588 ;
  assign n1589 = n1583 & n19111 ;
  assign n1590 = n1582 | n1589 ;
  assign n1591 = x70 & n1590 ;
  assign n1592 = x70 | n1590 ;
  assign n1593 = n1430 & n19051 ;
  assign n1594 = n175 & n1593 ;
  assign n19112 = ~n1436 ;
  assign n1595 = n19112 & n1594 ;
  assign n19113 = ~n1594 ;
  assign n1596 = n1436 & n19113 ;
  assign n1597 = n1595 | n1596 ;
  assign n19114 = ~n1597 ;
  assign n1598 = n1592 & n19114 ;
  assign n1599 = n1591 | n1598 ;
  assign n1600 = x71 & n1599 ;
  assign n1601 = x71 | n1599 ;
  assign n1602 = n1439 & n19055 ;
  assign n1603 = n175 & n1602 ;
  assign n1604 = n1445 & n1603 ;
  assign n1605 = n1445 | n1603 ;
  assign n19115 = ~n1604 ;
  assign n1606 = n19115 & n1605 ;
  assign n19116 = ~n1606 ;
  assign n1607 = n1601 & n19116 ;
  assign n1608 = n1600 | n1607 ;
  assign n1609 = x72 & n1608 ;
  assign n1610 = x72 | n1608 ;
  assign n1611 = n1448 & n19059 ;
  assign n1612 = n175 & n1611 ;
  assign n1613 = n1454 & n1612 ;
  assign n1614 = n1454 | n1612 ;
  assign n19117 = ~n1613 ;
  assign n1615 = n19117 & n1614 ;
  assign n19118 = ~n1615 ;
  assign n1616 = n1610 & n19118 ;
  assign n1617 = n1609 | n1616 ;
  assign n1618 = x73 & n1617 ;
  assign n1619 = x73 | n1617 ;
  assign n1620 = n1457 & n19063 ;
  assign n1621 = n175 & n1620 ;
  assign n1622 = n1463 & n1621 ;
  assign n1623 = n1463 | n1621 ;
  assign n19119 = ~n1622 ;
  assign n1624 = n19119 & n1623 ;
  assign n19120 = ~n1624 ;
  assign n1625 = n1619 & n19120 ;
  assign n1626 = n1618 | n1625 ;
  assign n1627 = x74 & n1626 ;
  assign n1628 = x74 | n1626 ;
  assign n1629 = n1466 & n19067 ;
  assign n1630 = n175 & n1629 ;
  assign n1631 = n1472 & n1630 ;
  assign n1632 = n1472 | n1630 ;
  assign n19121 = ~n1631 ;
  assign n1633 = n19121 & n1632 ;
  assign n19122 = ~n1633 ;
  assign n1634 = n1628 & n19122 ;
  assign n1635 = n1627 | n1634 ;
  assign n1636 = x75 & n1635 ;
  assign n1637 = x75 | n1635 ;
  assign n1638 = n1475 & n19071 ;
  assign n1639 = n175 & n1638 ;
  assign n1640 = n1481 & n1639 ;
  assign n1641 = n1481 | n1639 ;
  assign n19123 = ~n1640 ;
  assign n1642 = n19123 & n1641 ;
  assign n19124 = ~n1642 ;
  assign n1643 = n1637 & n19124 ;
  assign n1644 = n1636 | n1643 ;
  assign n1645 = x76 & n1644 ;
  assign n1646 = x76 | n1644 ;
  assign n1647 = n1484 & n19075 ;
  assign n1648 = n175 & n1647 ;
  assign n1649 = n1490 & n1648 ;
  assign n1650 = n1490 | n1648 ;
  assign n19125 = ~n1649 ;
  assign n1651 = n19125 & n1650 ;
  assign n19126 = ~n1651 ;
  assign n1652 = n1646 & n19126 ;
  assign n1653 = n1645 | n1652 ;
  assign n1654 = x77 & n1653 ;
  assign n1655 = x77 | n1653 ;
  assign n1656 = n1493 & n19079 ;
  assign n1657 = n175 & n1656 ;
  assign n1658 = n1499 & n1657 ;
  assign n1659 = n1499 | n1657 ;
  assign n19127 = ~n1658 ;
  assign n1660 = n19127 & n1659 ;
  assign n19128 = ~n1660 ;
  assign n1661 = n1655 & n19128 ;
  assign n1662 = n1654 | n1661 ;
  assign n1663 = x78 & n1662 ;
  assign n1664 = x78 | n1662 ;
  assign n1665 = n1502 & n19083 ;
  assign n1666 = n175 & n1665 ;
  assign n1667 = n1508 & n1666 ;
  assign n1668 = n1508 | n1666 ;
  assign n19129 = ~n1667 ;
  assign n1669 = n19129 & n1668 ;
  assign n19130 = ~n1669 ;
  assign n1670 = n1664 & n19130 ;
  assign n1671 = n1663 | n1670 ;
  assign n1672 = x79 & n1671 ;
  assign n1673 = x79 | n1671 ;
  assign n1674 = n1511 & n19087 ;
  assign n1675 = n175 & n1674 ;
  assign n1676 = n1517 & n1675 ;
  assign n1677 = n1517 | n1675 ;
  assign n19131 = ~n1676 ;
  assign n1678 = n19131 & n1677 ;
  assign n19132 = ~n1678 ;
  assign n1679 = n1673 & n19132 ;
  assign n1680 = n1672 | n1679 ;
  assign n1681 = x80 & n1680 ;
  assign n1682 = x80 | n1680 ;
  assign n1683 = n1520 & n19091 ;
  assign n1684 = n175 & n1683 ;
  assign n1685 = n1526 & n1684 ;
  assign n1686 = n1526 | n1684 ;
  assign n19133 = ~n1685 ;
  assign n1687 = n19133 & n1686 ;
  assign n19134 = ~n1687 ;
  assign n1688 = n1682 & n19134 ;
  assign n1689 = n1681 | n1688 ;
  assign n1690 = x81 & n1689 ;
  assign n19135 = ~n1690 ;
  assign n1691 = n1545 & n19135 ;
  assign n1694 = x81 | n1689 ;
  assign n1692 = n1535 & n1536 ;
  assign n1693 = n21884 | n1692 ;
  assign n19136 = ~x82 ;
  assign n1695 = n19136 & n1693 ;
  assign n19137 = ~n1695 ;
  assign n1696 = n1694 & n19137 ;
  assign n19138 = ~n1691 ;
  assign n1698 = n19138 & n1696 ;
  assign n1699 = n1697 | n1698 ;
  assign n1701 = n19135 & n1694 ;
  assign n174 = ~n1699 ;
  assign n1702 = n174 & n1701 ;
  assign n1703 = n1545 & n1702 ;
  assign n1704 = n1545 | n1702 ;
  assign n19140 = ~n1703 ;
  assign n1705 = n19140 & n1704 ;
  assign n19141 = ~x44 ;
  assign n1708 = n19141 & x64 ;
  assign n1709 = x65 | n1708 ;
  assign n1710 = x65 & n1708 ;
  assign n1711 = x64 & n174 ;
  assign n1712 = x45 & n1711 ;
  assign n1713 = x45 | n1711 ;
  assign n19142 = ~n1712 ;
  assign n1714 = n19142 & n1713 ;
  assign n19143 = ~n1710 ;
  assign n1715 = n19143 & n1714 ;
  assign n19144 = ~n1715 ;
  assign n1716 = n1709 & n19144 ;
  assign n1718 = x66 | n1716 ;
  assign n1717 = x66 & n1716 ;
  assign n1719 = n1547 & n19100 ;
  assign n1720 = n174 & n1719 ;
  assign n1721 = n1552 & n1720 ;
  assign n1722 = n1552 | n1720 ;
  assign n19145 = ~n1721 ;
  assign n1723 = n19145 & n1722 ;
  assign n19146 = ~n1717 ;
  assign n1724 = n19146 & n1723 ;
  assign n19147 = ~n1724 ;
  assign n1725 = n1718 & n19147 ;
  assign n1726 = x67 & n1725 ;
  assign n1727 = x67 | n1725 ;
  assign n1728 = n1556 & n174 ;
  assign n1729 = n1562 & n1728 ;
  assign n1730 = n19103 & n1728 ;
  assign n1731 = n1561 | n1730 ;
  assign n19148 = ~n1729 ;
  assign n1732 = n19148 & n1731 ;
  assign n19149 = ~n1732 ;
  assign n1733 = n1727 & n19149 ;
  assign n1734 = n1726 | n1733 ;
  assign n1735 = x68 | n1734 ;
  assign n1736 = x68 & n1734 ;
  assign n1737 = n1564 | n1699 ;
  assign n19150 = ~n1737 ;
  assign n1739 = n1571 & n19150 ;
  assign n1738 = n1565 & n19150 ;
  assign n19151 = ~n1738 ;
  assign n1740 = n1570 & n19151 ;
  assign n1741 = n1739 | n1740 ;
  assign n19152 = ~n1736 ;
  assign n1742 = n19152 & n1741 ;
  assign n19153 = ~n1742 ;
  assign n1743 = n1735 & n19153 ;
  assign n1744 = x69 | n1743 ;
  assign n1745 = x69 & n1743 ;
  assign n19154 = ~n1573 ;
  assign n1746 = n19154 & n1574 ;
  assign n1747 = n174 & n1746 ;
  assign n1748 = n1579 & n1747 ;
  assign n1749 = n1579 | n1747 ;
  assign n19155 = ~n1748 ;
  assign n1750 = n19155 & n1749 ;
  assign n19156 = ~n1745 ;
  assign n1751 = n19156 & n1750 ;
  assign n19157 = ~n1751 ;
  assign n1752 = n1744 & n19157 ;
  assign n1753 = x70 | n1752 ;
  assign n1754 = x70 & n1752 ;
  assign n19158 = ~n1582 ;
  assign n1755 = n19158 & n1583 ;
  assign n1756 = n174 & n1755 ;
  assign n1757 = n1588 & n1756 ;
  assign n1758 = n1588 | n1756 ;
  assign n19159 = ~n1757 ;
  assign n1759 = n19159 & n1758 ;
  assign n19160 = ~n1754 ;
  assign n1760 = n19160 & n1759 ;
  assign n19161 = ~n1760 ;
  assign n1761 = n1753 & n19161 ;
  assign n1762 = x71 | n1761 ;
  assign n1763 = x71 & n1761 ;
  assign n19162 = ~n1591 ;
  assign n1764 = n19162 & n1592 ;
  assign n1765 = n174 & n1764 ;
  assign n1766 = n1597 & n1765 ;
  assign n1767 = n1597 | n1765 ;
  assign n19163 = ~n1766 ;
  assign n1768 = n19163 & n1767 ;
  assign n19164 = ~n1763 ;
  assign n1769 = n19164 & n1768 ;
  assign n19165 = ~n1769 ;
  assign n1770 = n1762 & n19165 ;
  assign n1771 = x72 | n1770 ;
  assign n1772 = x72 & n1770 ;
  assign n19166 = ~n1600 ;
  assign n1773 = n19166 & n1601 ;
  assign n1774 = n174 & n1773 ;
  assign n1775 = n1606 & n1774 ;
  assign n1776 = n1606 | n1774 ;
  assign n19167 = ~n1775 ;
  assign n1777 = n19167 & n1776 ;
  assign n19168 = ~n1772 ;
  assign n1778 = n19168 & n1777 ;
  assign n19169 = ~n1778 ;
  assign n1779 = n1771 & n19169 ;
  assign n1780 = x73 | n1779 ;
  assign n1781 = x73 & n1779 ;
  assign n19170 = ~n1609 ;
  assign n1782 = n19170 & n1610 ;
  assign n1783 = n174 & n1782 ;
  assign n1784 = n1615 & n1783 ;
  assign n1785 = n1615 | n1783 ;
  assign n19171 = ~n1784 ;
  assign n1786 = n19171 & n1785 ;
  assign n19172 = ~n1781 ;
  assign n1787 = n19172 & n1786 ;
  assign n19173 = ~n1787 ;
  assign n1788 = n1780 & n19173 ;
  assign n1789 = x74 | n1788 ;
  assign n1790 = x74 & n1788 ;
  assign n19174 = ~n1618 ;
  assign n1791 = n19174 & n1619 ;
  assign n1792 = n174 & n1791 ;
  assign n1793 = n1624 & n1792 ;
  assign n1794 = n1624 | n1792 ;
  assign n19175 = ~n1793 ;
  assign n1795 = n19175 & n1794 ;
  assign n19176 = ~n1790 ;
  assign n1796 = n19176 & n1795 ;
  assign n19177 = ~n1796 ;
  assign n1797 = n1789 & n19177 ;
  assign n1798 = x75 | n1797 ;
  assign n1799 = x75 & n1797 ;
  assign n19178 = ~n1627 ;
  assign n1800 = n19178 & n1628 ;
  assign n1801 = n174 & n1800 ;
  assign n1802 = n1633 & n1801 ;
  assign n1803 = n1633 | n1801 ;
  assign n19179 = ~n1802 ;
  assign n1804 = n19179 & n1803 ;
  assign n19180 = ~n1799 ;
  assign n1805 = n19180 & n1804 ;
  assign n19181 = ~n1805 ;
  assign n1806 = n1798 & n19181 ;
  assign n1807 = x76 | n1806 ;
  assign n1808 = x76 & n1806 ;
  assign n19182 = ~n1636 ;
  assign n1809 = n19182 & n1637 ;
  assign n1810 = n174 & n1809 ;
  assign n1811 = n1642 & n1810 ;
  assign n1812 = n1642 | n1810 ;
  assign n19183 = ~n1811 ;
  assign n1813 = n19183 & n1812 ;
  assign n19184 = ~n1808 ;
  assign n1814 = n19184 & n1813 ;
  assign n19185 = ~n1814 ;
  assign n1815 = n1807 & n19185 ;
  assign n1816 = x77 | n1815 ;
  assign n1817 = x77 & n1815 ;
  assign n19186 = ~n1645 ;
  assign n1818 = n19186 & n1646 ;
  assign n1819 = n174 & n1818 ;
  assign n1820 = n1651 & n1819 ;
  assign n1821 = n1651 | n1819 ;
  assign n19187 = ~n1820 ;
  assign n1822 = n19187 & n1821 ;
  assign n19188 = ~n1817 ;
  assign n1823 = n19188 & n1822 ;
  assign n19189 = ~n1823 ;
  assign n1824 = n1816 & n19189 ;
  assign n1825 = x78 | n1824 ;
  assign n1826 = x78 & n1824 ;
  assign n19190 = ~n1654 ;
  assign n1827 = n19190 & n1655 ;
  assign n1828 = n174 & n1827 ;
  assign n1829 = n1660 & n1828 ;
  assign n1830 = n1660 | n1828 ;
  assign n19191 = ~n1829 ;
  assign n1831 = n19191 & n1830 ;
  assign n19192 = ~n1826 ;
  assign n1832 = n19192 & n1831 ;
  assign n19193 = ~n1832 ;
  assign n1833 = n1825 & n19193 ;
  assign n1834 = x79 | n1833 ;
  assign n1835 = x79 & n1833 ;
  assign n19194 = ~n1663 ;
  assign n1836 = n19194 & n1664 ;
  assign n1837 = n174 & n1836 ;
  assign n1838 = n1669 & n1837 ;
  assign n1839 = n1669 | n1837 ;
  assign n19195 = ~n1838 ;
  assign n1840 = n19195 & n1839 ;
  assign n19196 = ~n1835 ;
  assign n1841 = n19196 & n1840 ;
  assign n19197 = ~n1841 ;
  assign n1842 = n1834 & n19197 ;
  assign n1843 = x80 | n1842 ;
  assign n1844 = x80 & n1842 ;
  assign n19198 = ~n1672 ;
  assign n1845 = n19198 & n1673 ;
  assign n1846 = n174 & n1845 ;
  assign n1847 = n1678 & n1846 ;
  assign n1848 = n1678 | n1846 ;
  assign n19199 = ~n1847 ;
  assign n1849 = n19199 & n1848 ;
  assign n19200 = ~n1844 ;
  assign n1850 = n19200 & n1849 ;
  assign n19201 = ~n1850 ;
  assign n1851 = n1843 & n19201 ;
  assign n1852 = x81 | n1851 ;
  assign n1853 = x81 & n1851 ;
  assign n19202 = ~n1681 ;
  assign n1854 = n19202 & n1682 ;
  assign n1855 = n174 & n1854 ;
  assign n1856 = n1687 & n1855 ;
  assign n1857 = n1687 | n1855 ;
  assign n19203 = ~n1856 ;
  assign n1858 = n19203 & n1857 ;
  assign n19204 = ~n1853 ;
  assign n1859 = n19204 & n1858 ;
  assign n19205 = ~n1859 ;
  assign n1860 = n1852 & n19205 ;
  assign n1862 = x82 & n1860 ;
  assign n19206 = ~n1862 ;
  assign n1863 = n1705 & n19206 ;
  assign n1700 = n1692 & n1699 ;
  assign n1706 = n21884 | n1700 ;
  assign n19207 = ~x83 ;
  assign n1707 = n19207 & n1706 ;
  assign n1861 = x82 | n1860 ;
  assign n19208 = ~n1707 ;
  assign n1864 = n19208 & n1861 ;
  assign n19209 = ~n1863 ;
  assign n1865 = n19209 & n1864 ;
  assign n1866 = n18478 | n1865 ;
  assign n19210 = ~n1706 ;
  assign n1867 = x83 & n19210 ;
  assign n1868 = n1866 | n1867 ;
  assign n1869 = n1861 & n19206 ;
  assign n173 = ~n1868 ;
  assign n1870 = n173 & n1869 ;
  assign n1871 = n1705 & n1870 ;
  assign n1872 = n1705 | n1870 ;
  assign n19212 = ~n1871 ;
  assign n1873 = n19212 & n1872 ;
  assign n1874 = n1700 & n1866 ;
  assign n1875 = n21884 | n1874 ;
  assign n19213 = ~n18478 ;
  assign n1877 = n19213 & n1875 ;
  assign n19214 = ~x43 ;
  assign n1878 = n19214 & x64 ;
  assign n1879 = x65 | n1878 ;
  assign n1880 = x65 & n1878 ;
  assign n1881 = x64 & n173 ;
  assign n1882 = x44 & n1881 ;
  assign n1883 = x44 | n1881 ;
  assign n19215 = ~n1882 ;
  assign n1884 = n19215 & n1883 ;
  assign n19216 = ~n1880 ;
  assign n1885 = n19216 & n1884 ;
  assign n19217 = ~n1885 ;
  assign n1886 = n1879 & n19217 ;
  assign n1888 = x66 | n1886 ;
  assign n1887 = x66 & n1886 ;
  assign n1889 = n1709 & n19143 ;
  assign n1890 = n173 & n1889 ;
  assign n1891 = n1714 & n1890 ;
  assign n1892 = n1714 | n1890 ;
  assign n19218 = ~n1891 ;
  assign n1893 = n19218 & n1892 ;
  assign n19219 = ~n1887 ;
  assign n1894 = n19219 & n1893 ;
  assign n19220 = ~n1894 ;
  assign n1895 = n1888 & n19220 ;
  assign n1896 = x67 & n1895 ;
  assign n1897 = x67 | n1895 ;
  assign n1898 = n1718 & n173 ;
  assign n1899 = n1724 & n1898 ;
  assign n1900 = n19146 & n1898 ;
  assign n1901 = n1723 | n1900 ;
  assign n19221 = ~n1899 ;
  assign n1902 = n19221 & n1901 ;
  assign n19222 = ~n1902 ;
  assign n1903 = n1897 & n19222 ;
  assign n1904 = n1896 | n1903 ;
  assign n1905 = x68 | n1904 ;
  assign n1906 = x68 & n1904 ;
  assign n19223 = ~n1726 ;
  assign n1907 = n19223 & n1727 ;
  assign n1908 = n173 & n1907 ;
  assign n1909 = n1732 & n1908 ;
  assign n1910 = n1732 | n1908 ;
  assign n19224 = ~n1909 ;
  assign n1911 = n19224 & n1910 ;
  assign n19225 = ~n1906 ;
  assign n1912 = n19225 & n1911 ;
  assign n19226 = ~n1912 ;
  assign n1913 = n1905 & n19226 ;
  assign n1914 = x69 | n1913 ;
  assign n1915 = x69 & n1913 ;
  assign n1916 = n1735 & n19152 ;
  assign n1917 = n173 & n1916 ;
  assign n19227 = ~n1741 ;
  assign n1918 = n19227 & n1917 ;
  assign n19228 = ~n1917 ;
  assign n1919 = n1741 & n19228 ;
  assign n1920 = n1918 | n1919 ;
  assign n19229 = ~n1915 ;
  assign n1921 = n19229 & n1920 ;
  assign n19230 = ~n1921 ;
  assign n1922 = n1914 & n19230 ;
  assign n1923 = x70 | n1922 ;
  assign n1924 = x70 & n1922 ;
  assign n1925 = n1744 & n19156 ;
  assign n1926 = n173 & n1925 ;
  assign n1927 = n1750 & n1926 ;
  assign n1928 = n1750 | n1926 ;
  assign n19231 = ~n1927 ;
  assign n1929 = n19231 & n1928 ;
  assign n19232 = ~n1924 ;
  assign n1930 = n19232 & n1929 ;
  assign n19233 = ~n1930 ;
  assign n1931 = n1923 & n19233 ;
  assign n1932 = x71 | n1931 ;
  assign n1933 = x71 & n1931 ;
  assign n1934 = n1753 & n19160 ;
  assign n1935 = n173 & n1934 ;
  assign n1936 = n1759 & n1935 ;
  assign n1937 = n1759 | n1935 ;
  assign n19234 = ~n1936 ;
  assign n1938 = n19234 & n1937 ;
  assign n19235 = ~n1933 ;
  assign n1939 = n19235 & n1938 ;
  assign n19236 = ~n1939 ;
  assign n1940 = n1932 & n19236 ;
  assign n1941 = x72 | n1940 ;
  assign n1942 = x72 & n1940 ;
  assign n1943 = n1762 & n19164 ;
  assign n1944 = n173 & n1943 ;
  assign n1945 = n1768 & n1944 ;
  assign n1946 = n1768 | n1944 ;
  assign n19237 = ~n1945 ;
  assign n1947 = n19237 & n1946 ;
  assign n19238 = ~n1942 ;
  assign n1948 = n19238 & n1947 ;
  assign n19239 = ~n1948 ;
  assign n1949 = n1941 & n19239 ;
  assign n1950 = x73 | n1949 ;
  assign n1951 = x73 & n1949 ;
  assign n1952 = n1771 & n19168 ;
  assign n1953 = n173 & n1952 ;
  assign n1954 = n1777 & n1953 ;
  assign n1955 = n1777 | n1953 ;
  assign n19240 = ~n1954 ;
  assign n1956 = n19240 & n1955 ;
  assign n19241 = ~n1951 ;
  assign n1957 = n19241 & n1956 ;
  assign n19242 = ~n1957 ;
  assign n1958 = n1950 & n19242 ;
  assign n1959 = x74 | n1958 ;
  assign n1960 = x74 & n1958 ;
  assign n1961 = n1780 & n19172 ;
  assign n1962 = n173 & n1961 ;
  assign n1963 = n1786 & n1962 ;
  assign n1964 = n1786 | n1962 ;
  assign n19243 = ~n1963 ;
  assign n1965 = n19243 & n1964 ;
  assign n19244 = ~n1960 ;
  assign n1966 = n19244 & n1965 ;
  assign n19245 = ~n1966 ;
  assign n1967 = n1959 & n19245 ;
  assign n1968 = x75 | n1967 ;
  assign n1969 = x75 & n1967 ;
  assign n1970 = n1789 & n19176 ;
  assign n1971 = n173 & n1970 ;
  assign n1972 = n1795 & n1971 ;
  assign n1973 = n1795 | n1971 ;
  assign n19246 = ~n1972 ;
  assign n1974 = n19246 & n1973 ;
  assign n19247 = ~n1969 ;
  assign n1975 = n19247 & n1974 ;
  assign n19248 = ~n1975 ;
  assign n1976 = n1968 & n19248 ;
  assign n1977 = x76 | n1976 ;
  assign n1978 = x76 & n1976 ;
  assign n1979 = n1798 & n19180 ;
  assign n1980 = n173 & n1979 ;
  assign n1981 = n1804 & n1980 ;
  assign n1982 = n1804 | n1980 ;
  assign n19249 = ~n1981 ;
  assign n1983 = n19249 & n1982 ;
  assign n19250 = ~n1978 ;
  assign n1984 = n19250 & n1983 ;
  assign n19251 = ~n1984 ;
  assign n1985 = n1977 & n19251 ;
  assign n1986 = x77 | n1985 ;
  assign n1987 = x77 & n1985 ;
  assign n1988 = n1807 & n19184 ;
  assign n1989 = n173 & n1988 ;
  assign n1990 = n1813 & n1989 ;
  assign n1991 = n1813 | n1989 ;
  assign n19252 = ~n1990 ;
  assign n1992 = n19252 & n1991 ;
  assign n19253 = ~n1987 ;
  assign n1993 = n19253 & n1992 ;
  assign n19254 = ~n1993 ;
  assign n1994 = n1986 & n19254 ;
  assign n1995 = x78 | n1994 ;
  assign n1996 = x78 & n1994 ;
  assign n1997 = n1816 & n19188 ;
  assign n1998 = n173 & n1997 ;
  assign n1999 = n1822 & n1998 ;
  assign n2000 = n1822 | n1998 ;
  assign n19255 = ~n1999 ;
  assign n2001 = n19255 & n2000 ;
  assign n19256 = ~n1996 ;
  assign n2002 = n19256 & n2001 ;
  assign n19257 = ~n2002 ;
  assign n2003 = n1995 & n19257 ;
  assign n2004 = x79 | n2003 ;
  assign n2005 = x79 & n2003 ;
  assign n2006 = n1825 & n19192 ;
  assign n2007 = n173 & n2006 ;
  assign n2008 = n1831 & n2007 ;
  assign n2009 = n1831 | n2007 ;
  assign n19258 = ~n2008 ;
  assign n2010 = n19258 & n2009 ;
  assign n19259 = ~n2005 ;
  assign n2011 = n19259 & n2010 ;
  assign n19260 = ~n2011 ;
  assign n2012 = n2004 & n19260 ;
  assign n2013 = x80 | n2012 ;
  assign n2014 = x80 & n2012 ;
  assign n2015 = n1834 & n19196 ;
  assign n2016 = n173 & n2015 ;
  assign n2017 = n1840 & n2016 ;
  assign n2018 = n1840 | n2016 ;
  assign n19261 = ~n2017 ;
  assign n2019 = n19261 & n2018 ;
  assign n19262 = ~n2014 ;
  assign n2020 = n19262 & n2019 ;
  assign n19263 = ~n2020 ;
  assign n2021 = n2013 & n19263 ;
  assign n2022 = x81 | n2021 ;
  assign n2023 = x81 & n2021 ;
  assign n2024 = n1843 & n19200 ;
  assign n2025 = n173 & n2024 ;
  assign n2026 = n1849 & n2025 ;
  assign n2027 = n1849 | n2025 ;
  assign n19264 = ~n2026 ;
  assign n2028 = n19264 & n2027 ;
  assign n19265 = ~n2023 ;
  assign n2029 = n19265 & n2028 ;
  assign n19266 = ~n2029 ;
  assign n2030 = n2022 & n19266 ;
  assign n2031 = x82 | n2030 ;
  assign n2032 = x82 & n2030 ;
  assign n2033 = n1852 & n19204 ;
  assign n2034 = n173 & n2033 ;
  assign n2035 = n1858 & n2034 ;
  assign n2036 = n1858 | n2034 ;
  assign n19267 = ~n2035 ;
  assign n2037 = n19267 & n2036 ;
  assign n19268 = ~n2032 ;
  assign n2038 = n19268 & n2037 ;
  assign n19269 = ~n2038 ;
  assign n2039 = n2031 & n19269 ;
  assign n2041 = x83 | n2039 ;
  assign n19270 = ~n1873 ;
  assign n2042 = n19270 & n2041 ;
  assign n2040 = x83 & n2039 ;
  assign n19271 = ~n1875 ;
  assign n1876 = x84 & n19271 ;
  assign n2043 = n18473 | n1876 ;
  assign n19272 = ~x84 ;
  assign n2044 = n19272 & n1875 ;
  assign n2045 = n2043 | n2044 ;
  assign n2046 = n2040 | n2045 ;
  assign n2047 = n2042 | n2046 ;
  assign n19273 = ~n1877 ;
  assign n2048 = n19273 & n2047 ;
  assign n19274 = ~n2040 ;
  assign n2049 = n19274 & n2041 ;
  assign n172 = ~n2048 ;
  assign n2050 = n172 & n2049 ;
  assign n2051 = n19270 & n2050 ;
  assign n19276 = ~n2050 ;
  assign n2052 = n1873 & n19276 ;
  assign n2053 = n2051 | n2052 ;
  assign n19277 = ~x42 ;
  assign n2054 = n19277 & x64 ;
  assign n2055 = x65 | n2054 ;
  assign n2056 = x64 & n172 ;
  assign n19278 = ~n2056 ;
  assign n2057 = x43 & n19278 ;
  assign n2058 = n1878 & n172 ;
  assign n2059 = n2057 | n2058 ;
  assign n2060 = x65 & n2054 ;
  assign n19279 = ~n2060 ;
  assign n2061 = n2059 & n19279 ;
  assign n19280 = ~n2061 ;
  assign n2062 = n2055 & n19280 ;
  assign n2063 = x66 | n2062 ;
  assign n2064 = x66 & n2062 ;
  assign n2065 = n1879 & n19216 ;
  assign n2066 = n172 & n2065 ;
  assign n2067 = n1884 & n2066 ;
  assign n2068 = n1884 | n2066 ;
  assign n19281 = ~n2067 ;
  assign n2069 = n19281 & n2068 ;
  assign n19282 = ~n2064 ;
  assign n2070 = n19282 & n2069 ;
  assign n19283 = ~n2070 ;
  assign n2071 = n2063 & n19283 ;
  assign n2072 = x67 & n2071 ;
  assign n2073 = x67 | n2071 ;
  assign n2074 = n1888 & n172 ;
  assign n2075 = n1894 & n2074 ;
  assign n2076 = n19219 & n2074 ;
  assign n2077 = n1893 | n2076 ;
  assign n19284 = ~n2075 ;
  assign n2078 = n19284 & n2077 ;
  assign n19285 = ~n2078 ;
  assign n2079 = n2073 & n19285 ;
  assign n2080 = n2072 | n2079 ;
  assign n2081 = x68 | n2080 ;
  assign n2082 = x68 & n2080 ;
  assign n19286 = ~n1896 ;
  assign n2083 = n19286 & n1897 ;
  assign n2084 = n172 & n2083 ;
  assign n2085 = n1902 & n2084 ;
  assign n2086 = n1902 | n2084 ;
  assign n19287 = ~n2085 ;
  assign n2087 = n19287 & n2086 ;
  assign n19288 = ~n2082 ;
  assign n2088 = n19288 & n2087 ;
  assign n19289 = ~n2088 ;
  assign n2089 = n2081 & n19289 ;
  assign n2090 = x69 | n2089 ;
  assign n2091 = x69 & n2089 ;
  assign n2092 = n1905 & n19225 ;
  assign n2093 = n172 & n2092 ;
  assign n19290 = ~n1911 ;
  assign n2094 = n19290 & n2093 ;
  assign n19291 = ~n2093 ;
  assign n2095 = n1911 & n19291 ;
  assign n2096 = n2094 | n2095 ;
  assign n19292 = ~n2091 ;
  assign n2097 = n19292 & n2096 ;
  assign n19293 = ~n2097 ;
  assign n2098 = n2090 & n19293 ;
  assign n2099 = x70 | n2098 ;
  assign n2100 = x70 & n2098 ;
  assign n2101 = n1914 & n19229 ;
  assign n2102 = n172 & n2101 ;
  assign n2103 = n1920 & n2102 ;
  assign n2104 = n1920 | n2102 ;
  assign n19294 = ~n2103 ;
  assign n2105 = n19294 & n2104 ;
  assign n19295 = ~n2100 ;
  assign n2106 = n19295 & n2105 ;
  assign n19296 = ~n2106 ;
  assign n2107 = n2099 & n19296 ;
  assign n2108 = x71 | n2107 ;
  assign n2109 = x71 & n2107 ;
  assign n2110 = n1923 & n19232 ;
  assign n2111 = n172 & n2110 ;
  assign n2112 = n1929 & n2111 ;
  assign n2113 = n1929 | n2111 ;
  assign n19297 = ~n2112 ;
  assign n2114 = n19297 & n2113 ;
  assign n19298 = ~n2109 ;
  assign n2115 = n19298 & n2114 ;
  assign n19299 = ~n2115 ;
  assign n2116 = n2108 & n19299 ;
  assign n2117 = x72 | n2116 ;
  assign n2118 = x72 & n2116 ;
  assign n2119 = n1932 & n19235 ;
  assign n2120 = n172 & n2119 ;
  assign n2121 = n1938 & n2120 ;
  assign n2122 = n1938 | n2120 ;
  assign n19300 = ~n2121 ;
  assign n2123 = n19300 & n2122 ;
  assign n19301 = ~n2118 ;
  assign n2124 = n19301 & n2123 ;
  assign n19302 = ~n2124 ;
  assign n2125 = n2117 & n19302 ;
  assign n2126 = x73 | n2125 ;
  assign n2127 = x73 & n2125 ;
  assign n2128 = n1941 & n19238 ;
  assign n2129 = n172 & n2128 ;
  assign n2130 = n1947 & n2129 ;
  assign n2131 = n1947 | n2129 ;
  assign n19303 = ~n2130 ;
  assign n2132 = n19303 & n2131 ;
  assign n19304 = ~n2127 ;
  assign n2133 = n19304 & n2132 ;
  assign n19305 = ~n2133 ;
  assign n2134 = n2126 & n19305 ;
  assign n2135 = x74 | n2134 ;
  assign n2136 = x74 & n2134 ;
  assign n2137 = n1950 & n19241 ;
  assign n2138 = n172 & n2137 ;
  assign n2139 = n1956 & n2138 ;
  assign n2140 = n1956 | n2138 ;
  assign n19306 = ~n2139 ;
  assign n2141 = n19306 & n2140 ;
  assign n19307 = ~n2136 ;
  assign n2142 = n19307 & n2141 ;
  assign n19308 = ~n2142 ;
  assign n2143 = n2135 & n19308 ;
  assign n2144 = x75 | n2143 ;
  assign n2145 = x75 & n2143 ;
  assign n2146 = n1959 & n19244 ;
  assign n2147 = n172 & n2146 ;
  assign n2148 = n1965 & n2147 ;
  assign n2149 = n1965 | n2147 ;
  assign n19309 = ~n2148 ;
  assign n2150 = n19309 & n2149 ;
  assign n19310 = ~n2145 ;
  assign n2151 = n19310 & n2150 ;
  assign n19311 = ~n2151 ;
  assign n2152 = n2144 & n19311 ;
  assign n2153 = x76 | n2152 ;
  assign n2154 = x76 & n2152 ;
  assign n2155 = n1968 & n19247 ;
  assign n2156 = n172 & n2155 ;
  assign n2157 = n1974 & n2156 ;
  assign n2158 = n1974 | n2156 ;
  assign n19312 = ~n2157 ;
  assign n2159 = n19312 & n2158 ;
  assign n19313 = ~n2154 ;
  assign n2160 = n19313 & n2159 ;
  assign n19314 = ~n2160 ;
  assign n2161 = n2153 & n19314 ;
  assign n2162 = x77 | n2161 ;
  assign n2163 = x77 & n2161 ;
  assign n2164 = n1977 & n19250 ;
  assign n2165 = n172 & n2164 ;
  assign n2166 = n1983 & n2165 ;
  assign n2167 = n1983 | n2165 ;
  assign n19315 = ~n2166 ;
  assign n2168 = n19315 & n2167 ;
  assign n19316 = ~n2163 ;
  assign n2169 = n19316 & n2168 ;
  assign n19317 = ~n2169 ;
  assign n2170 = n2162 & n19317 ;
  assign n2171 = x78 | n2170 ;
  assign n2172 = x78 & n2170 ;
  assign n2173 = n1986 & n19253 ;
  assign n2174 = n172 & n2173 ;
  assign n2175 = n1992 & n2174 ;
  assign n2176 = n1992 | n2174 ;
  assign n19318 = ~n2175 ;
  assign n2177 = n19318 & n2176 ;
  assign n19319 = ~n2172 ;
  assign n2178 = n19319 & n2177 ;
  assign n19320 = ~n2178 ;
  assign n2179 = n2171 & n19320 ;
  assign n2180 = x79 | n2179 ;
  assign n2181 = x79 & n2179 ;
  assign n2182 = n1995 & n19256 ;
  assign n2183 = n172 & n2182 ;
  assign n2184 = n2001 & n2183 ;
  assign n2185 = n2001 | n2183 ;
  assign n19321 = ~n2184 ;
  assign n2186 = n19321 & n2185 ;
  assign n19322 = ~n2181 ;
  assign n2187 = n19322 & n2186 ;
  assign n19323 = ~n2187 ;
  assign n2188 = n2180 & n19323 ;
  assign n2189 = x80 | n2188 ;
  assign n2190 = x80 & n2188 ;
  assign n2191 = n2004 & n19259 ;
  assign n2192 = n172 & n2191 ;
  assign n2193 = n2010 & n2192 ;
  assign n2194 = n2010 | n2192 ;
  assign n19324 = ~n2193 ;
  assign n2195 = n19324 & n2194 ;
  assign n19325 = ~n2190 ;
  assign n2196 = n19325 & n2195 ;
  assign n19326 = ~n2196 ;
  assign n2197 = n2189 & n19326 ;
  assign n2198 = x81 | n2197 ;
  assign n2199 = x81 & n2197 ;
  assign n2200 = n2013 & n19262 ;
  assign n2201 = n172 & n2200 ;
  assign n2202 = n2019 & n2201 ;
  assign n2203 = n2019 | n2201 ;
  assign n19327 = ~n2202 ;
  assign n2204 = n19327 & n2203 ;
  assign n19328 = ~n2199 ;
  assign n2205 = n19328 & n2204 ;
  assign n19329 = ~n2205 ;
  assign n2206 = n2198 & n19329 ;
  assign n2207 = x82 | n2206 ;
  assign n2208 = x82 & n2206 ;
  assign n2209 = n2022 & n19265 ;
  assign n2210 = n172 & n2209 ;
  assign n2211 = n2028 & n2210 ;
  assign n2212 = n2028 | n2210 ;
  assign n19330 = ~n2211 ;
  assign n2213 = n19330 & n2212 ;
  assign n19331 = ~n2208 ;
  assign n2214 = n19331 & n2213 ;
  assign n19332 = ~n2214 ;
  assign n2215 = n2207 & n19332 ;
  assign n2216 = x83 | n2215 ;
  assign n2217 = x83 & n2215 ;
  assign n2218 = n2031 & n19268 ;
  assign n2219 = n172 & n2218 ;
  assign n2220 = n2037 & n2219 ;
  assign n2221 = n2037 | n2219 ;
  assign n19333 = ~n2220 ;
  assign n2222 = n19333 & n2221 ;
  assign n19334 = ~n2217 ;
  assign n2223 = n19334 & n2222 ;
  assign n19335 = ~n2223 ;
  assign n2224 = n2216 & n19335 ;
  assign n2225 = x84 | n2224 ;
  assign n2226 = x84 & n2224 ;
  assign n19336 = ~n2226 ;
  assign n2227 = n2053 & n19336 ;
  assign n19337 = ~n2227 ;
  assign n2228 = n2225 & n19337 ;
  assign n2230 = x85 & n2228 ;
  assign n2231 = n18468 | n2230 ;
  assign n2229 = x85 | n2228 ;
  assign n2232 = n18478 & n1706 ;
  assign n2233 = n2047 & n2232 ;
  assign n2234 = n21884 | n2233 ;
  assign n19338 = ~n2234 ;
  assign n2235 = n2229 & n19338 ;
  assign n2236 = n2231 | n2235 ;
  assign n2237 = n2225 & n19336 ;
  assign n171 = ~n2236 ;
  assign n2238 = n171 & n2237 ;
  assign n19340 = ~n2053 ;
  assign n2239 = n19340 & n2238 ;
  assign n19341 = ~n2238 ;
  assign n2240 = n2053 & n19341 ;
  assign n2241 = n2239 | n2240 ;
  assign n19342 = ~x41 ;
  assign n2245 = n19342 & x64 ;
  assign n2247 = x65 | n2245 ;
  assign n2246 = x65 & n2245 ;
  assign n2248 = x64 & n171 ;
  assign n2249 = x42 & n2248 ;
  assign n2250 = x42 | n2248 ;
  assign n19343 = ~n2249 ;
  assign n2251 = n19343 & n2250 ;
  assign n19344 = ~n2246 ;
  assign n2252 = n19344 & n2251 ;
  assign n19345 = ~n2252 ;
  assign n2253 = n2247 & n19345 ;
  assign n2254 = x66 & n2253 ;
  assign n2255 = x66 | n2253 ;
  assign n2256 = n2055 & n171 ;
  assign n2257 = n2061 & n2256 ;
  assign n2258 = n19279 & n2256 ;
  assign n2259 = n2059 | n2258 ;
  assign n19346 = ~n2257 ;
  assign n2260 = n19346 & n2259 ;
  assign n19347 = ~n2260 ;
  assign n2261 = n2255 & n19347 ;
  assign n2262 = n2254 | n2261 ;
  assign n2263 = x67 & n2262 ;
  assign n2264 = x67 | n2262 ;
  assign n2265 = n2063 & n171 ;
  assign n2266 = n2070 & n2265 ;
  assign n2267 = n19282 & n2265 ;
  assign n2268 = n2069 | n2267 ;
  assign n19348 = ~n2266 ;
  assign n2269 = n19348 & n2268 ;
  assign n19349 = ~n2269 ;
  assign n2270 = n2264 & n19349 ;
  assign n2271 = n2263 | n2270 ;
  assign n2273 = x68 | n2271 ;
  assign n2272 = x68 & n2271 ;
  assign n19350 = ~n2072 ;
  assign n2274 = n19350 & n2073 ;
  assign n2275 = n171 & n2274 ;
  assign n2276 = n2078 & n2275 ;
  assign n2277 = n2078 | n2275 ;
  assign n19351 = ~n2276 ;
  assign n2278 = n19351 & n2277 ;
  assign n19352 = ~n2272 ;
  assign n2279 = n19352 & n2278 ;
  assign n19353 = ~n2279 ;
  assign n2280 = n2273 & n19353 ;
  assign n2281 = x69 | n2280 ;
  assign n2282 = x69 & n2280 ;
  assign n2283 = n2081 & n19288 ;
  assign n2284 = n171 & n2283 ;
  assign n19354 = ~n2087 ;
  assign n2285 = n19354 & n2284 ;
  assign n19355 = ~n2284 ;
  assign n2286 = n2087 & n19355 ;
  assign n2287 = n2285 | n2286 ;
  assign n19356 = ~n2282 ;
  assign n2288 = n19356 & n2287 ;
  assign n19357 = ~n2288 ;
  assign n2289 = n2281 & n19357 ;
  assign n2290 = x70 | n2289 ;
  assign n2291 = x70 & n2289 ;
  assign n2292 = n2090 & n19292 ;
  assign n2293 = n171 & n2292 ;
  assign n19358 = ~n2096 ;
  assign n2294 = n19358 & n2293 ;
  assign n19359 = ~n2293 ;
  assign n2295 = n2096 & n19359 ;
  assign n2296 = n2294 | n2295 ;
  assign n19360 = ~n2291 ;
  assign n2297 = n19360 & n2296 ;
  assign n19361 = ~n2297 ;
  assign n2298 = n2290 & n19361 ;
  assign n2299 = x71 | n2298 ;
  assign n2300 = x71 & n2298 ;
  assign n2301 = n2099 & n19295 ;
  assign n2302 = n171 & n2301 ;
  assign n2303 = n2105 & n2302 ;
  assign n2304 = n2105 | n2302 ;
  assign n19362 = ~n2303 ;
  assign n2305 = n19362 & n2304 ;
  assign n19363 = ~n2300 ;
  assign n2306 = n19363 & n2305 ;
  assign n19364 = ~n2306 ;
  assign n2307 = n2299 & n19364 ;
  assign n2308 = x72 | n2307 ;
  assign n2309 = x72 & n2307 ;
  assign n2310 = n2108 & n19298 ;
  assign n2311 = n171 & n2310 ;
  assign n2312 = n2114 & n2311 ;
  assign n2313 = n2114 | n2311 ;
  assign n19365 = ~n2312 ;
  assign n2314 = n19365 & n2313 ;
  assign n19366 = ~n2309 ;
  assign n2315 = n19366 & n2314 ;
  assign n19367 = ~n2315 ;
  assign n2316 = n2308 & n19367 ;
  assign n2317 = x73 | n2316 ;
  assign n2318 = x73 & n2316 ;
  assign n2319 = n2117 & n19301 ;
  assign n2320 = n171 & n2319 ;
  assign n2321 = n2123 & n2320 ;
  assign n2322 = n2123 | n2320 ;
  assign n19368 = ~n2321 ;
  assign n2323 = n19368 & n2322 ;
  assign n19369 = ~n2318 ;
  assign n2324 = n19369 & n2323 ;
  assign n19370 = ~n2324 ;
  assign n2325 = n2317 & n19370 ;
  assign n2326 = x74 | n2325 ;
  assign n2327 = x74 & n2325 ;
  assign n2328 = n2126 & n19304 ;
  assign n2329 = n171 & n2328 ;
  assign n2330 = n2132 & n2329 ;
  assign n2331 = n2132 | n2329 ;
  assign n19371 = ~n2330 ;
  assign n2332 = n19371 & n2331 ;
  assign n19372 = ~n2327 ;
  assign n2333 = n19372 & n2332 ;
  assign n19373 = ~n2333 ;
  assign n2334 = n2326 & n19373 ;
  assign n2335 = x75 | n2334 ;
  assign n2336 = x75 & n2334 ;
  assign n2337 = n2135 & n19307 ;
  assign n2338 = n171 & n2337 ;
  assign n2339 = n2141 & n2338 ;
  assign n2340 = n2141 | n2338 ;
  assign n19374 = ~n2339 ;
  assign n2341 = n19374 & n2340 ;
  assign n19375 = ~n2336 ;
  assign n2342 = n19375 & n2341 ;
  assign n19376 = ~n2342 ;
  assign n2343 = n2335 & n19376 ;
  assign n2344 = x76 | n2343 ;
  assign n2345 = x76 & n2343 ;
  assign n2346 = n2144 & n19310 ;
  assign n2347 = n171 & n2346 ;
  assign n2348 = n2150 & n2347 ;
  assign n2349 = n2150 | n2347 ;
  assign n19377 = ~n2348 ;
  assign n2350 = n19377 & n2349 ;
  assign n19378 = ~n2345 ;
  assign n2351 = n19378 & n2350 ;
  assign n19379 = ~n2351 ;
  assign n2352 = n2344 & n19379 ;
  assign n2353 = x77 | n2352 ;
  assign n2354 = x77 & n2352 ;
  assign n2355 = n2153 & n19313 ;
  assign n2356 = n171 & n2355 ;
  assign n2357 = n2159 & n2356 ;
  assign n2358 = n2159 | n2356 ;
  assign n19380 = ~n2357 ;
  assign n2359 = n19380 & n2358 ;
  assign n19381 = ~n2354 ;
  assign n2360 = n19381 & n2359 ;
  assign n19382 = ~n2360 ;
  assign n2361 = n2353 & n19382 ;
  assign n2362 = x78 | n2361 ;
  assign n2363 = x78 & n2361 ;
  assign n2364 = n2162 & n19316 ;
  assign n2365 = n171 & n2364 ;
  assign n2366 = n2168 & n2365 ;
  assign n2367 = n2168 | n2365 ;
  assign n19383 = ~n2366 ;
  assign n2368 = n19383 & n2367 ;
  assign n19384 = ~n2363 ;
  assign n2369 = n19384 & n2368 ;
  assign n19385 = ~n2369 ;
  assign n2370 = n2362 & n19385 ;
  assign n2371 = x79 | n2370 ;
  assign n2372 = x79 & n2370 ;
  assign n2373 = n2171 & n19319 ;
  assign n2374 = n171 & n2373 ;
  assign n2375 = n2177 & n2374 ;
  assign n2376 = n2177 | n2374 ;
  assign n19386 = ~n2375 ;
  assign n2377 = n19386 & n2376 ;
  assign n19387 = ~n2372 ;
  assign n2378 = n19387 & n2377 ;
  assign n19388 = ~n2378 ;
  assign n2379 = n2371 & n19388 ;
  assign n2380 = x80 | n2379 ;
  assign n2381 = x80 & n2379 ;
  assign n2382 = n2180 & n19322 ;
  assign n2383 = n171 & n2382 ;
  assign n2384 = n2186 & n2383 ;
  assign n2385 = n2186 | n2383 ;
  assign n19389 = ~n2384 ;
  assign n2386 = n19389 & n2385 ;
  assign n19390 = ~n2381 ;
  assign n2387 = n19390 & n2386 ;
  assign n19391 = ~n2387 ;
  assign n2388 = n2380 & n19391 ;
  assign n2389 = x81 | n2388 ;
  assign n2390 = x81 & n2388 ;
  assign n2391 = n2189 & n19325 ;
  assign n2392 = n171 & n2391 ;
  assign n2393 = n2195 & n2392 ;
  assign n2394 = n2195 | n2392 ;
  assign n19392 = ~n2393 ;
  assign n2395 = n19392 & n2394 ;
  assign n19393 = ~n2390 ;
  assign n2396 = n19393 & n2395 ;
  assign n19394 = ~n2396 ;
  assign n2397 = n2389 & n19394 ;
  assign n2398 = x82 | n2397 ;
  assign n2399 = x82 & n2397 ;
  assign n2400 = n2198 & n19328 ;
  assign n2401 = n171 & n2400 ;
  assign n2402 = n2204 & n2401 ;
  assign n2403 = n2204 | n2401 ;
  assign n19395 = ~n2402 ;
  assign n2404 = n19395 & n2403 ;
  assign n19396 = ~n2399 ;
  assign n2405 = n19396 & n2404 ;
  assign n19397 = ~n2405 ;
  assign n2406 = n2398 & n19397 ;
  assign n2407 = x83 | n2406 ;
  assign n2408 = x83 & n2406 ;
  assign n2409 = n2207 & n19331 ;
  assign n2410 = n171 & n2409 ;
  assign n2411 = n2213 & n2410 ;
  assign n2412 = n2213 | n2410 ;
  assign n19398 = ~n2411 ;
  assign n2413 = n19398 & n2412 ;
  assign n19399 = ~n2408 ;
  assign n2414 = n19399 & n2413 ;
  assign n19400 = ~n2414 ;
  assign n2415 = n2407 & n19400 ;
  assign n2416 = x84 | n2415 ;
  assign n2417 = x84 & n2415 ;
  assign n2418 = n2216 & n19334 ;
  assign n2419 = n171 & n2418 ;
  assign n2420 = n2222 & n2419 ;
  assign n2421 = n2222 | n2419 ;
  assign n19401 = ~n2420 ;
  assign n2422 = n19401 & n2421 ;
  assign n19402 = ~n2417 ;
  assign n2423 = n19402 & n2422 ;
  assign n19403 = ~n2423 ;
  assign n2424 = n2416 & n19403 ;
  assign n2426 = x85 & n2424 ;
  assign n19404 = ~n2426 ;
  assign n2427 = n2241 & n19404 ;
  assign n2242 = n21884 | n2231 ;
  assign n2243 = n2234 & n2242 ;
  assign n19405 = ~x86 ;
  assign n2244 = n19405 & n2243 ;
  assign n2425 = x85 | n2424 ;
  assign n19406 = ~n2244 ;
  assign n2428 = n19406 & n2425 ;
  assign n19407 = ~n2427 ;
  assign n2429 = n19407 & n2428 ;
  assign n2430 = n18463 | n2429 ;
  assign n19408 = ~n2243 ;
  assign n2432 = x86 & n19408 ;
  assign n2433 = n2430 | n2432 ;
  assign n2434 = n2425 & n19404 ;
  assign n170 = ~n2433 ;
  assign n2435 = n170 & n2434 ;
  assign n19410 = ~n2241 ;
  assign n2436 = n19410 & n2435 ;
  assign n19411 = ~n2435 ;
  assign n2437 = n2241 & n19411 ;
  assign n2438 = n2436 | n2437 ;
  assign n19412 = ~x40 ;
  assign n2439 = n19412 & x64 ;
  assign n2441 = x65 | n2439 ;
  assign n2440 = x65 & n2439 ;
  assign n2442 = x64 & n170 ;
  assign n2443 = x41 & n2442 ;
  assign n2444 = x41 | n2442 ;
  assign n19413 = ~n2443 ;
  assign n2445 = n19413 & n2444 ;
  assign n19414 = ~n2440 ;
  assign n2446 = n19414 & n2445 ;
  assign n19415 = ~n2446 ;
  assign n2447 = n2441 & n19415 ;
  assign n2448 = x66 & n2447 ;
  assign n2449 = x66 | n2447 ;
  assign n2450 = n19344 & n2247 ;
  assign n2451 = n170 & n2450 ;
  assign n2452 = n2251 & n2451 ;
  assign n2453 = n2251 | n2451 ;
  assign n19416 = ~n2452 ;
  assign n2454 = n19416 & n2453 ;
  assign n19417 = ~n2454 ;
  assign n2455 = n2449 & n19417 ;
  assign n2456 = n2448 | n2455 ;
  assign n2457 = x67 & n2456 ;
  assign n2458 = x67 | n2456 ;
  assign n19418 = ~n2254 ;
  assign n2459 = n19418 & n2255 ;
  assign n2460 = n170 & n2459 ;
  assign n2461 = n2260 & n2460 ;
  assign n2462 = n2260 | n2460 ;
  assign n19419 = ~n2461 ;
  assign n2463 = n19419 & n2462 ;
  assign n19420 = ~n2463 ;
  assign n2464 = n2458 & n19420 ;
  assign n2465 = n2457 | n2464 ;
  assign n2466 = x68 & n2465 ;
  assign n2467 = x68 | n2465 ;
  assign n19421 = ~n2263 ;
  assign n2468 = n19421 & n2264 ;
  assign n2469 = n170 & n2468 ;
  assign n2470 = n19349 & n2469 ;
  assign n19422 = ~n2469 ;
  assign n2471 = n2269 & n19422 ;
  assign n2472 = n2470 | n2471 ;
  assign n19423 = ~n2472 ;
  assign n2473 = n2467 & n19423 ;
  assign n2474 = n2466 | n2473 ;
  assign n2475 = x69 & n2474 ;
  assign n2476 = x69 | n2474 ;
  assign n2477 = n19352 & n2273 ;
  assign n2478 = n170 & n2477 ;
  assign n19424 = ~n2278 ;
  assign n2479 = n19424 & n2478 ;
  assign n19425 = ~n2478 ;
  assign n2480 = n2278 & n19425 ;
  assign n2481 = n2479 | n2480 ;
  assign n19426 = ~n2481 ;
  assign n2482 = n2476 & n19426 ;
  assign n2483 = n2475 | n2482 ;
  assign n2484 = x70 & n2483 ;
  assign n2485 = x70 | n2483 ;
  assign n2486 = n2281 & n19356 ;
  assign n2487 = n170 & n2486 ;
  assign n19427 = ~n2287 ;
  assign n2488 = n19427 & n2487 ;
  assign n19428 = ~n2487 ;
  assign n2489 = n2287 & n19428 ;
  assign n2490 = n2488 | n2489 ;
  assign n19429 = ~n2490 ;
  assign n2491 = n2485 & n19429 ;
  assign n2492 = n2484 | n2491 ;
  assign n2493 = x71 & n2492 ;
  assign n2494 = x71 | n2492 ;
  assign n2495 = n2290 & n19360 ;
  assign n2496 = n170 & n2495 ;
  assign n19430 = ~n2296 ;
  assign n2497 = n19430 & n2496 ;
  assign n19431 = ~n2496 ;
  assign n2498 = n2296 & n19431 ;
  assign n2499 = n2497 | n2498 ;
  assign n19432 = ~n2499 ;
  assign n2500 = n2494 & n19432 ;
  assign n2501 = n2493 | n2500 ;
  assign n2502 = x72 & n2501 ;
  assign n2503 = x72 | n2501 ;
  assign n2504 = n2299 & n19363 ;
  assign n2505 = n170 & n2504 ;
  assign n2506 = n2305 & n2505 ;
  assign n2507 = n2305 | n2505 ;
  assign n19433 = ~n2506 ;
  assign n2508 = n19433 & n2507 ;
  assign n19434 = ~n2508 ;
  assign n2509 = n2503 & n19434 ;
  assign n2510 = n2502 | n2509 ;
  assign n2511 = x73 & n2510 ;
  assign n2512 = x73 | n2510 ;
  assign n2513 = n2308 & n19366 ;
  assign n2514 = n170 & n2513 ;
  assign n2515 = n2314 & n2514 ;
  assign n2516 = n2314 | n2514 ;
  assign n19435 = ~n2515 ;
  assign n2517 = n19435 & n2516 ;
  assign n19436 = ~n2517 ;
  assign n2518 = n2512 & n19436 ;
  assign n2519 = n2511 | n2518 ;
  assign n2520 = x74 & n2519 ;
  assign n2521 = x74 | n2519 ;
  assign n2522 = n2317 & n19369 ;
  assign n2523 = n170 & n2522 ;
  assign n2524 = n2323 & n2523 ;
  assign n2525 = n2323 | n2523 ;
  assign n19437 = ~n2524 ;
  assign n2526 = n19437 & n2525 ;
  assign n19438 = ~n2526 ;
  assign n2527 = n2521 & n19438 ;
  assign n2528 = n2520 | n2527 ;
  assign n2529 = x75 & n2528 ;
  assign n2530 = x75 | n2528 ;
  assign n2531 = n2326 & n19372 ;
  assign n2532 = n170 & n2531 ;
  assign n2533 = n2332 & n2532 ;
  assign n2534 = n2332 | n2532 ;
  assign n19439 = ~n2533 ;
  assign n2535 = n19439 & n2534 ;
  assign n19440 = ~n2535 ;
  assign n2536 = n2530 & n19440 ;
  assign n2537 = n2529 | n2536 ;
  assign n2538 = x76 & n2537 ;
  assign n2539 = x76 | n2537 ;
  assign n2540 = n2335 & n19375 ;
  assign n2541 = n170 & n2540 ;
  assign n2542 = n2341 & n2541 ;
  assign n2543 = n2341 | n2541 ;
  assign n19441 = ~n2542 ;
  assign n2544 = n19441 & n2543 ;
  assign n19442 = ~n2544 ;
  assign n2545 = n2539 & n19442 ;
  assign n2546 = n2538 | n2545 ;
  assign n2547 = x77 & n2546 ;
  assign n2548 = x77 | n2546 ;
  assign n2549 = n2344 & n19378 ;
  assign n2550 = n170 & n2549 ;
  assign n2551 = n2350 & n2550 ;
  assign n2552 = n2350 | n2550 ;
  assign n19443 = ~n2551 ;
  assign n2553 = n19443 & n2552 ;
  assign n19444 = ~n2553 ;
  assign n2554 = n2548 & n19444 ;
  assign n2555 = n2547 | n2554 ;
  assign n2556 = x78 & n2555 ;
  assign n2557 = x78 | n2555 ;
  assign n2558 = n2353 & n19381 ;
  assign n2559 = n170 & n2558 ;
  assign n2560 = n2359 & n2559 ;
  assign n2561 = n2359 | n2559 ;
  assign n19445 = ~n2560 ;
  assign n2562 = n19445 & n2561 ;
  assign n19446 = ~n2562 ;
  assign n2563 = n2557 & n19446 ;
  assign n2564 = n2556 | n2563 ;
  assign n2565 = x79 & n2564 ;
  assign n2566 = x79 | n2564 ;
  assign n2567 = n2362 & n19384 ;
  assign n2568 = n170 & n2567 ;
  assign n2569 = n2368 & n2568 ;
  assign n2570 = n2368 | n2568 ;
  assign n19447 = ~n2569 ;
  assign n2571 = n19447 & n2570 ;
  assign n19448 = ~n2571 ;
  assign n2572 = n2566 & n19448 ;
  assign n2573 = n2565 | n2572 ;
  assign n2574 = x80 & n2573 ;
  assign n2575 = x80 | n2573 ;
  assign n2576 = n2371 & n19387 ;
  assign n2577 = n170 & n2576 ;
  assign n2578 = n2377 & n2577 ;
  assign n2579 = n2377 | n2577 ;
  assign n19449 = ~n2578 ;
  assign n2580 = n19449 & n2579 ;
  assign n19450 = ~n2580 ;
  assign n2581 = n2575 & n19450 ;
  assign n2582 = n2574 | n2581 ;
  assign n2583 = x81 & n2582 ;
  assign n2584 = x81 | n2582 ;
  assign n2585 = n2380 & n19390 ;
  assign n2586 = n170 & n2585 ;
  assign n2587 = n2386 & n2586 ;
  assign n2588 = n2386 | n2586 ;
  assign n19451 = ~n2587 ;
  assign n2589 = n19451 & n2588 ;
  assign n19452 = ~n2589 ;
  assign n2590 = n2584 & n19452 ;
  assign n2591 = n2583 | n2590 ;
  assign n2592 = x82 & n2591 ;
  assign n2593 = x82 | n2591 ;
  assign n2594 = n2389 & n19393 ;
  assign n2595 = n170 & n2594 ;
  assign n2596 = n2395 & n2595 ;
  assign n2597 = n2395 | n2595 ;
  assign n19453 = ~n2596 ;
  assign n2598 = n19453 & n2597 ;
  assign n19454 = ~n2598 ;
  assign n2599 = n2593 & n19454 ;
  assign n2600 = n2592 | n2599 ;
  assign n2601 = x83 & n2600 ;
  assign n2602 = x83 | n2600 ;
  assign n2603 = n2398 & n19396 ;
  assign n2604 = n170 & n2603 ;
  assign n2605 = n2404 & n2604 ;
  assign n2606 = n2404 | n2604 ;
  assign n19455 = ~n2605 ;
  assign n2607 = n19455 & n2606 ;
  assign n19456 = ~n2607 ;
  assign n2608 = n2602 & n19456 ;
  assign n2609 = n2601 | n2608 ;
  assign n2610 = x84 & n2609 ;
  assign n2611 = x84 | n2609 ;
  assign n2612 = n2407 & n19399 ;
  assign n2613 = n170 & n2612 ;
  assign n2614 = n2413 & n2613 ;
  assign n2615 = n2413 | n2613 ;
  assign n19457 = ~n2614 ;
  assign n2616 = n19457 & n2615 ;
  assign n19458 = ~n2616 ;
  assign n2617 = n2611 & n19458 ;
  assign n2618 = n2610 | n2617 ;
  assign n2619 = x85 & n2618 ;
  assign n2620 = x85 | n2618 ;
  assign n2621 = n2416 & n19402 ;
  assign n2622 = n170 & n2621 ;
  assign n2623 = n2422 & n2622 ;
  assign n2624 = n2422 | n2622 ;
  assign n19459 = ~n2623 ;
  assign n2625 = n19459 & n2624 ;
  assign n19460 = ~n2625 ;
  assign n2626 = n2620 & n19460 ;
  assign n2627 = n2619 | n2626 ;
  assign n2628 = x86 & n2627 ;
  assign n2629 = x86 | n2627 ;
  assign n19461 = ~n2438 ;
  assign n2630 = n19461 & n2629 ;
  assign n2631 = n2628 | n2630 ;
  assign n2633 = x87 & n2631 ;
  assign n2634 = n18458 | n2633 ;
  assign n2632 = x87 | n2631 ;
  assign n2431 = n21884 | n2430 ;
  assign n2635 = n2243 & n2431 ;
  assign n19462 = ~n2635 ;
  assign n2636 = n2632 & n19462 ;
  assign n2637 = n2634 | n2636 ;
  assign n19463 = ~n2628 ;
  assign n2638 = n19463 & n2629 ;
  assign n169 = ~n2637 ;
  assign n2639 = n169 & n2638 ;
  assign n2640 = n19461 & n2639 ;
  assign n19465 = ~n2639 ;
  assign n2641 = n2438 & n19465 ;
  assign n2642 = n2640 | n2641 ;
  assign n19466 = ~x39 ;
  assign n2646 = n19466 & x64 ;
  assign n2648 = x65 | n2646 ;
  assign n2647 = x65 & n2646 ;
  assign n2649 = x64 & n169 ;
  assign n2650 = x40 & n2649 ;
  assign n2651 = x40 | n2649 ;
  assign n19467 = ~n2650 ;
  assign n2652 = n19467 & n2651 ;
  assign n19468 = ~n2647 ;
  assign n2653 = n19468 & n2652 ;
  assign n19469 = ~n2653 ;
  assign n2654 = n2648 & n19469 ;
  assign n2655 = x66 & n2654 ;
  assign n2656 = x66 | n2654 ;
  assign n2657 = n19414 & n2441 ;
  assign n2658 = n169 & n2657 ;
  assign n2659 = n2445 & n2658 ;
  assign n2660 = n2445 | n2658 ;
  assign n19470 = ~n2659 ;
  assign n2661 = n19470 & n2660 ;
  assign n19471 = ~n2661 ;
  assign n2662 = n2656 & n19471 ;
  assign n2663 = n2655 | n2662 ;
  assign n2664 = x67 & n2663 ;
  assign n2665 = x67 | n2663 ;
  assign n19472 = ~n2448 ;
  assign n2666 = n19472 & n2449 ;
  assign n2667 = n169 & n2666 ;
  assign n2668 = n2454 & n2667 ;
  assign n2669 = n2454 | n2667 ;
  assign n19473 = ~n2668 ;
  assign n2670 = n19473 & n2669 ;
  assign n19474 = ~n2670 ;
  assign n2671 = n2665 & n19474 ;
  assign n2672 = n2664 | n2671 ;
  assign n2673 = x68 & n2672 ;
  assign n2674 = x68 | n2672 ;
  assign n19475 = ~n2457 ;
  assign n2675 = n19475 & n2458 ;
  assign n2676 = n169 & n2675 ;
  assign n2677 = n2463 & n2676 ;
  assign n2678 = n2463 | n2676 ;
  assign n19476 = ~n2677 ;
  assign n2679 = n19476 & n2678 ;
  assign n19477 = ~n2679 ;
  assign n2680 = n2674 & n19477 ;
  assign n2681 = n2673 | n2680 ;
  assign n2682 = x69 & n2681 ;
  assign n2683 = x69 | n2681 ;
  assign n19478 = ~n2466 ;
  assign n2684 = n19478 & n2467 ;
  assign n2685 = n169 & n2684 ;
  assign n2686 = n19423 & n2685 ;
  assign n19479 = ~n2685 ;
  assign n2687 = n2472 & n19479 ;
  assign n2688 = n2686 | n2687 ;
  assign n19480 = ~n2688 ;
  assign n2689 = n2683 & n19480 ;
  assign n2690 = n2682 | n2689 ;
  assign n2691 = x70 & n2690 ;
  assign n2692 = x70 | n2690 ;
  assign n19481 = ~n2475 ;
  assign n2693 = n19481 & n2476 ;
  assign n2694 = n169 & n2693 ;
  assign n2695 = n19426 & n2694 ;
  assign n19482 = ~n2694 ;
  assign n2696 = n2481 & n19482 ;
  assign n2697 = n2695 | n2696 ;
  assign n19483 = ~n2697 ;
  assign n2698 = n2692 & n19483 ;
  assign n2699 = n2691 | n2698 ;
  assign n2700 = x71 & n2699 ;
  assign n2701 = x71 | n2699 ;
  assign n19484 = ~n2484 ;
  assign n2702 = n19484 & n2485 ;
  assign n2703 = n169 & n2702 ;
  assign n2704 = n2490 & n2703 ;
  assign n2705 = n2490 | n2703 ;
  assign n19485 = ~n2704 ;
  assign n2706 = n19485 & n2705 ;
  assign n19486 = ~n2706 ;
  assign n2707 = n2701 & n19486 ;
  assign n2708 = n2700 | n2707 ;
  assign n2709 = x72 & n2708 ;
  assign n2710 = x72 | n2708 ;
  assign n19487 = ~n2493 ;
  assign n2711 = n19487 & n2494 ;
  assign n2712 = n169 & n2711 ;
  assign n2713 = n2499 & n2712 ;
  assign n2714 = n2499 | n2712 ;
  assign n19488 = ~n2713 ;
  assign n2715 = n19488 & n2714 ;
  assign n19489 = ~n2715 ;
  assign n2716 = n2710 & n19489 ;
  assign n2717 = n2709 | n2716 ;
  assign n2718 = x73 & n2717 ;
  assign n2719 = x73 | n2717 ;
  assign n19490 = ~n2502 ;
  assign n2720 = n19490 & n2503 ;
  assign n2721 = n169 & n2720 ;
  assign n2722 = n2508 & n2721 ;
  assign n2723 = n2508 | n2721 ;
  assign n19491 = ~n2722 ;
  assign n2724 = n19491 & n2723 ;
  assign n19492 = ~n2724 ;
  assign n2725 = n2719 & n19492 ;
  assign n2726 = n2718 | n2725 ;
  assign n2727 = x74 & n2726 ;
  assign n2728 = x74 | n2726 ;
  assign n19493 = ~n2511 ;
  assign n2729 = n19493 & n2512 ;
  assign n2730 = n169 & n2729 ;
  assign n2731 = n2517 & n2730 ;
  assign n2732 = n2517 | n2730 ;
  assign n19494 = ~n2731 ;
  assign n2733 = n19494 & n2732 ;
  assign n19495 = ~n2733 ;
  assign n2734 = n2728 & n19495 ;
  assign n2735 = n2727 | n2734 ;
  assign n2736 = x75 & n2735 ;
  assign n2737 = x75 | n2735 ;
  assign n19496 = ~n2520 ;
  assign n2738 = n19496 & n2521 ;
  assign n2739 = n169 & n2738 ;
  assign n2740 = n2526 & n2739 ;
  assign n2741 = n2526 | n2739 ;
  assign n19497 = ~n2740 ;
  assign n2742 = n19497 & n2741 ;
  assign n19498 = ~n2742 ;
  assign n2743 = n2737 & n19498 ;
  assign n2744 = n2736 | n2743 ;
  assign n2745 = x76 & n2744 ;
  assign n2746 = x76 | n2744 ;
  assign n19499 = ~n2529 ;
  assign n2747 = n19499 & n2530 ;
  assign n2748 = n169 & n2747 ;
  assign n2749 = n2535 & n2748 ;
  assign n2750 = n2535 | n2748 ;
  assign n19500 = ~n2749 ;
  assign n2751 = n19500 & n2750 ;
  assign n19501 = ~n2751 ;
  assign n2752 = n2746 & n19501 ;
  assign n2753 = n2745 | n2752 ;
  assign n2754 = x77 & n2753 ;
  assign n2755 = x77 | n2753 ;
  assign n19502 = ~n2538 ;
  assign n2756 = n19502 & n2539 ;
  assign n2757 = n169 & n2756 ;
  assign n2758 = n2544 & n2757 ;
  assign n2759 = n2544 | n2757 ;
  assign n19503 = ~n2758 ;
  assign n2760 = n19503 & n2759 ;
  assign n19504 = ~n2760 ;
  assign n2761 = n2755 & n19504 ;
  assign n2762 = n2754 | n2761 ;
  assign n2763 = x78 & n2762 ;
  assign n2764 = x78 | n2762 ;
  assign n19505 = ~n2547 ;
  assign n2765 = n19505 & n2548 ;
  assign n2766 = n169 & n2765 ;
  assign n2767 = n2553 & n2766 ;
  assign n2768 = n2553 | n2766 ;
  assign n19506 = ~n2767 ;
  assign n2769 = n19506 & n2768 ;
  assign n19507 = ~n2769 ;
  assign n2770 = n2764 & n19507 ;
  assign n2771 = n2763 | n2770 ;
  assign n2772 = x79 & n2771 ;
  assign n2773 = x79 | n2771 ;
  assign n19508 = ~n2556 ;
  assign n2774 = n19508 & n2557 ;
  assign n2775 = n169 & n2774 ;
  assign n2776 = n2562 & n2775 ;
  assign n2777 = n2562 | n2775 ;
  assign n19509 = ~n2776 ;
  assign n2778 = n19509 & n2777 ;
  assign n19510 = ~n2778 ;
  assign n2779 = n2773 & n19510 ;
  assign n2780 = n2772 | n2779 ;
  assign n2781 = x80 & n2780 ;
  assign n2782 = x80 | n2780 ;
  assign n19511 = ~n2565 ;
  assign n2783 = n19511 & n2566 ;
  assign n2784 = n169 & n2783 ;
  assign n2785 = n2571 & n2784 ;
  assign n2786 = n2571 | n2784 ;
  assign n19512 = ~n2785 ;
  assign n2787 = n19512 & n2786 ;
  assign n19513 = ~n2787 ;
  assign n2788 = n2782 & n19513 ;
  assign n2789 = n2781 | n2788 ;
  assign n2790 = x81 & n2789 ;
  assign n2791 = x81 | n2789 ;
  assign n19514 = ~n2574 ;
  assign n2792 = n19514 & n2575 ;
  assign n2793 = n169 & n2792 ;
  assign n2794 = n2580 & n2793 ;
  assign n2795 = n2580 | n2793 ;
  assign n19515 = ~n2794 ;
  assign n2796 = n19515 & n2795 ;
  assign n19516 = ~n2796 ;
  assign n2797 = n2791 & n19516 ;
  assign n2798 = n2790 | n2797 ;
  assign n2799 = x82 & n2798 ;
  assign n2800 = x82 | n2798 ;
  assign n19517 = ~n2583 ;
  assign n2801 = n19517 & n2584 ;
  assign n2802 = n169 & n2801 ;
  assign n2803 = n2589 & n2802 ;
  assign n2804 = n2589 | n2802 ;
  assign n19518 = ~n2803 ;
  assign n2805 = n19518 & n2804 ;
  assign n19519 = ~n2805 ;
  assign n2806 = n2800 & n19519 ;
  assign n2807 = n2799 | n2806 ;
  assign n2808 = x83 & n2807 ;
  assign n2809 = x83 | n2807 ;
  assign n19520 = ~n2592 ;
  assign n2810 = n19520 & n2593 ;
  assign n2811 = n169 & n2810 ;
  assign n2812 = n2598 & n2811 ;
  assign n2813 = n2598 | n2811 ;
  assign n19521 = ~n2812 ;
  assign n2814 = n19521 & n2813 ;
  assign n19522 = ~n2814 ;
  assign n2815 = n2809 & n19522 ;
  assign n2816 = n2808 | n2815 ;
  assign n2817 = x84 & n2816 ;
  assign n2818 = x84 | n2816 ;
  assign n19523 = ~n2601 ;
  assign n2819 = n19523 & n2602 ;
  assign n2820 = n169 & n2819 ;
  assign n2821 = n2607 & n2820 ;
  assign n2822 = n2607 | n2820 ;
  assign n19524 = ~n2821 ;
  assign n2823 = n19524 & n2822 ;
  assign n19525 = ~n2823 ;
  assign n2824 = n2818 & n19525 ;
  assign n2825 = n2817 | n2824 ;
  assign n2826 = x85 & n2825 ;
  assign n2827 = x85 | n2825 ;
  assign n19526 = ~n2610 ;
  assign n2828 = n19526 & n2611 ;
  assign n2829 = n169 & n2828 ;
  assign n2830 = n2616 & n2829 ;
  assign n2831 = n2616 | n2829 ;
  assign n19527 = ~n2830 ;
  assign n2832 = n19527 & n2831 ;
  assign n19528 = ~n2832 ;
  assign n2833 = n2827 & n19528 ;
  assign n2834 = n2826 | n2833 ;
  assign n2835 = x86 & n2834 ;
  assign n2836 = x86 | n2834 ;
  assign n19529 = ~n2619 ;
  assign n2837 = n19529 & n2620 ;
  assign n2838 = n169 & n2837 ;
  assign n2839 = n2625 & n2838 ;
  assign n2840 = n2625 | n2838 ;
  assign n19530 = ~n2839 ;
  assign n2841 = n19530 & n2840 ;
  assign n19531 = ~n2841 ;
  assign n2842 = n2836 & n19531 ;
  assign n2843 = n2835 | n2842 ;
  assign n2845 = x87 & n2843 ;
  assign n19532 = ~n2845 ;
  assign n2846 = n2642 & n19532 ;
  assign n2643 = n21884 | n2634 ;
  assign n2644 = n2635 & n2643 ;
  assign n19533 = ~x88 ;
  assign n2645 = n19533 & n2644 ;
  assign n2844 = x87 | n2843 ;
  assign n19534 = ~n2645 ;
  assign n2847 = n19534 & n2844 ;
  assign n19535 = ~n2846 ;
  assign n2848 = n19535 & n2847 ;
  assign n2849 = n18453 | n2848 ;
  assign n19536 = ~n2644 ;
  assign n2851 = x88 & n19536 ;
  assign n2852 = n2849 | n2851 ;
  assign n2853 = n2844 & n19532 ;
  assign n168 = ~n2852 ;
  assign n2854 = n168 & n2853 ;
  assign n2855 = n2642 & n2854 ;
  assign n2856 = n2642 | n2854 ;
  assign n19538 = ~n2855 ;
  assign n2857 = n19538 & n2856 ;
  assign n19539 = ~x38 ;
  assign n2858 = n19539 & x64 ;
  assign n2860 = x65 | n2858 ;
  assign n2859 = x65 & n2858 ;
  assign n2861 = x64 & n168 ;
  assign n2862 = x39 & n2861 ;
  assign n2863 = x39 | n2861 ;
  assign n19540 = ~n2862 ;
  assign n2864 = n19540 & n2863 ;
  assign n19541 = ~n2859 ;
  assign n2865 = n19541 & n2864 ;
  assign n19542 = ~n2865 ;
  assign n2866 = n2860 & n19542 ;
  assign n2867 = x66 & n2866 ;
  assign n2868 = x66 | n2866 ;
  assign n2869 = n19468 & n2648 ;
  assign n2870 = n168 & n2869 ;
  assign n2871 = n2652 & n2870 ;
  assign n2872 = n2652 | n2870 ;
  assign n19543 = ~n2871 ;
  assign n2873 = n19543 & n2872 ;
  assign n19544 = ~n2873 ;
  assign n2874 = n2868 & n19544 ;
  assign n2875 = n2867 | n2874 ;
  assign n2876 = x67 & n2875 ;
  assign n2877 = x67 | n2875 ;
  assign n19545 = ~n2655 ;
  assign n2878 = n19545 & n2656 ;
  assign n2879 = n168 & n2878 ;
  assign n2880 = n2661 & n2879 ;
  assign n2881 = n2661 | n2879 ;
  assign n19546 = ~n2880 ;
  assign n2882 = n19546 & n2881 ;
  assign n19547 = ~n2882 ;
  assign n2883 = n2877 & n19547 ;
  assign n2884 = n2876 | n2883 ;
  assign n2885 = x68 & n2884 ;
  assign n2886 = x68 | n2884 ;
  assign n19548 = ~n2664 ;
  assign n2887 = n19548 & n2665 ;
  assign n2888 = n168 & n2887 ;
  assign n2889 = n2670 & n2888 ;
  assign n2890 = n2670 | n2888 ;
  assign n19549 = ~n2889 ;
  assign n2891 = n19549 & n2890 ;
  assign n19550 = ~n2891 ;
  assign n2892 = n2886 & n19550 ;
  assign n2893 = n2885 | n2892 ;
  assign n2894 = x69 & n2893 ;
  assign n2895 = x69 | n2893 ;
  assign n19551 = ~n2673 ;
  assign n2896 = n19551 & n2674 ;
  assign n2897 = n168 & n2896 ;
  assign n2898 = n19477 & n2897 ;
  assign n19552 = ~n2897 ;
  assign n2899 = n2679 & n19552 ;
  assign n2900 = n2898 | n2899 ;
  assign n19553 = ~n2900 ;
  assign n2901 = n2895 & n19553 ;
  assign n2902 = n2894 | n2901 ;
  assign n2903 = x70 & n2902 ;
  assign n2904 = x70 | n2902 ;
  assign n19554 = ~n2682 ;
  assign n2905 = n19554 & n2683 ;
  assign n2906 = n168 & n2905 ;
  assign n2907 = n19480 & n2906 ;
  assign n19555 = ~n2906 ;
  assign n2908 = n2688 & n19555 ;
  assign n2909 = n2907 | n2908 ;
  assign n19556 = ~n2909 ;
  assign n2910 = n2904 & n19556 ;
  assign n2911 = n2903 | n2910 ;
  assign n2912 = x71 & n2911 ;
  assign n2913 = x71 | n2911 ;
  assign n19557 = ~n2691 ;
  assign n2914 = n19557 & n2692 ;
  assign n2915 = n168 & n2914 ;
  assign n2916 = n2697 & n2915 ;
  assign n2917 = n2697 | n2915 ;
  assign n19558 = ~n2916 ;
  assign n2918 = n19558 & n2917 ;
  assign n19559 = ~n2918 ;
  assign n2919 = n2913 & n19559 ;
  assign n2920 = n2912 | n2919 ;
  assign n2921 = x72 & n2920 ;
  assign n2922 = x72 | n2920 ;
  assign n19560 = ~n2700 ;
  assign n2923 = n19560 & n2701 ;
  assign n2924 = n168 & n2923 ;
  assign n2925 = n2706 & n2924 ;
  assign n2926 = n2706 | n2924 ;
  assign n19561 = ~n2925 ;
  assign n2927 = n19561 & n2926 ;
  assign n19562 = ~n2927 ;
  assign n2928 = n2922 & n19562 ;
  assign n2929 = n2921 | n2928 ;
  assign n2930 = x73 & n2929 ;
  assign n2931 = x73 | n2929 ;
  assign n19563 = ~n2709 ;
  assign n2932 = n19563 & n2710 ;
  assign n2933 = n168 & n2932 ;
  assign n2934 = n2715 & n2933 ;
  assign n2935 = n2715 | n2933 ;
  assign n19564 = ~n2934 ;
  assign n2936 = n19564 & n2935 ;
  assign n19565 = ~n2936 ;
  assign n2937 = n2931 & n19565 ;
  assign n2938 = n2930 | n2937 ;
  assign n2939 = x74 & n2938 ;
  assign n2940 = x74 | n2938 ;
  assign n19566 = ~n2718 ;
  assign n2941 = n19566 & n2719 ;
  assign n2942 = n168 & n2941 ;
  assign n2943 = n19492 & n2942 ;
  assign n19567 = ~n2942 ;
  assign n2944 = n2724 & n19567 ;
  assign n2945 = n2943 | n2944 ;
  assign n19568 = ~n2945 ;
  assign n2946 = n2940 & n19568 ;
  assign n2947 = n2939 | n2946 ;
  assign n2948 = x75 & n2947 ;
  assign n2949 = x75 | n2947 ;
  assign n19569 = ~n2727 ;
  assign n2950 = n19569 & n2728 ;
  assign n2951 = n168 & n2950 ;
  assign n2952 = n19495 & n2951 ;
  assign n19570 = ~n2951 ;
  assign n2953 = n2733 & n19570 ;
  assign n2954 = n2952 | n2953 ;
  assign n19571 = ~n2954 ;
  assign n2955 = n2949 & n19571 ;
  assign n2956 = n2948 | n2955 ;
  assign n2957 = x76 & n2956 ;
  assign n2958 = x76 | n2956 ;
  assign n19572 = ~n2736 ;
  assign n2959 = n19572 & n2737 ;
  assign n2960 = n168 & n2959 ;
  assign n2961 = n19498 & n2960 ;
  assign n19573 = ~n2960 ;
  assign n2962 = n2742 & n19573 ;
  assign n2963 = n2961 | n2962 ;
  assign n19574 = ~n2963 ;
  assign n2964 = n2958 & n19574 ;
  assign n2965 = n2957 | n2964 ;
  assign n2966 = x77 & n2965 ;
  assign n2967 = x77 | n2965 ;
  assign n19575 = ~n2745 ;
  assign n2968 = n19575 & n2746 ;
  assign n2969 = n168 & n2968 ;
  assign n2970 = n19501 & n2969 ;
  assign n19576 = ~n2969 ;
  assign n2971 = n2751 & n19576 ;
  assign n2972 = n2970 | n2971 ;
  assign n19577 = ~n2972 ;
  assign n2973 = n2967 & n19577 ;
  assign n2974 = n2966 | n2973 ;
  assign n2975 = x78 & n2974 ;
  assign n2976 = x78 | n2974 ;
  assign n19578 = ~n2754 ;
  assign n2977 = n19578 & n2755 ;
  assign n2978 = n168 & n2977 ;
  assign n2979 = n19504 & n2978 ;
  assign n19579 = ~n2978 ;
  assign n2980 = n2760 & n19579 ;
  assign n2981 = n2979 | n2980 ;
  assign n19580 = ~n2981 ;
  assign n2982 = n2976 & n19580 ;
  assign n2983 = n2975 | n2982 ;
  assign n2984 = x79 & n2983 ;
  assign n2985 = x79 | n2983 ;
  assign n19581 = ~n2763 ;
  assign n2986 = n19581 & n2764 ;
  assign n2987 = n168 & n2986 ;
  assign n2988 = n19507 & n2987 ;
  assign n19582 = ~n2987 ;
  assign n2989 = n2769 & n19582 ;
  assign n2990 = n2988 | n2989 ;
  assign n19583 = ~n2990 ;
  assign n2991 = n2985 & n19583 ;
  assign n2992 = n2984 | n2991 ;
  assign n2993 = x80 & n2992 ;
  assign n2994 = x80 | n2992 ;
  assign n19584 = ~n2772 ;
  assign n2995 = n19584 & n2773 ;
  assign n2996 = n168 & n2995 ;
  assign n2997 = n19510 & n2996 ;
  assign n19585 = ~n2996 ;
  assign n2998 = n2778 & n19585 ;
  assign n2999 = n2997 | n2998 ;
  assign n19586 = ~n2999 ;
  assign n3000 = n2994 & n19586 ;
  assign n3001 = n2993 | n3000 ;
  assign n3002 = x81 & n3001 ;
  assign n3003 = x81 | n3001 ;
  assign n19587 = ~n2781 ;
  assign n3004 = n19587 & n2782 ;
  assign n3005 = n168 & n3004 ;
  assign n3006 = n19513 & n3005 ;
  assign n19588 = ~n3005 ;
  assign n3007 = n2787 & n19588 ;
  assign n3008 = n3006 | n3007 ;
  assign n19589 = ~n3008 ;
  assign n3009 = n3003 & n19589 ;
  assign n3010 = n3002 | n3009 ;
  assign n3011 = x82 & n3010 ;
  assign n3012 = x82 | n3010 ;
  assign n19590 = ~n2790 ;
  assign n3013 = n19590 & n2791 ;
  assign n3014 = n168 & n3013 ;
  assign n3015 = n19516 & n3014 ;
  assign n19591 = ~n3014 ;
  assign n3016 = n2796 & n19591 ;
  assign n3017 = n3015 | n3016 ;
  assign n19592 = ~n3017 ;
  assign n3018 = n3012 & n19592 ;
  assign n3019 = n3011 | n3018 ;
  assign n3020 = x83 & n3019 ;
  assign n3021 = x83 | n3019 ;
  assign n19593 = ~n2799 ;
  assign n3022 = n19593 & n2800 ;
  assign n3023 = n168 & n3022 ;
  assign n3024 = n19519 & n3023 ;
  assign n19594 = ~n3023 ;
  assign n3025 = n2805 & n19594 ;
  assign n3026 = n3024 | n3025 ;
  assign n19595 = ~n3026 ;
  assign n3027 = n3021 & n19595 ;
  assign n3028 = n3020 | n3027 ;
  assign n3029 = x84 & n3028 ;
  assign n3030 = x84 | n3028 ;
  assign n19596 = ~n2808 ;
  assign n3031 = n19596 & n2809 ;
  assign n3032 = n168 & n3031 ;
  assign n3033 = n19522 & n3032 ;
  assign n19597 = ~n3032 ;
  assign n3034 = n2814 & n19597 ;
  assign n3035 = n3033 | n3034 ;
  assign n19598 = ~n3035 ;
  assign n3036 = n3030 & n19598 ;
  assign n3037 = n3029 | n3036 ;
  assign n3038 = x85 & n3037 ;
  assign n3039 = x85 | n3037 ;
  assign n19599 = ~n2817 ;
  assign n3040 = n19599 & n2818 ;
  assign n3041 = n168 & n3040 ;
  assign n3042 = n19525 & n3041 ;
  assign n19600 = ~n3041 ;
  assign n3043 = n2823 & n19600 ;
  assign n3044 = n3042 | n3043 ;
  assign n19601 = ~n3044 ;
  assign n3045 = n3039 & n19601 ;
  assign n3046 = n3038 | n3045 ;
  assign n3047 = x86 & n3046 ;
  assign n3048 = x86 | n3046 ;
  assign n19602 = ~n2826 ;
  assign n3049 = n19602 & n2827 ;
  assign n3050 = n168 & n3049 ;
  assign n3051 = n19528 & n3050 ;
  assign n19603 = ~n3050 ;
  assign n3052 = n2832 & n19603 ;
  assign n3053 = n3051 | n3052 ;
  assign n19604 = ~n3053 ;
  assign n3054 = n3048 & n19604 ;
  assign n3055 = n3047 | n3054 ;
  assign n3056 = x87 & n3055 ;
  assign n3057 = x87 | n3055 ;
  assign n19605 = ~n2835 ;
  assign n3058 = n19605 & n2836 ;
  assign n3059 = n168 & n3058 ;
  assign n3060 = n19531 & n3059 ;
  assign n19606 = ~n3059 ;
  assign n3061 = n2841 & n19606 ;
  assign n3062 = n3060 | n3061 ;
  assign n19607 = ~n3062 ;
  assign n3063 = n3057 & n19607 ;
  assign n3064 = n3056 | n3063 ;
  assign n3065 = x88 & n3064 ;
  assign n19608 = ~n3065 ;
  assign n3066 = n2857 & n19608 ;
  assign n3070 = x88 | n3064 ;
  assign n2850 = n21884 | n2849 ;
  assign n3067 = n2644 & n2850 ;
  assign n19609 = ~x89 ;
  assign n3071 = n19609 & n3067 ;
  assign n19610 = ~n3071 ;
  assign n3072 = n3070 & n19610 ;
  assign n19611 = ~n3066 ;
  assign n3074 = n19611 & n3072 ;
  assign n19612 = ~n18448 ;
  assign n3073 = n19612 & n3067 ;
  assign n19613 = ~n3073 ;
  assign n3075 = n18453 & n19613 ;
  assign n3076 = n3074 | n3075 ;
  assign n3077 = n19608 & n3070 ;
  assign n167 = ~n3076 ;
  assign n3078 = n167 & n3077 ;
  assign n3079 = n2857 & n3078 ;
  assign n3080 = n2857 | n3078 ;
  assign n19615 = ~n3079 ;
  assign n3081 = n19615 & n3080 ;
  assign n19616 = ~x37 ;
  assign n3082 = n19616 & x64 ;
  assign n3084 = x65 | n3082 ;
  assign n3083 = x65 & n3082 ;
  assign n3085 = x64 & n167 ;
  assign n3086 = x38 & n3085 ;
  assign n3087 = x38 | n3085 ;
  assign n19617 = ~n3086 ;
  assign n3088 = n19617 & n3087 ;
  assign n19618 = ~n3083 ;
  assign n3089 = n19618 & n3088 ;
  assign n19619 = ~n3089 ;
  assign n3090 = n3084 & n19619 ;
  assign n3091 = x66 & n3090 ;
  assign n3092 = x66 | n3090 ;
  assign n3093 = n19541 & n2860 ;
  assign n3094 = n167 & n3093 ;
  assign n3095 = n2864 & n3094 ;
  assign n3096 = n2864 | n3094 ;
  assign n19620 = ~n3095 ;
  assign n3097 = n19620 & n3096 ;
  assign n19621 = ~n3097 ;
  assign n3098 = n3092 & n19621 ;
  assign n3099 = n3091 | n3098 ;
  assign n3100 = x67 & n3099 ;
  assign n3101 = x67 | n3099 ;
  assign n19622 = ~n2867 ;
  assign n3102 = n19622 & n2868 ;
  assign n3103 = n167 & n3102 ;
  assign n3104 = n2873 & n3103 ;
  assign n3105 = n2873 | n3103 ;
  assign n19623 = ~n3104 ;
  assign n3106 = n19623 & n3105 ;
  assign n19624 = ~n3106 ;
  assign n3107 = n3101 & n19624 ;
  assign n3108 = n3100 | n3107 ;
  assign n3110 = x68 | n3108 ;
  assign n3109 = x68 & n3108 ;
  assign n19625 = ~n2876 ;
  assign n3111 = n19625 & n2877 ;
  assign n3112 = n167 & n3111 ;
  assign n3113 = n2882 & n3112 ;
  assign n3114 = n2882 | n3112 ;
  assign n19626 = ~n3113 ;
  assign n3115 = n19626 & n3114 ;
  assign n19627 = ~n3109 ;
  assign n3116 = n19627 & n3115 ;
  assign n19628 = ~n3116 ;
  assign n3117 = n3110 & n19628 ;
  assign n3118 = x69 | n3117 ;
  assign n3119 = x69 & n3117 ;
  assign n19629 = ~n2885 ;
  assign n3120 = n19629 & n2886 ;
  assign n3121 = n167 & n3120 ;
  assign n3122 = n2891 & n3121 ;
  assign n3123 = n2891 | n3121 ;
  assign n19630 = ~n3122 ;
  assign n3124 = n19630 & n3123 ;
  assign n19631 = ~n3119 ;
  assign n3125 = n19631 & n3124 ;
  assign n19632 = ~n3125 ;
  assign n3126 = n3118 & n19632 ;
  assign n3127 = x70 | n3126 ;
  assign n3128 = x70 & n3126 ;
  assign n19633 = ~n2894 ;
  assign n3129 = n19633 & n2895 ;
  assign n3130 = n167 & n3129 ;
  assign n3131 = n2900 & n3130 ;
  assign n3132 = n2900 | n3130 ;
  assign n19634 = ~n3131 ;
  assign n3133 = n19634 & n3132 ;
  assign n19635 = ~n3128 ;
  assign n3134 = n19635 & n3133 ;
  assign n19636 = ~n3134 ;
  assign n3135 = n3127 & n19636 ;
  assign n3136 = x71 | n3135 ;
  assign n3137 = x71 & n3135 ;
  assign n19637 = ~n2903 ;
  assign n3138 = n19637 & n2904 ;
  assign n3139 = n167 & n3138 ;
  assign n3140 = n2909 & n3139 ;
  assign n3141 = n2909 | n3139 ;
  assign n19638 = ~n3140 ;
  assign n3142 = n19638 & n3141 ;
  assign n19639 = ~n3137 ;
  assign n3143 = n19639 & n3142 ;
  assign n19640 = ~n3143 ;
  assign n3144 = n3136 & n19640 ;
  assign n3146 = x72 & n3144 ;
  assign n3145 = x72 | n3144 ;
  assign n19641 = ~n2912 ;
  assign n3147 = n19641 & n2913 ;
  assign n3148 = n167 & n3147 ;
  assign n3149 = n2918 & n3148 ;
  assign n3150 = n2918 | n3148 ;
  assign n19642 = ~n3149 ;
  assign n3151 = n19642 & n3150 ;
  assign n19643 = ~n3151 ;
  assign n3152 = n3145 & n19643 ;
  assign n3153 = n3146 | n3152 ;
  assign n3154 = x73 & n3153 ;
  assign n3155 = x73 | n3153 ;
  assign n19644 = ~n2921 ;
  assign n3156 = n19644 & n2922 ;
  assign n3157 = n167 & n3156 ;
  assign n3158 = n2927 & n3157 ;
  assign n3159 = n2927 | n3157 ;
  assign n19645 = ~n3158 ;
  assign n3160 = n19645 & n3159 ;
  assign n19646 = ~n3160 ;
  assign n3161 = n3155 & n19646 ;
  assign n3162 = n3154 | n3161 ;
  assign n3163 = x74 & n3162 ;
  assign n3164 = x74 | n3162 ;
  assign n19647 = ~n2930 ;
  assign n3165 = n19647 & n2931 ;
  assign n3166 = n167 & n3165 ;
  assign n3167 = n2936 & n3166 ;
  assign n3168 = n2936 | n3166 ;
  assign n19648 = ~n3167 ;
  assign n3169 = n19648 & n3168 ;
  assign n19649 = ~n3169 ;
  assign n3170 = n3164 & n19649 ;
  assign n3171 = n3163 | n3170 ;
  assign n3172 = x75 & n3171 ;
  assign n3173 = x75 | n3171 ;
  assign n19650 = ~n2939 ;
  assign n3174 = n19650 & n2940 ;
  assign n3175 = n167 & n3174 ;
  assign n3176 = n19568 & n3175 ;
  assign n19651 = ~n3175 ;
  assign n3177 = n2945 & n19651 ;
  assign n3178 = n3176 | n3177 ;
  assign n19652 = ~n3178 ;
  assign n3179 = n3173 & n19652 ;
  assign n3180 = n3172 | n3179 ;
  assign n3181 = x76 & n3180 ;
  assign n3182 = x76 | n3180 ;
  assign n19653 = ~n2948 ;
  assign n3183 = n19653 & n2949 ;
  assign n3184 = n167 & n3183 ;
  assign n3185 = n19571 & n3184 ;
  assign n19654 = ~n3184 ;
  assign n3186 = n2954 & n19654 ;
  assign n3187 = n3185 | n3186 ;
  assign n19655 = ~n3187 ;
  assign n3188 = n3182 & n19655 ;
  assign n3189 = n3181 | n3188 ;
  assign n3190 = x77 & n3189 ;
  assign n3191 = x77 | n3189 ;
  assign n19656 = ~n2957 ;
  assign n3192 = n19656 & n2958 ;
  assign n3193 = n167 & n3192 ;
  assign n3194 = n19574 & n3193 ;
  assign n19657 = ~n3193 ;
  assign n3195 = n2963 & n19657 ;
  assign n3196 = n3194 | n3195 ;
  assign n19658 = ~n3196 ;
  assign n3197 = n3191 & n19658 ;
  assign n3198 = n3190 | n3197 ;
  assign n3199 = x78 & n3198 ;
  assign n3200 = x78 | n3198 ;
  assign n19659 = ~n2966 ;
  assign n3201 = n19659 & n2967 ;
  assign n3202 = n167 & n3201 ;
  assign n3203 = n19577 & n3202 ;
  assign n19660 = ~n3202 ;
  assign n3204 = n2972 & n19660 ;
  assign n3205 = n3203 | n3204 ;
  assign n19661 = ~n3205 ;
  assign n3206 = n3200 & n19661 ;
  assign n3207 = n3199 | n3206 ;
  assign n3208 = x79 & n3207 ;
  assign n3209 = x79 | n3207 ;
  assign n19662 = ~n2975 ;
  assign n3210 = n19662 & n2976 ;
  assign n3211 = n167 & n3210 ;
  assign n3212 = n19580 & n3211 ;
  assign n19663 = ~n3211 ;
  assign n3213 = n2981 & n19663 ;
  assign n3214 = n3212 | n3213 ;
  assign n19664 = ~n3214 ;
  assign n3215 = n3209 & n19664 ;
  assign n3216 = n3208 | n3215 ;
  assign n3217 = x80 & n3216 ;
  assign n3218 = x80 | n3216 ;
  assign n19665 = ~n2984 ;
  assign n3219 = n19665 & n2985 ;
  assign n3220 = n167 & n3219 ;
  assign n3221 = n19583 & n3220 ;
  assign n19666 = ~n3220 ;
  assign n3222 = n2990 & n19666 ;
  assign n3223 = n3221 | n3222 ;
  assign n19667 = ~n3223 ;
  assign n3224 = n3218 & n19667 ;
  assign n3225 = n3217 | n3224 ;
  assign n3226 = x81 & n3225 ;
  assign n3227 = x81 | n3225 ;
  assign n19668 = ~n2993 ;
  assign n3228 = n19668 & n2994 ;
  assign n3229 = n167 & n3228 ;
  assign n3230 = n19586 & n3229 ;
  assign n19669 = ~n3229 ;
  assign n3231 = n2999 & n19669 ;
  assign n3232 = n3230 | n3231 ;
  assign n19670 = ~n3232 ;
  assign n3233 = n3227 & n19670 ;
  assign n3234 = n3226 | n3233 ;
  assign n3235 = x82 & n3234 ;
  assign n3236 = x82 | n3234 ;
  assign n19671 = ~n3002 ;
  assign n3237 = n19671 & n3003 ;
  assign n3238 = n167 & n3237 ;
  assign n3239 = n19589 & n3238 ;
  assign n19672 = ~n3238 ;
  assign n3240 = n3008 & n19672 ;
  assign n3241 = n3239 | n3240 ;
  assign n19673 = ~n3241 ;
  assign n3242 = n3236 & n19673 ;
  assign n3243 = n3235 | n3242 ;
  assign n3244 = x83 & n3243 ;
  assign n3245 = x83 | n3243 ;
  assign n19674 = ~n3011 ;
  assign n3246 = n19674 & n3012 ;
  assign n3247 = n167 & n3246 ;
  assign n3248 = n19592 & n3247 ;
  assign n19675 = ~n3247 ;
  assign n3249 = n3017 & n19675 ;
  assign n3250 = n3248 | n3249 ;
  assign n19676 = ~n3250 ;
  assign n3251 = n3245 & n19676 ;
  assign n3252 = n3244 | n3251 ;
  assign n3253 = x84 & n3252 ;
  assign n3254 = x84 | n3252 ;
  assign n19677 = ~n3020 ;
  assign n3255 = n19677 & n3021 ;
  assign n3256 = n167 & n3255 ;
  assign n3257 = n19595 & n3256 ;
  assign n19678 = ~n3256 ;
  assign n3258 = n3026 & n19678 ;
  assign n3259 = n3257 | n3258 ;
  assign n19679 = ~n3259 ;
  assign n3260 = n3254 & n19679 ;
  assign n3261 = n3253 | n3260 ;
  assign n3262 = x85 & n3261 ;
  assign n3263 = x85 | n3261 ;
  assign n19680 = ~n3029 ;
  assign n3264 = n19680 & n3030 ;
  assign n3265 = n167 & n3264 ;
  assign n3266 = n19598 & n3265 ;
  assign n19681 = ~n3265 ;
  assign n3267 = n3035 & n19681 ;
  assign n3268 = n3266 | n3267 ;
  assign n19682 = ~n3268 ;
  assign n3269 = n3263 & n19682 ;
  assign n3270 = n3262 | n3269 ;
  assign n3271 = x86 & n3270 ;
  assign n3272 = x86 | n3270 ;
  assign n19683 = ~n3038 ;
  assign n3273 = n19683 & n3039 ;
  assign n3274 = n167 & n3273 ;
  assign n3275 = n19601 & n3274 ;
  assign n19684 = ~n3274 ;
  assign n3276 = n3044 & n19684 ;
  assign n3277 = n3275 | n3276 ;
  assign n19685 = ~n3277 ;
  assign n3278 = n3272 & n19685 ;
  assign n3279 = n3271 | n3278 ;
  assign n3280 = x87 & n3279 ;
  assign n3281 = x87 | n3279 ;
  assign n19686 = ~n3047 ;
  assign n3282 = n19686 & n3048 ;
  assign n3283 = n167 & n3282 ;
  assign n3284 = n19604 & n3283 ;
  assign n19687 = ~n3283 ;
  assign n3285 = n3053 & n19687 ;
  assign n3286 = n3284 | n3285 ;
  assign n19688 = ~n3286 ;
  assign n3287 = n3281 & n19688 ;
  assign n3288 = n3280 | n3287 ;
  assign n3289 = x88 & n3288 ;
  assign n3290 = x88 | n3288 ;
  assign n19689 = ~n3056 ;
  assign n3291 = n19689 & n3057 ;
  assign n3292 = n167 & n3291 ;
  assign n3293 = n19607 & n3292 ;
  assign n19690 = ~n3292 ;
  assign n3294 = n3062 & n19690 ;
  assign n3295 = n3293 | n3294 ;
  assign n19691 = ~n3295 ;
  assign n3296 = n3290 & n19691 ;
  assign n3297 = n3289 | n3296 ;
  assign n3299 = x89 | n3297 ;
  assign n19692 = ~n3081 ;
  assign n3300 = n19692 & n3299 ;
  assign n3298 = x89 & n3297 ;
  assign n19693 = ~n3067 ;
  assign n3068 = x90 & n19693 ;
  assign n3301 = n18443 | n3068 ;
  assign n3302 = n3298 | n3301 ;
  assign n3303 = n3300 | n3302 ;
  assign n3304 = n21884 | n3074 ;
  assign n3305 = n3073 & n3304 ;
  assign n19694 = ~n3305 ;
  assign n3306 = n3303 & n19694 ;
  assign n19695 = ~n3298 ;
  assign n3307 = n19695 & n3299 ;
  assign n166 = ~n3306 ;
  assign n3308 = n166 & n3307 ;
  assign n3309 = n3081 & n3308 ;
  assign n3310 = n3081 | n3308 ;
  assign n19697 = ~n3309 ;
  assign n3311 = n19697 & n3310 ;
  assign n19698 = ~x36 ;
  assign n3312 = n19698 & x64 ;
  assign n3313 = x65 | n3312 ;
  assign n3314 = x64 & n166 ;
  assign n19699 = ~n3314 ;
  assign n3315 = x37 & n19699 ;
  assign n3316 = n3082 & n166 ;
  assign n3317 = n3315 | n3316 ;
  assign n3318 = x65 & n3312 ;
  assign n19700 = ~n3318 ;
  assign n3319 = n3317 & n19700 ;
  assign n19701 = ~n3319 ;
  assign n3320 = n3313 & n19701 ;
  assign n3321 = x66 & n3320 ;
  assign n3322 = n19618 & n3084 ;
  assign n3323 = n166 & n3322 ;
  assign n3324 = n3088 & n3323 ;
  assign n3325 = n3088 | n3323 ;
  assign n19702 = ~n3324 ;
  assign n3326 = n19702 & n3325 ;
  assign n3327 = x66 | n3320 ;
  assign n19703 = ~n3326 ;
  assign n3328 = n19703 & n3327 ;
  assign n3329 = n3321 | n3328 ;
  assign n3330 = x67 & n3329 ;
  assign n3331 = x67 | n3329 ;
  assign n19704 = ~n3091 ;
  assign n3332 = n19704 & n3092 ;
  assign n3333 = n166 & n3332 ;
  assign n3334 = n3097 & n3333 ;
  assign n3335 = n3097 | n3333 ;
  assign n19705 = ~n3334 ;
  assign n3336 = n19705 & n3335 ;
  assign n19706 = ~n3336 ;
  assign n3337 = n3331 & n19706 ;
  assign n3338 = n3330 | n3337 ;
  assign n3339 = x68 & n3338 ;
  assign n3340 = x68 | n3338 ;
  assign n19707 = ~n3100 ;
  assign n3341 = n19707 & n3101 ;
  assign n3342 = n166 & n3341 ;
  assign n3343 = n3106 & n3342 ;
  assign n3344 = n3106 | n3342 ;
  assign n19708 = ~n3343 ;
  assign n3345 = n19708 & n3344 ;
  assign n19709 = ~n3345 ;
  assign n3346 = n3340 & n19709 ;
  assign n3347 = n3339 | n3346 ;
  assign n3348 = x69 & n3347 ;
  assign n3349 = x69 | n3347 ;
  assign n3350 = n19627 & n3110 ;
  assign n3351 = n166 & n3350 ;
  assign n19710 = ~n3115 ;
  assign n3352 = n19710 & n3351 ;
  assign n19711 = ~n3351 ;
  assign n3353 = n3115 & n19711 ;
  assign n3354 = n3352 | n3353 ;
  assign n19712 = ~n3354 ;
  assign n3355 = n3349 & n19712 ;
  assign n3356 = n3348 | n3355 ;
  assign n3357 = x70 & n3356 ;
  assign n3358 = x70 | n3356 ;
  assign n3359 = n3118 & n19631 ;
  assign n3360 = n166 & n3359 ;
  assign n3361 = n3124 & n3360 ;
  assign n3362 = n3124 | n3360 ;
  assign n19713 = ~n3361 ;
  assign n3363 = n19713 & n3362 ;
  assign n19714 = ~n3363 ;
  assign n3364 = n3358 & n19714 ;
  assign n3365 = n3357 | n3364 ;
  assign n3366 = x71 & n3365 ;
  assign n3367 = x71 | n3365 ;
  assign n3368 = n3127 & n19635 ;
  assign n3369 = n166 & n3368 ;
  assign n3370 = n3133 & n3369 ;
  assign n3371 = n3133 | n3369 ;
  assign n19715 = ~n3370 ;
  assign n3372 = n19715 & n3371 ;
  assign n19716 = ~n3372 ;
  assign n3373 = n3367 & n19716 ;
  assign n3374 = n3366 | n3373 ;
  assign n3375 = x72 & n3374 ;
  assign n3376 = x72 | n3374 ;
  assign n3377 = n3136 & n19639 ;
  assign n3378 = n166 & n3377 ;
  assign n3379 = n3142 & n3378 ;
  assign n3380 = n3142 | n3378 ;
  assign n19717 = ~n3379 ;
  assign n3381 = n19717 & n3380 ;
  assign n19718 = ~n3381 ;
  assign n3382 = n3376 & n19718 ;
  assign n3383 = n3375 | n3382 ;
  assign n3384 = x73 & n3383 ;
  assign n3385 = x73 | n3383 ;
  assign n19719 = ~n3146 ;
  assign n3386 = n3145 & n19719 ;
  assign n3387 = n166 & n3386 ;
  assign n3388 = n3151 & n3387 ;
  assign n3389 = n3151 | n3387 ;
  assign n19720 = ~n3388 ;
  assign n3390 = n19720 & n3389 ;
  assign n19721 = ~n3390 ;
  assign n3391 = n3385 & n19721 ;
  assign n3392 = n3384 | n3391 ;
  assign n3393 = x74 & n3392 ;
  assign n3394 = x74 | n3392 ;
  assign n19722 = ~n3154 ;
  assign n3395 = n19722 & n3155 ;
  assign n3396 = n166 & n3395 ;
  assign n3397 = n3160 & n3396 ;
  assign n3398 = n3160 | n3396 ;
  assign n19723 = ~n3397 ;
  assign n3399 = n19723 & n3398 ;
  assign n19724 = ~n3399 ;
  assign n3400 = n3394 & n19724 ;
  assign n3401 = n3393 | n3400 ;
  assign n3402 = x75 & n3401 ;
  assign n3403 = x75 | n3401 ;
  assign n19725 = ~n3163 ;
  assign n3404 = n19725 & n3164 ;
  assign n3405 = n166 & n3404 ;
  assign n3406 = n19649 & n3405 ;
  assign n19726 = ~n3405 ;
  assign n3407 = n3169 & n19726 ;
  assign n3408 = n3406 | n3407 ;
  assign n19727 = ~n3408 ;
  assign n3409 = n3403 & n19727 ;
  assign n3410 = n3402 | n3409 ;
  assign n3411 = x76 & n3410 ;
  assign n3412 = x76 | n3410 ;
  assign n19728 = ~n3172 ;
  assign n3413 = n19728 & n3173 ;
  assign n3414 = n166 & n3413 ;
  assign n3415 = n3178 & n3414 ;
  assign n3416 = n3178 | n3414 ;
  assign n19729 = ~n3415 ;
  assign n3417 = n19729 & n3416 ;
  assign n19730 = ~n3417 ;
  assign n3418 = n3412 & n19730 ;
  assign n3419 = n3411 | n3418 ;
  assign n3420 = x77 & n3419 ;
  assign n3421 = x77 | n3419 ;
  assign n19731 = ~n3181 ;
  assign n3422 = n19731 & n3182 ;
  assign n3423 = n166 & n3422 ;
  assign n3424 = n3187 & n3423 ;
  assign n3425 = n3187 | n3423 ;
  assign n19732 = ~n3424 ;
  assign n3426 = n19732 & n3425 ;
  assign n19733 = ~n3426 ;
  assign n3427 = n3421 & n19733 ;
  assign n3428 = n3420 | n3427 ;
  assign n3429 = x78 & n3428 ;
  assign n3430 = x78 | n3428 ;
  assign n19734 = ~n3190 ;
  assign n3431 = n19734 & n3191 ;
  assign n3432 = n166 & n3431 ;
  assign n3433 = n3196 & n3432 ;
  assign n3434 = n3196 | n3432 ;
  assign n19735 = ~n3433 ;
  assign n3435 = n19735 & n3434 ;
  assign n19736 = ~n3435 ;
  assign n3436 = n3430 & n19736 ;
  assign n3437 = n3429 | n3436 ;
  assign n3438 = x79 & n3437 ;
  assign n3439 = x79 | n3437 ;
  assign n19737 = ~n3199 ;
  assign n3440 = n19737 & n3200 ;
  assign n3441 = n166 & n3440 ;
  assign n3442 = n3205 & n3441 ;
  assign n3443 = n3205 | n3441 ;
  assign n19738 = ~n3442 ;
  assign n3444 = n19738 & n3443 ;
  assign n19739 = ~n3444 ;
  assign n3445 = n3439 & n19739 ;
  assign n3446 = n3438 | n3445 ;
  assign n3447 = x80 & n3446 ;
  assign n3448 = x80 | n3446 ;
  assign n19740 = ~n3208 ;
  assign n3449 = n19740 & n3209 ;
  assign n3450 = n166 & n3449 ;
  assign n3451 = n3214 & n3450 ;
  assign n3452 = n3214 | n3450 ;
  assign n19741 = ~n3451 ;
  assign n3453 = n19741 & n3452 ;
  assign n19742 = ~n3453 ;
  assign n3454 = n3448 & n19742 ;
  assign n3455 = n3447 | n3454 ;
  assign n3456 = x81 & n3455 ;
  assign n3457 = x81 | n3455 ;
  assign n19743 = ~n3217 ;
  assign n3458 = n19743 & n3218 ;
  assign n3459 = n166 & n3458 ;
  assign n3460 = n3223 & n3459 ;
  assign n3461 = n3223 | n3459 ;
  assign n19744 = ~n3460 ;
  assign n3462 = n19744 & n3461 ;
  assign n19745 = ~n3462 ;
  assign n3463 = n3457 & n19745 ;
  assign n3464 = n3456 | n3463 ;
  assign n3465 = x82 & n3464 ;
  assign n3466 = x82 | n3464 ;
  assign n19746 = ~n3226 ;
  assign n3467 = n19746 & n3227 ;
  assign n3468 = n166 & n3467 ;
  assign n3469 = n3232 & n3468 ;
  assign n3470 = n3232 | n3468 ;
  assign n19747 = ~n3469 ;
  assign n3471 = n19747 & n3470 ;
  assign n19748 = ~n3471 ;
  assign n3472 = n3466 & n19748 ;
  assign n3473 = n3465 | n3472 ;
  assign n3474 = x83 & n3473 ;
  assign n3475 = x83 | n3473 ;
  assign n19749 = ~n3235 ;
  assign n3476 = n19749 & n3236 ;
  assign n3477 = n166 & n3476 ;
  assign n3478 = n3241 & n3477 ;
  assign n3479 = n3241 | n3477 ;
  assign n19750 = ~n3478 ;
  assign n3480 = n19750 & n3479 ;
  assign n19751 = ~n3480 ;
  assign n3481 = n3475 & n19751 ;
  assign n3482 = n3474 | n3481 ;
  assign n3483 = x84 & n3482 ;
  assign n3484 = x84 | n3482 ;
  assign n19752 = ~n3244 ;
  assign n3485 = n19752 & n3245 ;
  assign n3486 = n166 & n3485 ;
  assign n3487 = n3250 & n3486 ;
  assign n3488 = n3250 | n3486 ;
  assign n19753 = ~n3487 ;
  assign n3489 = n19753 & n3488 ;
  assign n19754 = ~n3489 ;
  assign n3490 = n3484 & n19754 ;
  assign n3491 = n3483 | n3490 ;
  assign n3492 = x85 & n3491 ;
  assign n3493 = x85 | n3491 ;
  assign n19755 = ~n3253 ;
  assign n3494 = n19755 & n3254 ;
  assign n3495 = n166 & n3494 ;
  assign n3496 = n3259 & n3495 ;
  assign n3497 = n3259 | n3495 ;
  assign n19756 = ~n3496 ;
  assign n3498 = n19756 & n3497 ;
  assign n19757 = ~n3498 ;
  assign n3499 = n3493 & n19757 ;
  assign n3500 = n3492 | n3499 ;
  assign n3501 = x86 & n3500 ;
  assign n3502 = x86 | n3500 ;
  assign n19758 = ~n3262 ;
  assign n3503 = n19758 & n3263 ;
  assign n3504 = n166 & n3503 ;
  assign n3505 = n3268 & n3504 ;
  assign n3506 = n3268 | n3504 ;
  assign n19759 = ~n3505 ;
  assign n3507 = n19759 & n3506 ;
  assign n19760 = ~n3507 ;
  assign n3508 = n3502 & n19760 ;
  assign n3509 = n3501 | n3508 ;
  assign n3510 = x87 & n3509 ;
  assign n3511 = x87 | n3509 ;
  assign n19761 = ~n3271 ;
  assign n3512 = n19761 & n3272 ;
  assign n3513 = n166 & n3512 ;
  assign n3514 = n3277 & n3513 ;
  assign n3515 = n3277 | n3513 ;
  assign n19762 = ~n3514 ;
  assign n3516 = n19762 & n3515 ;
  assign n19763 = ~n3516 ;
  assign n3517 = n3511 & n19763 ;
  assign n3518 = n3510 | n3517 ;
  assign n3519 = x88 & n3518 ;
  assign n3520 = x88 | n3518 ;
  assign n19764 = ~n3280 ;
  assign n3521 = n19764 & n3281 ;
  assign n3522 = n166 & n3521 ;
  assign n3523 = n3286 & n3522 ;
  assign n3524 = n3286 | n3522 ;
  assign n19765 = ~n3523 ;
  assign n3525 = n19765 & n3524 ;
  assign n19766 = ~n3525 ;
  assign n3526 = n3520 & n19766 ;
  assign n3527 = n3519 | n3526 ;
  assign n3528 = x89 & n3527 ;
  assign n3529 = x89 | n3527 ;
  assign n19767 = ~n3289 ;
  assign n3530 = n19767 & n3290 ;
  assign n3531 = n166 & n3530 ;
  assign n3532 = n3295 & n3531 ;
  assign n3533 = n3295 | n3531 ;
  assign n19768 = ~n3532 ;
  assign n3534 = n19768 & n3533 ;
  assign n19769 = ~n3534 ;
  assign n3535 = n3529 & n19769 ;
  assign n3536 = n3528 | n3535 ;
  assign n3537 = x90 & n3536 ;
  assign n3538 = x90 | n3536 ;
  assign n19770 = ~n3311 ;
  assign n3539 = n19770 & n3538 ;
  assign n3540 = n3537 | n3539 ;
  assign n3542 = x91 & n3540 ;
  assign n3543 = n18438 | n3542 ;
  assign n3541 = x91 | n3540 ;
  assign n3069 = n18448 & n3067 ;
  assign n3544 = n3069 & n3303 ;
  assign n3546 = n21884 | n3544 ;
  assign n19771 = ~n3546 ;
  assign n3547 = n3541 & n19771 ;
  assign n3548 = n3543 | n3547 ;
  assign n19772 = ~n3537 ;
  assign n3549 = n19772 & n3538 ;
  assign n165 = ~n3548 ;
  assign n3550 = n165 & n3549 ;
  assign n3551 = n19770 & n3550 ;
  assign n19774 = ~n3550 ;
  assign n3552 = n3311 & n19774 ;
  assign n3553 = n3551 | n3552 ;
  assign n19775 = ~x35 ;
  assign n3554 = n19775 & x64 ;
  assign n3556 = x65 | n3554 ;
  assign n3555 = x65 & n3554 ;
  assign n3557 = x64 & n165 ;
  assign n3558 = x36 & n3557 ;
  assign n3559 = x36 | n3557 ;
  assign n19776 = ~n3558 ;
  assign n3560 = n19776 & n3559 ;
  assign n19777 = ~n3555 ;
  assign n3561 = n19777 & n3560 ;
  assign n19778 = ~n3561 ;
  assign n3562 = n3556 & n19778 ;
  assign n3563 = x66 | n3562 ;
  assign n3564 = x66 & n3562 ;
  assign n3565 = n3313 & n165 ;
  assign n3566 = n19700 & n3565 ;
  assign n3567 = n3317 | n3566 ;
  assign n3568 = n3319 & n3565 ;
  assign n19779 = ~n3568 ;
  assign n3569 = n3567 & n19779 ;
  assign n19780 = ~n3564 ;
  assign n3570 = n19780 & n3569 ;
  assign n19781 = ~n3570 ;
  assign n3571 = n3563 & n19781 ;
  assign n3572 = x67 | n3571 ;
  assign n3573 = x67 & n3571 ;
  assign n19782 = ~n3321 ;
  assign n3574 = n19782 & n3327 ;
  assign n3575 = n165 & n3574 ;
  assign n3576 = n3326 & n3575 ;
  assign n3577 = n3326 | n3575 ;
  assign n19783 = ~n3576 ;
  assign n3578 = n19783 & n3577 ;
  assign n19784 = ~n3573 ;
  assign n3579 = n19784 & n3578 ;
  assign n19785 = ~n3579 ;
  assign n3580 = n3572 & n19785 ;
  assign n3581 = x68 | n3580 ;
  assign n3582 = x68 & n3580 ;
  assign n19786 = ~n3330 ;
  assign n3583 = n19786 & n3331 ;
  assign n3584 = n165 & n3583 ;
  assign n3585 = n3336 & n3584 ;
  assign n3586 = n3336 | n3584 ;
  assign n19787 = ~n3585 ;
  assign n3587 = n19787 & n3586 ;
  assign n19788 = ~n3582 ;
  assign n3588 = n19788 & n3587 ;
  assign n19789 = ~n3588 ;
  assign n3589 = n3581 & n19789 ;
  assign n3590 = x69 | n3589 ;
  assign n3591 = x69 & n3589 ;
  assign n19790 = ~n3339 ;
  assign n3592 = n19790 & n3340 ;
  assign n3593 = n165 & n3592 ;
  assign n3594 = n3345 & n3593 ;
  assign n3595 = n3345 | n3593 ;
  assign n19791 = ~n3594 ;
  assign n3596 = n19791 & n3595 ;
  assign n19792 = ~n3591 ;
  assign n3597 = n19792 & n3596 ;
  assign n19793 = ~n3597 ;
  assign n3598 = n3590 & n19793 ;
  assign n3599 = x70 | n3598 ;
  assign n3600 = x70 & n3598 ;
  assign n19794 = ~n3348 ;
  assign n3601 = n19794 & n3349 ;
  assign n3602 = n165 & n3601 ;
  assign n3603 = n19712 & n3602 ;
  assign n19795 = ~n3602 ;
  assign n3604 = n3354 & n19795 ;
  assign n3605 = n3603 | n3604 ;
  assign n19796 = ~n3600 ;
  assign n3606 = n19796 & n3605 ;
  assign n19797 = ~n3606 ;
  assign n3607 = n3599 & n19797 ;
  assign n3608 = x71 | n3607 ;
  assign n3609 = x71 & n3607 ;
  assign n19798 = ~n3357 ;
  assign n3610 = n19798 & n3358 ;
  assign n3611 = n165 & n3610 ;
  assign n3612 = n3363 & n3611 ;
  assign n3613 = n3363 | n3611 ;
  assign n19799 = ~n3612 ;
  assign n3614 = n19799 & n3613 ;
  assign n19800 = ~n3609 ;
  assign n3615 = n19800 & n3614 ;
  assign n19801 = ~n3615 ;
  assign n3616 = n3608 & n19801 ;
  assign n3617 = x72 | n3616 ;
  assign n3618 = x72 & n3616 ;
  assign n19802 = ~n3366 ;
  assign n3619 = n19802 & n3367 ;
  assign n3620 = n165 & n3619 ;
  assign n3621 = n3372 & n3620 ;
  assign n3622 = n3372 | n3620 ;
  assign n19803 = ~n3621 ;
  assign n3623 = n19803 & n3622 ;
  assign n19804 = ~n3618 ;
  assign n3624 = n19804 & n3623 ;
  assign n19805 = ~n3624 ;
  assign n3625 = n3617 & n19805 ;
  assign n3626 = x73 | n3625 ;
  assign n3627 = x73 & n3625 ;
  assign n19806 = ~n3375 ;
  assign n3628 = n19806 & n3376 ;
  assign n3629 = n165 & n3628 ;
  assign n3630 = n3381 & n3629 ;
  assign n3631 = n3381 | n3629 ;
  assign n19807 = ~n3630 ;
  assign n3632 = n19807 & n3631 ;
  assign n19808 = ~n3627 ;
  assign n3633 = n19808 & n3632 ;
  assign n19809 = ~n3633 ;
  assign n3634 = n3626 & n19809 ;
  assign n3635 = x74 | n3634 ;
  assign n3636 = x74 & n3634 ;
  assign n19810 = ~n3384 ;
  assign n3637 = n19810 & n3385 ;
  assign n3638 = n165 & n3637 ;
  assign n3639 = n3390 & n3638 ;
  assign n3640 = n3390 | n3638 ;
  assign n19811 = ~n3639 ;
  assign n3641 = n19811 & n3640 ;
  assign n19812 = ~n3636 ;
  assign n3642 = n19812 & n3641 ;
  assign n19813 = ~n3642 ;
  assign n3643 = n3635 & n19813 ;
  assign n3644 = x75 | n3643 ;
  assign n3645 = x75 & n3643 ;
  assign n19814 = ~n3393 ;
  assign n3646 = n19814 & n3394 ;
  assign n3647 = n165 & n3646 ;
  assign n3648 = n19724 & n3647 ;
  assign n19815 = ~n3647 ;
  assign n3649 = n3399 & n19815 ;
  assign n3650 = n3648 | n3649 ;
  assign n19816 = ~n3645 ;
  assign n3651 = n19816 & n3650 ;
  assign n19817 = ~n3651 ;
  assign n3652 = n3644 & n19817 ;
  assign n3653 = x76 | n3652 ;
  assign n3654 = x76 & n3652 ;
  assign n19818 = ~n3402 ;
  assign n3655 = n19818 & n3403 ;
  assign n3656 = n165 & n3655 ;
  assign n3657 = n19727 & n3656 ;
  assign n19819 = ~n3656 ;
  assign n3658 = n3408 & n19819 ;
  assign n3659 = n3657 | n3658 ;
  assign n19820 = ~n3654 ;
  assign n3660 = n19820 & n3659 ;
  assign n19821 = ~n3660 ;
  assign n3661 = n3653 & n19821 ;
  assign n3662 = x77 | n3661 ;
  assign n3663 = x77 & n3661 ;
  assign n19822 = ~n3411 ;
  assign n3664 = n19822 & n3412 ;
  assign n3665 = n165 & n3664 ;
  assign n3666 = n3417 & n3665 ;
  assign n3667 = n3417 | n3665 ;
  assign n19823 = ~n3666 ;
  assign n3668 = n19823 & n3667 ;
  assign n19824 = ~n3663 ;
  assign n3669 = n19824 & n3668 ;
  assign n19825 = ~n3669 ;
  assign n3670 = n3662 & n19825 ;
  assign n3671 = x78 | n3670 ;
  assign n3672 = x78 & n3670 ;
  assign n19826 = ~n3420 ;
  assign n3673 = n19826 & n3421 ;
  assign n3674 = n165 & n3673 ;
  assign n3675 = n3426 & n3674 ;
  assign n3676 = n3426 | n3674 ;
  assign n19827 = ~n3675 ;
  assign n3677 = n19827 & n3676 ;
  assign n19828 = ~n3672 ;
  assign n3678 = n19828 & n3677 ;
  assign n19829 = ~n3678 ;
  assign n3679 = n3671 & n19829 ;
  assign n3680 = x79 | n3679 ;
  assign n3681 = x79 & n3679 ;
  assign n19830 = ~n3429 ;
  assign n3682 = n19830 & n3430 ;
  assign n3683 = n165 & n3682 ;
  assign n3684 = n3435 & n3683 ;
  assign n3685 = n3435 | n3683 ;
  assign n19831 = ~n3684 ;
  assign n3686 = n19831 & n3685 ;
  assign n19832 = ~n3681 ;
  assign n3687 = n19832 & n3686 ;
  assign n19833 = ~n3687 ;
  assign n3688 = n3680 & n19833 ;
  assign n3689 = x80 | n3688 ;
  assign n3690 = x80 & n3688 ;
  assign n19834 = ~n3438 ;
  assign n3691 = n19834 & n3439 ;
  assign n3692 = n165 & n3691 ;
  assign n3693 = n3444 & n3692 ;
  assign n3694 = n3444 | n3692 ;
  assign n19835 = ~n3693 ;
  assign n3695 = n19835 & n3694 ;
  assign n19836 = ~n3690 ;
  assign n3696 = n19836 & n3695 ;
  assign n19837 = ~n3696 ;
  assign n3697 = n3689 & n19837 ;
  assign n3698 = x81 | n3697 ;
  assign n3699 = x81 & n3697 ;
  assign n19838 = ~n3447 ;
  assign n3700 = n19838 & n3448 ;
  assign n3701 = n165 & n3700 ;
  assign n3702 = n3453 & n3701 ;
  assign n3703 = n3453 | n3701 ;
  assign n19839 = ~n3702 ;
  assign n3704 = n19839 & n3703 ;
  assign n19840 = ~n3699 ;
  assign n3705 = n19840 & n3704 ;
  assign n19841 = ~n3705 ;
  assign n3706 = n3698 & n19841 ;
  assign n3707 = x82 | n3706 ;
  assign n3708 = x82 & n3706 ;
  assign n19842 = ~n3456 ;
  assign n3709 = n19842 & n3457 ;
  assign n3710 = n165 & n3709 ;
  assign n3711 = n3462 & n3710 ;
  assign n3712 = n3462 | n3710 ;
  assign n19843 = ~n3711 ;
  assign n3713 = n19843 & n3712 ;
  assign n19844 = ~n3708 ;
  assign n3714 = n19844 & n3713 ;
  assign n19845 = ~n3714 ;
  assign n3715 = n3707 & n19845 ;
  assign n3716 = x83 | n3715 ;
  assign n3717 = x83 & n3715 ;
  assign n19846 = ~n3465 ;
  assign n3718 = n19846 & n3466 ;
  assign n3719 = n165 & n3718 ;
  assign n3720 = n3471 & n3719 ;
  assign n3721 = n3471 | n3719 ;
  assign n19847 = ~n3720 ;
  assign n3722 = n19847 & n3721 ;
  assign n19848 = ~n3717 ;
  assign n3723 = n19848 & n3722 ;
  assign n19849 = ~n3723 ;
  assign n3724 = n3716 & n19849 ;
  assign n3725 = x84 | n3724 ;
  assign n3726 = x84 & n3724 ;
  assign n19850 = ~n3474 ;
  assign n3727 = n19850 & n3475 ;
  assign n3728 = n165 & n3727 ;
  assign n3729 = n3480 & n3728 ;
  assign n3730 = n3480 | n3728 ;
  assign n19851 = ~n3729 ;
  assign n3731 = n19851 & n3730 ;
  assign n19852 = ~n3726 ;
  assign n3732 = n19852 & n3731 ;
  assign n19853 = ~n3732 ;
  assign n3733 = n3725 & n19853 ;
  assign n3734 = x85 | n3733 ;
  assign n3735 = x85 & n3733 ;
  assign n19854 = ~n3483 ;
  assign n3736 = n19854 & n3484 ;
  assign n3737 = n165 & n3736 ;
  assign n3738 = n3489 & n3737 ;
  assign n3739 = n3489 | n3737 ;
  assign n19855 = ~n3738 ;
  assign n3740 = n19855 & n3739 ;
  assign n19856 = ~n3735 ;
  assign n3741 = n19856 & n3740 ;
  assign n19857 = ~n3741 ;
  assign n3742 = n3734 & n19857 ;
  assign n3743 = x86 | n3742 ;
  assign n3744 = x86 & n3742 ;
  assign n19858 = ~n3492 ;
  assign n3745 = n19858 & n3493 ;
  assign n3746 = n165 & n3745 ;
  assign n3747 = n3498 & n3746 ;
  assign n3748 = n3498 | n3746 ;
  assign n19859 = ~n3747 ;
  assign n3749 = n19859 & n3748 ;
  assign n19860 = ~n3744 ;
  assign n3750 = n19860 & n3749 ;
  assign n19861 = ~n3750 ;
  assign n3751 = n3743 & n19861 ;
  assign n3752 = x87 | n3751 ;
  assign n3753 = x87 & n3751 ;
  assign n19862 = ~n3501 ;
  assign n3754 = n19862 & n3502 ;
  assign n3755 = n165 & n3754 ;
  assign n3756 = n3507 & n3755 ;
  assign n3757 = n3507 | n3755 ;
  assign n19863 = ~n3756 ;
  assign n3758 = n19863 & n3757 ;
  assign n19864 = ~n3753 ;
  assign n3759 = n19864 & n3758 ;
  assign n19865 = ~n3759 ;
  assign n3760 = n3752 & n19865 ;
  assign n3761 = x88 | n3760 ;
  assign n3762 = x88 & n3760 ;
  assign n19866 = ~n3510 ;
  assign n3763 = n19866 & n3511 ;
  assign n3764 = n165 & n3763 ;
  assign n3765 = n3516 & n3764 ;
  assign n3766 = n3516 | n3764 ;
  assign n19867 = ~n3765 ;
  assign n3767 = n19867 & n3766 ;
  assign n19868 = ~n3762 ;
  assign n3768 = n19868 & n3767 ;
  assign n19869 = ~n3768 ;
  assign n3769 = n3761 & n19869 ;
  assign n3770 = x89 | n3769 ;
  assign n3771 = x89 & n3769 ;
  assign n19870 = ~n3519 ;
  assign n3772 = n19870 & n3520 ;
  assign n3773 = n165 & n3772 ;
  assign n3774 = n3525 & n3773 ;
  assign n3775 = n3525 | n3773 ;
  assign n19871 = ~n3774 ;
  assign n3776 = n19871 & n3775 ;
  assign n19872 = ~n3771 ;
  assign n3777 = n19872 & n3776 ;
  assign n19873 = ~n3777 ;
  assign n3778 = n3770 & n19873 ;
  assign n3779 = x90 | n3778 ;
  assign n3780 = x90 & n3778 ;
  assign n19874 = ~n3528 ;
  assign n3781 = n19874 & n3529 ;
  assign n3782 = n165 & n3781 ;
  assign n3783 = n3534 & n3782 ;
  assign n3784 = n3534 | n3782 ;
  assign n19875 = ~n3783 ;
  assign n3785 = n19875 & n3784 ;
  assign n19876 = ~n3780 ;
  assign n3786 = n19876 & n3785 ;
  assign n19877 = ~n3786 ;
  assign n3787 = n3779 & n19877 ;
  assign n3789 = x91 & n3787 ;
  assign n19878 = ~n3789 ;
  assign n3790 = n3553 & n19878 ;
  assign n3788 = x91 | n3787 ;
  assign n3545 = n3543 & n3544 ;
  assign n3791 = n21884 | n3545 ;
  assign n19879 = ~x92 ;
  assign n3792 = n19879 & n3791 ;
  assign n19880 = ~n3792 ;
  assign n3793 = n3788 & n19880 ;
  assign n19881 = ~n3790 ;
  assign n3794 = n19881 & n3793 ;
  assign n3795 = n18433 | n3794 ;
  assign n3796 = x92 & n19771 ;
  assign n3797 = n3795 | n3796 ;
  assign n3798 = n3788 & n19878 ;
  assign n164 = ~n3797 ;
  assign n3799 = n164 & n3798 ;
  assign n19883 = ~n3553 ;
  assign n3800 = n19883 & n3799 ;
  assign n19884 = ~n3799 ;
  assign n3801 = n3553 & n19884 ;
  assign n3802 = n3800 | n3801 ;
  assign n19885 = ~x34 ;
  assign n3803 = n19885 & x64 ;
  assign n3805 = x65 | n3803 ;
  assign n3804 = x65 & n3803 ;
  assign n3806 = x64 & n164 ;
  assign n3807 = x35 & n3806 ;
  assign n3808 = x35 | n3806 ;
  assign n19886 = ~n3807 ;
  assign n3809 = n19886 & n3808 ;
  assign n19887 = ~n3804 ;
  assign n3810 = n19887 & n3809 ;
  assign n19888 = ~n3810 ;
  assign n3811 = n3805 & n19888 ;
  assign n3812 = x66 & n3811 ;
  assign n3813 = x66 | n3811 ;
  assign n3814 = n19777 & n3556 ;
  assign n3815 = n164 & n3814 ;
  assign n3816 = n3560 & n3815 ;
  assign n3817 = n3560 | n3815 ;
  assign n19889 = ~n3816 ;
  assign n3818 = n19889 & n3817 ;
  assign n19890 = ~n3818 ;
  assign n3819 = n3813 & n19890 ;
  assign n3820 = n3812 | n3819 ;
  assign n3821 = x67 & n3820 ;
  assign n3822 = x67 | n3820 ;
  assign n3823 = n3563 & n19780 ;
  assign n3824 = n164 & n3823 ;
  assign n19891 = ~n3569 ;
  assign n3825 = n19891 & n3824 ;
  assign n19892 = ~n3824 ;
  assign n3826 = n3569 & n19892 ;
  assign n3827 = n3825 | n3826 ;
  assign n19893 = ~n3827 ;
  assign n3828 = n3822 & n19893 ;
  assign n3829 = n3821 | n3828 ;
  assign n3830 = x68 & n3829 ;
  assign n3831 = x68 | n3829 ;
  assign n3832 = n3572 & n19784 ;
  assign n3833 = n164 & n3832 ;
  assign n19894 = ~n3578 ;
  assign n3834 = n19894 & n3833 ;
  assign n19895 = ~n3833 ;
  assign n3835 = n3578 & n19895 ;
  assign n3836 = n3834 | n3835 ;
  assign n19896 = ~n3836 ;
  assign n3837 = n3831 & n19896 ;
  assign n3838 = n3830 | n3837 ;
  assign n3839 = x69 & n3838 ;
  assign n3840 = x69 | n3838 ;
  assign n3841 = n3581 & n19788 ;
  assign n3842 = n164 & n3841 ;
  assign n19897 = ~n3587 ;
  assign n3843 = n19897 & n3842 ;
  assign n19898 = ~n3842 ;
  assign n3844 = n3587 & n19898 ;
  assign n3845 = n3843 | n3844 ;
  assign n19899 = ~n3845 ;
  assign n3846 = n3840 & n19899 ;
  assign n3847 = n3839 | n3846 ;
  assign n3848 = x70 & n3847 ;
  assign n3849 = x70 | n3847 ;
  assign n3850 = n3590 & n19792 ;
  assign n3851 = n164 & n3850 ;
  assign n3852 = n3596 & n3851 ;
  assign n3853 = n3596 | n3851 ;
  assign n19900 = ~n3852 ;
  assign n3854 = n19900 & n3853 ;
  assign n19901 = ~n3854 ;
  assign n3855 = n3849 & n19901 ;
  assign n3856 = n3848 | n3855 ;
  assign n3857 = x71 & n3856 ;
  assign n3858 = x71 | n3856 ;
  assign n3859 = n3599 & n19796 ;
  assign n3860 = n164 & n3859 ;
  assign n19902 = ~n3605 ;
  assign n3861 = n19902 & n3860 ;
  assign n19903 = ~n3860 ;
  assign n3862 = n3605 & n19903 ;
  assign n3863 = n3861 | n3862 ;
  assign n19904 = ~n3863 ;
  assign n3864 = n3858 & n19904 ;
  assign n3865 = n3857 | n3864 ;
  assign n3866 = x72 & n3865 ;
  assign n3867 = x72 | n3865 ;
  assign n3868 = n3608 & n19800 ;
  assign n3869 = n164 & n3868 ;
  assign n19905 = ~n3614 ;
  assign n3870 = n19905 & n3869 ;
  assign n19906 = ~n3869 ;
  assign n3871 = n3614 & n19906 ;
  assign n3872 = n3870 | n3871 ;
  assign n19907 = ~n3872 ;
  assign n3873 = n3867 & n19907 ;
  assign n3874 = n3866 | n3873 ;
  assign n3875 = x73 & n3874 ;
  assign n3876 = x73 | n3874 ;
  assign n3877 = n3617 & n19804 ;
  assign n3878 = n164 & n3877 ;
  assign n19908 = ~n3623 ;
  assign n3879 = n19908 & n3878 ;
  assign n19909 = ~n3878 ;
  assign n3880 = n3623 & n19909 ;
  assign n3881 = n3879 | n3880 ;
  assign n19910 = ~n3881 ;
  assign n3882 = n3876 & n19910 ;
  assign n3883 = n3875 | n3882 ;
  assign n3884 = x74 & n3883 ;
  assign n3885 = x74 | n3883 ;
  assign n3886 = n3626 & n19808 ;
  assign n3887 = n164 & n3886 ;
  assign n19911 = ~n3632 ;
  assign n3888 = n19911 & n3887 ;
  assign n19912 = ~n3887 ;
  assign n3889 = n3632 & n19912 ;
  assign n3890 = n3888 | n3889 ;
  assign n19913 = ~n3890 ;
  assign n3891 = n3885 & n19913 ;
  assign n3892 = n3884 | n3891 ;
  assign n3893 = x75 & n3892 ;
  assign n3894 = x75 | n3892 ;
  assign n3895 = n3635 & n19812 ;
  assign n3896 = n164 & n3895 ;
  assign n19914 = ~n3641 ;
  assign n3897 = n19914 & n3896 ;
  assign n19915 = ~n3896 ;
  assign n3898 = n3641 & n19915 ;
  assign n3899 = n3897 | n3898 ;
  assign n19916 = ~n3899 ;
  assign n3900 = n3894 & n19916 ;
  assign n3901 = n3893 | n3900 ;
  assign n3902 = x76 & n3901 ;
  assign n3903 = x76 | n3901 ;
  assign n3904 = n3644 & n19816 ;
  assign n3905 = n164 & n3904 ;
  assign n19917 = ~n3650 ;
  assign n3906 = n19917 & n3905 ;
  assign n19918 = ~n3905 ;
  assign n3907 = n3650 & n19918 ;
  assign n3908 = n3906 | n3907 ;
  assign n19919 = ~n3908 ;
  assign n3909 = n3903 & n19919 ;
  assign n3910 = n3902 | n3909 ;
  assign n3911 = x77 & n3910 ;
  assign n3912 = x77 | n3910 ;
  assign n3913 = n3653 & n19820 ;
  assign n3914 = n164 & n3913 ;
  assign n19920 = ~n3659 ;
  assign n3915 = n19920 & n3914 ;
  assign n19921 = ~n3914 ;
  assign n3916 = n3659 & n19921 ;
  assign n3917 = n3915 | n3916 ;
  assign n19922 = ~n3917 ;
  assign n3918 = n3912 & n19922 ;
  assign n3919 = n3911 | n3918 ;
  assign n3920 = x78 & n3919 ;
  assign n3921 = x78 | n3919 ;
  assign n3922 = n3662 & n19824 ;
  assign n3923 = n164 & n3922 ;
  assign n3924 = n3668 & n3923 ;
  assign n3925 = n3668 | n3923 ;
  assign n19923 = ~n3924 ;
  assign n3926 = n19923 & n3925 ;
  assign n19924 = ~n3926 ;
  assign n3927 = n3921 & n19924 ;
  assign n3928 = n3920 | n3927 ;
  assign n3929 = x79 & n3928 ;
  assign n3930 = x79 | n3928 ;
  assign n3931 = n3671 & n19828 ;
  assign n3932 = n164 & n3931 ;
  assign n3933 = n3677 & n3932 ;
  assign n3934 = n3677 | n3932 ;
  assign n19925 = ~n3933 ;
  assign n3935 = n19925 & n3934 ;
  assign n19926 = ~n3935 ;
  assign n3936 = n3930 & n19926 ;
  assign n3937 = n3929 | n3936 ;
  assign n3938 = x80 & n3937 ;
  assign n3939 = x80 | n3937 ;
  assign n3940 = n3680 & n19832 ;
  assign n3941 = n164 & n3940 ;
  assign n3942 = n3686 & n3941 ;
  assign n3943 = n3686 | n3941 ;
  assign n19927 = ~n3942 ;
  assign n3944 = n19927 & n3943 ;
  assign n19928 = ~n3944 ;
  assign n3945 = n3939 & n19928 ;
  assign n3946 = n3938 | n3945 ;
  assign n3947 = x81 & n3946 ;
  assign n3948 = x81 | n3946 ;
  assign n3949 = n3689 & n19836 ;
  assign n3950 = n164 & n3949 ;
  assign n3951 = n3695 & n3950 ;
  assign n3952 = n3695 | n3950 ;
  assign n19929 = ~n3951 ;
  assign n3953 = n19929 & n3952 ;
  assign n19930 = ~n3953 ;
  assign n3954 = n3948 & n19930 ;
  assign n3955 = n3947 | n3954 ;
  assign n3956 = x82 & n3955 ;
  assign n3957 = x82 | n3955 ;
  assign n3958 = n3698 & n19840 ;
  assign n3959 = n164 & n3958 ;
  assign n3960 = n3704 & n3959 ;
  assign n3961 = n3704 | n3959 ;
  assign n19931 = ~n3960 ;
  assign n3962 = n19931 & n3961 ;
  assign n19932 = ~n3962 ;
  assign n3963 = n3957 & n19932 ;
  assign n3964 = n3956 | n3963 ;
  assign n3965 = x83 & n3964 ;
  assign n3966 = x83 | n3964 ;
  assign n3967 = n3707 & n19844 ;
  assign n3968 = n164 & n3967 ;
  assign n3969 = n3713 & n3968 ;
  assign n3970 = n3713 | n3968 ;
  assign n19933 = ~n3969 ;
  assign n3971 = n19933 & n3970 ;
  assign n19934 = ~n3971 ;
  assign n3972 = n3966 & n19934 ;
  assign n3973 = n3965 | n3972 ;
  assign n3974 = x84 & n3973 ;
  assign n3975 = x84 | n3973 ;
  assign n3976 = n3716 & n19848 ;
  assign n3977 = n164 & n3976 ;
  assign n3978 = n3722 & n3977 ;
  assign n3979 = n3722 | n3977 ;
  assign n19935 = ~n3978 ;
  assign n3980 = n19935 & n3979 ;
  assign n19936 = ~n3980 ;
  assign n3981 = n3975 & n19936 ;
  assign n3982 = n3974 | n3981 ;
  assign n3983 = x85 & n3982 ;
  assign n3984 = x85 | n3982 ;
  assign n3985 = n3725 & n19852 ;
  assign n3986 = n164 & n3985 ;
  assign n3987 = n3731 & n3986 ;
  assign n3988 = n3731 | n3986 ;
  assign n19937 = ~n3987 ;
  assign n3989 = n19937 & n3988 ;
  assign n19938 = ~n3989 ;
  assign n3990 = n3984 & n19938 ;
  assign n3991 = n3983 | n3990 ;
  assign n3992 = x86 & n3991 ;
  assign n3993 = x86 | n3991 ;
  assign n3994 = n3734 & n19856 ;
  assign n3995 = n164 & n3994 ;
  assign n3996 = n3740 & n3995 ;
  assign n3997 = n3740 | n3995 ;
  assign n19939 = ~n3996 ;
  assign n3998 = n19939 & n3997 ;
  assign n19940 = ~n3998 ;
  assign n3999 = n3993 & n19940 ;
  assign n4000 = n3992 | n3999 ;
  assign n4001 = x87 & n4000 ;
  assign n4002 = x87 | n4000 ;
  assign n4003 = n3743 & n19860 ;
  assign n4004 = n164 & n4003 ;
  assign n4005 = n3749 & n4004 ;
  assign n4006 = n3749 | n4004 ;
  assign n19941 = ~n4005 ;
  assign n4007 = n19941 & n4006 ;
  assign n19942 = ~n4007 ;
  assign n4008 = n4002 & n19942 ;
  assign n4009 = n4001 | n4008 ;
  assign n4010 = x88 & n4009 ;
  assign n4011 = x88 | n4009 ;
  assign n4012 = n3752 & n19864 ;
  assign n4013 = n164 & n4012 ;
  assign n4014 = n3758 & n4013 ;
  assign n4015 = n3758 | n4013 ;
  assign n19943 = ~n4014 ;
  assign n4016 = n19943 & n4015 ;
  assign n19944 = ~n4016 ;
  assign n4017 = n4011 & n19944 ;
  assign n4018 = n4010 | n4017 ;
  assign n4019 = x89 & n4018 ;
  assign n4020 = x89 | n4018 ;
  assign n4021 = n3761 & n19868 ;
  assign n4022 = n164 & n4021 ;
  assign n4023 = n3767 & n4022 ;
  assign n4024 = n3767 | n4022 ;
  assign n19945 = ~n4023 ;
  assign n4025 = n19945 & n4024 ;
  assign n19946 = ~n4025 ;
  assign n4026 = n4020 & n19946 ;
  assign n4027 = n4019 | n4026 ;
  assign n4028 = x90 & n4027 ;
  assign n4029 = x90 | n4027 ;
  assign n4030 = n3770 & n19872 ;
  assign n4031 = n164 & n4030 ;
  assign n4032 = n3776 & n4031 ;
  assign n4033 = n3776 | n4031 ;
  assign n19947 = ~n4032 ;
  assign n4034 = n19947 & n4033 ;
  assign n19948 = ~n4034 ;
  assign n4035 = n4029 & n19948 ;
  assign n4036 = n4028 | n4035 ;
  assign n4037 = x91 & n4036 ;
  assign n4038 = x91 | n4036 ;
  assign n4039 = n3779 & n19876 ;
  assign n4040 = n164 & n4039 ;
  assign n4041 = n3785 & n4040 ;
  assign n4042 = n3785 | n4040 ;
  assign n19949 = ~n4041 ;
  assign n4043 = n19949 & n4042 ;
  assign n19950 = ~n4043 ;
  assign n4044 = n4038 & n19950 ;
  assign n4045 = n4037 | n4044 ;
  assign n4046 = x92 & n4045 ;
  assign n19951 = ~n4046 ;
  assign n4047 = n3802 & n19951 ;
  assign n4048 = x92 | n4045 ;
  assign n19952 = ~n4047 ;
  assign n4049 = n19952 & n4048 ;
  assign n4051 = x93 & n4049 ;
  assign n4052 = n18428 | n4051 ;
  assign n4050 = x93 | n4049 ;
  assign n4053 = n3545 & n3795 ;
  assign n4054 = n21884 | n4053 ;
  assign n19953 = ~n4054 ;
  assign n4055 = n4050 & n19953 ;
  assign n4056 = n4052 | n4055 ;
  assign n163 = ~n4056 ;
  assign n4058 = n4048 & n163 ;
  assign n4059 = n4047 & n4058 ;
  assign n4060 = n19951 & n4058 ;
  assign n4061 = n3802 | n4060 ;
  assign n19955 = ~n4059 ;
  assign n4062 = n19955 & n4061 ;
  assign n19956 = ~x33 ;
  assign n4066 = n19956 & x64 ;
  assign n4067 = x65 | n4066 ;
  assign n4057 = n3803 & n163 ;
  assign n4068 = x64 & n163 ;
  assign n19957 = ~n4068 ;
  assign n4069 = x34 & n19957 ;
  assign n4070 = n4057 | n4069 ;
  assign n4071 = x65 & n4066 ;
  assign n19958 = ~n4071 ;
  assign n4072 = n4070 & n19958 ;
  assign n19959 = ~n4072 ;
  assign n4073 = n4067 & n19959 ;
  assign n4074 = x66 & n4073 ;
  assign n4075 = n19887 & n3805 ;
  assign n4076 = n163 & n4075 ;
  assign n4077 = n3809 & n4076 ;
  assign n4078 = n3809 | n4076 ;
  assign n19960 = ~n4077 ;
  assign n4079 = n19960 & n4078 ;
  assign n4080 = x66 | n4073 ;
  assign n19961 = ~n4079 ;
  assign n4081 = n19961 & n4080 ;
  assign n4082 = n4074 | n4081 ;
  assign n4083 = x67 & n4082 ;
  assign n4084 = x67 | n4082 ;
  assign n19962 = ~n3812 ;
  assign n4085 = n19962 & n3813 ;
  assign n4086 = n163 & n4085 ;
  assign n4087 = n3818 & n4086 ;
  assign n4088 = n3818 | n4086 ;
  assign n19963 = ~n4087 ;
  assign n4089 = n19963 & n4088 ;
  assign n19964 = ~n4089 ;
  assign n4090 = n4084 & n19964 ;
  assign n4091 = n4083 | n4090 ;
  assign n4092 = x68 & n4091 ;
  assign n4093 = x68 | n4091 ;
  assign n19965 = ~n3821 ;
  assign n4094 = n19965 & n3822 ;
  assign n4095 = n163 & n4094 ;
  assign n4096 = n3827 & n4095 ;
  assign n4097 = n3827 | n4095 ;
  assign n19966 = ~n4096 ;
  assign n4098 = n19966 & n4097 ;
  assign n19967 = ~n4098 ;
  assign n4099 = n4093 & n19967 ;
  assign n4100 = n4092 | n4099 ;
  assign n4101 = x69 & n4100 ;
  assign n4102 = x69 | n4100 ;
  assign n19968 = ~n3830 ;
  assign n4103 = n19968 & n3831 ;
  assign n4104 = n163 & n4103 ;
  assign n4105 = n3836 & n4104 ;
  assign n4106 = n3836 | n4104 ;
  assign n19969 = ~n4105 ;
  assign n4107 = n19969 & n4106 ;
  assign n19970 = ~n4107 ;
  assign n4108 = n4102 & n19970 ;
  assign n4109 = n4101 | n4108 ;
  assign n4110 = x70 & n4109 ;
  assign n4111 = x70 | n4109 ;
  assign n19971 = ~n3839 ;
  assign n4112 = n19971 & n3840 ;
  assign n4113 = n163 & n4112 ;
  assign n4114 = n3845 & n4113 ;
  assign n4115 = n3845 | n4113 ;
  assign n19972 = ~n4114 ;
  assign n4116 = n19972 & n4115 ;
  assign n19973 = ~n4116 ;
  assign n4117 = n4111 & n19973 ;
  assign n4118 = n4110 | n4117 ;
  assign n4119 = x71 & n4118 ;
  assign n4120 = x71 | n4118 ;
  assign n19974 = ~n3848 ;
  assign n4121 = n19974 & n3849 ;
  assign n4122 = n163 & n4121 ;
  assign n4123 = n3854 & n4122 ;
  assign n4124 = n3854 | n4122 ;
  assign n19975 = ~n4123 ;
  assign n4125 = n19975 & n4124 ;
  assign n19976 = ~n4125 ;
  assign n4126 = n4120 & n19976 ;
  assign n4127 = n4119 | n4126 ;
  assign n4128 = x72 & n4127 ;
  assign n4129 = x72 | n4127 ;
  assign n19977 = ~n3857 ;
  assign n4130 = n19977 & n3858 ;
  assign n4131 = n163 & n4130 ;
  assign n4132 = n3863 & n4131 ;
  assign n4133 = n3863 | n4131 ;
  assign n19978 = ~n4132 ;
  assign n4134 = n19978 & n4133 ;
  assign n19979 = ~n4134 ;
  assign n4135 = n4129 & n19979 ;
  assign n4136 = n4128 | n4135 ;
  assign n4137 = x73 & n4136 ;
  assign n4138 = x73 | n4136 ;
  assign n19980 = ~n3866 ;
  assign n4139 = n19980 & n3867 ;
  assign n4140 = n163 & n4139 ;
  assign n4141 = n19907 & n4140 ;
  assign n19981 = ~n4140 ;
  assign n4142 = n3872 & n19981 ;
  assign n4143 = n4141 | n4142 ;
  assign n19982 = ~n4143 ;
  assign n4144 = n4138 & n19982 ;
  assign n4145 = n4137 | n4144 ;
  assign n4146 = x74 & n4145 ;
  assign n4147 = x74 | n4145 ;
  assign n19983 = ~n3875 ;
  assign n4148 = n19983 & n3876 ;
  assign n4149 = n163 & n4148 ;
  assign n4150 = n19910 & n4149 ;
  assign n19984 = ~n4149 ;
  assign n4151 = n3881 & n19984 ;
  assign n4152 = n4150 | n4151 ;
  assign n19985 = ~n4152 ;
  assign n4153 = n4147 & n19985 ;
  assign n4154 = n4146 | n4153 ;
  assign n4155 = x75 & n4154 ;
  assign n4156 = x75 | n4154 ;
  assign n19986 = ~n3884 ;
  assign n4157 = n19986 & n3885 ;
  assign n4158 = n163 & n4157 ;
  assign n4159 = n19913 & n4158 ;
  assign n19987 = ~n4158 ;
  assign n4160 = n3890 & n19987 ;
  assign n4161 = n4159 | n4160 ;
  assign n19988 = ~n4161 ;
  assign n4162 = n4156 & n19988 ;
  assign n4163 = n4155 | n4162 ;
  assign n4164 = x76 & n4163 ;
  assign n4165 = x76 | n4163 ;
  assign n19989 = ~n3893 ;
  assign n4166 = n19989 & n3894 ;
  assign n4167 = n163 & n4166 ;
  assign n4168 = n19916 & n4167 ;
  assign n19990 = ~n4167 ;
  assign n4169 = n3899 & n19990 ;
  assign n4170 = n4168 | n4169 ;
  assign n19991 = ~n4170 ;
  assign n4171 = n4165 & n19991 ;
  assign n4172 = n4164 | n4171 ;
  assign n4173 = x77 & n4172 ;
  assign n4174 = x77 | n4172 ;
  assign n19992 = ~n3902 ;
  assign n4175 = n19992 & n3903 ;
  assign n4176 = n163 & n4175 ;
  assign n4177 = n3908 & n4176 ;
  assign n4178 = n3908 | n4176 ;
  assign n19993 = ~n4177 ;
  assign n4179 = n19993 & n4178 ;
  assign n19994 = ~n4179 ;
  assign n4180 = n4174 & n19994 ;
  assign n4181 = n4173 | n4180 ;
  assign n4182 = x78 & n4181 ;
  assign n4183 = x78 | n4181 ;
  assign n19995 = ~n3911 ;
  assign n4184 = n19995 & n3912 ;
  assign n4185 = n163 & n4184 ;
  assign n4186 = n3917 & n4185 ;
  assign n4187 = n3917 | n4185 ;
  assign n19996 = ~n4186 ;
  assign n4188 = n19996 & n4187 ;
  assign n19997 = ~n4188 ;
  assign n4189 = n4183 & n19997 ;
  assign n4190 = n4182 | n4189 ;
  assign n4191 = x79 & n4190 ;
  assign n4192 = x79 | n4190 ;
  assign n19998 = ~n3920 ;
  assign n4193 = n19998 & n3921 ;
  assign n4194 = n163 & n4193 ;
  assign n4195 = n3926 & n4194 ;
  assign n4196 = n3926 | n4194 ;
  assign n19999 = ~n4195 ;
  assign n4197 = n19999 & n4196 ;
  assign n20000 = ~n4197 ;
  assign n4198 = n4192 & n20000 ;
  assign n4199 = n4191 | n4198 ;
  assign n4200 = x80 & n4199 ;
  assign n4201 = x80 | n4199 ;
  assign n20001 = ~n3929 ;
  assign n4202 = n20001 & n3930 ;
  assign n4203 = n163 & n4202 ;
  assign n4204 = n3935 & n4203 ;
  assign n4205 = n3935 | n4203 ;
  assign n20002 = ~n4204 ;
  assign n4206 = n20002 & n4205 ;
  assign n20003 = ~n4206 ;
  assign n4207 = n4201 & n20003 ;
  assign n4208 = n4200 | n4207 ;
  assign n4209 = x81 & n4208 ;
  assign n4210 = x81 | n4208 ;
  assign n20004 = ~n3938 ;
  assign n4211 = n20004 & n3939 ;
  assign n4212 = n163 & n4211 ;
  assign n4213 = n3944 & n4212 ;
  assign n4214 = n3944 | n4212 ;
  assign n20005 = ~n4213 ;
  assign n4215 = n20005 & n4214 ;
  assign n20006 = ~n4215 ;
  assign n4216 = n4210 & n20006 ;
  assign n4217 = n4209 | n4216 ;
  assign n4218 = x82 & n4217 ;
  assign n4219 = x82 | n4217 ;
  assign n20007 = ~n3947 ;
  assign n4220 = n20007 & n3948 ;
  assign n4221 = n163 & n4220 ;
  assign n4222 = n3953 & n4221 ;
  assign n4223 = n3953 | n4221 ;
  assign n20008 = ~n4222 ;
  assign n4224 = n20008 & n4223 ;
  assign n20009 = ~n4224 ;
  assign n4225 = n4219 & n20009 ;
  assign n4226 = n4218 | n4225 ;
  assign n4227 = x83 & n4226 ;
  assign n4228 = x83 | n4226 ;
  assign n20010 = ~n3956 ;
  assign n4229 = n20010 & n3957 ;
  assign n4230 = n163 & n4229 ;
  assign n4231 = n3962 & n4230 ;
  assign n4232 = n3962 | n4230 ;
  assign n20011 = ~n4231 ;
  assign n4233 = n20011 & n4232 ;
  assign n20012 = ~n4233 ;
  assign n4234 = n4228 & n20012 ;
  assign n4235 = n4227 | n4234 ;
  assign n4236 = x84 & n4235 ;
  assign n4237 = x84 | n4235 ;
  assign n20013 = ~n3965 ;
  assign n4238 = n20013 & n3966 ;
  assign n4239 = n163 & n4238 ;
  assign n4240 = n3971 & n4239 ;
  assign n4241 = n3971 | n4239 ;
  assign n20014 = ~n4240 ;
  assign n4242 = n20014 & n4241 ;
  assign n20015 = ~n4242 ;
  assign n4243 = n4237 & n20015 ;
  assign n4244 = n4236 | n4243 ;
  assign n4245 = x85 & n4244 ;
  assign n4246 = x85 | n4244 ;
  assign n20016 = ~n3974 ;
  assign n4247 = n20016 & n3975 ;
  assign n4248 = n163 & n4247 ;
  assign n4249 = n3980 & n4248 ;
  assign n4250 = n3980 | n4248 ;
  assign n20017 = ~n4249 ;
  assign n4251 = n20017 & n4250 ;
  assign n20018 = ~n4251 ;
  assign n4252 = n4246 & n20018 ;
  assign n4253 = n4245 | n4252 ;
  assign n4254 = x86 & n4253 ;
  assign n4255 = x86 | n4253 ;
  assign n20019 = ~n3983 ;
  assign n4256 = n20019 & n3984 ;
  assign n4257 = n163 & n4256 ;
  assign n4258 = n3989 & n4257 ;
  assign n4259 = n3989 | n4257 ;
  assign n20020 = ~n4258 ;
  assign n4260 = n20020 & n4259 ;
  assign n20021 = ~n4260 ;
  assign n4261 = n4255 & n20021 ;
  assign n4262 = n4254 | n4261 ;
  assign n4263 = x87 & n4262 ;
  assign n4264 = x87 | n4262 ;
  assign n20022 = ~n3992 ;
  assign n4265 = n20022 & n3993 ;
  assign n4266 = n163 & n4265 ;
  assign n4267 = n3998 & n4266 ;
  assign n4268 = n3998 | n4266 ;
  assign n20023 = ~n4267 ;
  assign n4269 = n20023 & n4268 ;
  assign n20024 = ~n4269 ;
  assign n4270 = n4264 & n20024 ;
  assign n4271 = n4263 | n4270 ;
  assign n4272 = x88 & n4271 ;
  assign n4273 = x88 | n4271 ;
  assign n20025 = ~n4001 ;
  assign n4274 = n20025 & n4002 ;
  assign n4275 = n163 & n4274 ;
  assign n4276 = n4007 & n4275 ;
  assign n4277 = n4007 | n4275 ;
  assign n20026 = ~n4276 ;
  assign n4278 = n20026 & n4277 ;
  assign n20027 = ~n4278 ;
  assign n4279 = n4273 & n20027 ;
  assign n4280 = n4272 | n4279 ;
  assign n4281 = x89 & n4280 ;
  assign n4282 = x89 | n4280 ;
  assign n20028 = ~n4010 ;
  assign n4283 = n20028 & n4011 ;
  assign n4284 = n163 & n4283 ;
  assign n4285 = n4016 & n4284 ;
  assign n4286 = n4016 | n4284 ;
  assign n20029 = ~n4285 ;
  assign n4287 = n20029 & n4286 ;
  assign n20030 = ~n4287 ;
  assign n4288 = n4282 & n20030 ;
  assign n4289 = n4281 | n4288 ;
  assign n4290 = x90 & n4289 ;
  assign n4291 = x90 | n4289 ;
  assign n20031 = ~n4019 ;
  assign n4292 = n20031 & n4020 ;
  assign n4293 = n163 & n4292 ;
  assign n4294 = n4025 & n4293 ;
  assign n4295 = n4025 | n4293 ;
  assign n20032 = ~n4294 ;
  assign n4296 = n20032 & n4295 ;
  assign n20033 = ~n4296 ;
  assign n4297 = n4291 & n20033 ;
  assign n4298 = n4290 | n4297 ;
  assign n4299 = x91 & n4298 ;
  assign n4300 = x91 | n4298 ;
  assign n20034 = ~n4028 ;
  assign n4301 = n20034 & n4029 ;
  assign n4302 = n163 & n4301 ;
  assign n4303 = n4034 & n4302 ;
  assign n4304 = n4034 | n4302 ;
  assign n20035 = ~n4303 ;
  assign n4305 = n20035 & n4304 ;
  assign n20036 = ~n4305 ;
  assign n4306 = n4300 & n20036 ;
  assign n4307 = n4299 | n4306 ;
  assign n4308 = x92 & n4307 ;
  assign n4309 = x92 | n4307 ;
  assign n20037 = ~n4037 ;
  assign n4310 = n20037 & n4038 ;
  assign n4311 = n163 & n4310 ;
  assign n4312 = n4043 & n4311 ;
  assign n4313 = n4043 | n4311 ;
  assign n20038 = ~n4312 ;
  assign n4314 = n20038 & n4313 ;
  assign n20039 = ~n4314 ;
  assign n4315 = n4309 & n20039 ;
  assign n4316 = n4308 | n4315 ;
  assign n4318 = x93 & n4316 ;
  assign n20040 = ~n4318 ;
  assign n4319 = n4062 & n20040 ;
  assign n4063 = n21884 | n4052 ;
  assign n4064 = n4054 & n4063 ;
  assign n20041 = ~x94 ;
  assign n4065 = n20041 & n4064 ;
  assign n4317 = x93 | n4316 ;
  assign n20042 = ~n4065 ;
  assign n4320 = n20042 & n4317 ;
  assign n20043 = ~n4319 ;
  assign n4321 = n20043 & n4320 ;
  assign n4322 = n18423 | n4321 ;
  assign n20044 = ~n4064 ;
  assign n4324 = x94 & n20044 ;
  assign n4325 = n4322 | n4324 ;
  assign n4326 = n4317 & n20040 ;
  assign n162 = ~n4325 ;
  assign n4327 = n162 & n4326 ;
  assign n4328 = n4062 & n4327 ;
  assign n4329 = n4062 | n4327 ;
  assign n20046 = ~n4328 ;
  assign n4330 = n20046 & n4329 ;
  assign n4323 = n21884 | n4322 ;
  assign n4331 = n4064 & n4323 ;
  assign n20047 = ~n18418 ;
  assign n4334 = n20047 & n4331 ;
  assign n20048 = ~n4334 ;
  assign n4601 = n18423 & n20048 ;
  assign n20049 = ~x32 ;
  assign n4335 = n20049 & x64 ;
  assign n4337 = x65 | n4335 ;
  assign n4336 = x65 & n4335 ;
  assign n4338 = x64 & n162 ;
  assign n4339 = x33 & n4338 ;
  assign n4340 = x33 | n4338 ;
  assign n20050 = ~n4339 ;
  assign n4341 = n20050 & n4340 ;
  assign n20051 = ~n4336 ;
  assign n4342 = n20051 & n4341 ;
  assign n20052 = ~n4342 ;
  assign n4343 = n4337 & n20052 ;
  assign n4344 = x66 | n4343 ;
  assign n4345 = x66 & n4343 ;
  assign n4346 = n4067 & n162 ;
  assign n4347 = n19958 & n4346 ;
  assign n4348 = n4070 | n4347 ;
  assign n4349 = n4072 & n4346 ;
  assign n20053 = ~n4349 ;
  assign n4350 = n4348 & n20053 ;
  assign n20054 = ~n4345 ;
  assign n4351 = n20054 & n4350 ;
  assign n20055 = ~n4351 ;
  assign n4352 = n4344 & n20055 ;
  assign n4353 = x67 | n4352 ;
  assign n4354 = x67 & n4352 ;
  assign n20056 = ~n4074 ;
  assign n4355 = n20056 & n4080 ;
  assign n4356 = n162 & n4355 ;
  assign n4357 = n4079 & n4356 ;
  assign n4358 = n4079 | n4356 ;
  assign n20057 = ~n4357 ;
  assign n4359 = n20057 & n4358 ;
  assign n20058 = ~n4354 ;
  assign n4360 = n20058 & n4359 ;
  assign n20059 = ~n4360 ;
  assign n4361 = n4353 & n20059 ;
  assign n4362 = x68 | n4361 ;
  assign n4363 = x68 & n4361 ;
  assign n20060 = ~n4083 ;
  assign n4364 = n20060 & n4084 ;
  assign n4365 = n162 & n4364 ;
  assign n4366 = n4089 & n4365 ;
  assign n4367 = n4089 | n4365 ;
  assign n20061 = ~n4366 ;
  assign n4368 = n20061 & n4367 ;
  assign n20062 = ~n4363 ;
  assign n4369 = n20062 & n4368 ;
  assign n20063 = ~n4369 ;
  assign n4370 = n4362 & n20063 ;
  assign n4371 = x69 | n4370 ;
  assign n4372 = x69 & n4370 ;
  assign n20064 = ~n4092 ;
  assign n4373 = n20064 & n4093 ;
  assign n4374 = n162 & n4373 ;
  assign n4375 = n19967 & n4374 ;
  assign n20065 = ~n4374 ;
  assign n4376 = n4098 & n20065 ;
  assign n4377 = n4375 | n4376 ;
  assign n20066 = ~n4372 ;
  assign n4378 = n20066 & n4377 ;
  assign n20067 = ~n4378 ;
  assign n4379 = n4371 & n20067 ;
  assign n4380 = x70 | n4379 ;
  assign n4381 = x70 & n4379 ;
  assign n20068 = ~n4101 ;
  assign n4382 = n20068 & n4102 ;
  assign n4383 = n162 & n4382 ;
  assign n4384 = n4107 & n4383 ;
  assign n4385 = n4107 | n4383 ;
  assign n20069 = ~n4384 ;
  assign n4386 = n20069 & n4385 ;
  assign n20070 = ~n4381 ;
  assign n4387 = n20070 & n4386 ;
  assign n20071 = ~n4387 ;
  assign n4388 = n4380 & n20071 ;
  assign n4389 = x71 | n4388 ;
  assign n4390 = x71 & n4388 ;
  assign n20072 = ~n4110 ;
  assign n4391 = n20072 & n4111 ;
  assign n4392 = n162 & n4391 ;
  assign n4393 = n4116 & n4392 ;
  assign n4394 = n4116 | n4392 ;
  assign n20073 = ~n4393 ;
  assign n4395 = n20073 & n4394 ;
  assign n20074 = ~n4390 ;
  assign n4396 = n20074 & n4395 ;
  assign n20075 = ~n4396 ;
  assign n4397 = n4389 & n20075 ;
  assign n4398 = x72 | n4397 ;
  assign n4399 = x72 & n4397 ;
  assign n20076 = ~n4119 ;
  assign n4400 = n20076 & n4120 ;
  assign n4401 = n162 & n4400 ;
  assign n4402 = n4125 & n4401 ;
  assign n4403 = n4125 | n4401 ;
  assign n20077 = ~n4402 ;
  assign n4404 = n20077 & n4403 ;
  assign n20078 = ~n4399 ;
  assign n4405 = n20078 & n4404 ;
  assign n20079 = ~n4405 ;
  assign n4406 = n4398 & n20079 ;
  assign n4407 = x73 | n4406 ;
  assign n4408 = x73 & n4406 ;
  assign n20080 = ~n4128 ;
  assign n4409 = n20080 & n4129 ;
  assign n4410 = n162 & n4409 ;
  assign n4411 = n4134 & n4410 ;
  assign n4412 = n4134 | n4410 ;
  assign n20081 = ~n4411 ;
  assign n4413 = n20081 & n4412 ;
  assign n20082 = ~n4408 ;
  assign n4414 = n20082 & n4413 ;
  assign n20083 = ~n4414 ;
  assign n4415 = n4407 & n20083 ;
  assign n4416 = x74 | n4415 ;
  assign n4417 = x74 & n4415 ;
  assign n20084 = ~n4137 ;
  assign n4418 = n20084 & n4138 ;
  assign n4419 = n162 & n4418 ;
  assign n4420 = n19982 & n4419 ;
  assign n20085 = ~n4419 ;
  assign n4421 = n4143 & n20085 ;
  assign n4422 = n4420 | n4421 ;
  assign n20086 = ~n4417 ;
  assign n4423 = n20086 & n4422 ;
  assign n20087 = ~n4423 ;
  assign n4424 = n4416 & n20087 ;
  assign n4425 = x75 | n4424 ;
  assign n4426 = x75 & n4424 ;
  assign n20088 = ~n4146 ;
  assign n4427 = n20088 & n4147 ;
  assign n4428 = n162 & n4427 ;
  assign n4429 = n19985 & n4428 ;
  assign n20089 = ~n4428 ;
  assign n4430 = n4152 & n20089 ;
  assign n4431 = n4429 | n4430 ;
  assign n20090 = ~n4426 ;
  assign n4432 = n20090 & n4431 ;
  assign n20091 = ~n4432 ;
  assign n4433 = n4425 & n20091 ;
  assign n4434 = x76 | n4433 ;
  assign n4435 = x76 & n4433 ;
  assign n20092 = ~n4155 ;
  assign n4436 = n20092 & n4156 ;
  assign n4437 = n162 & n4436 ;
  assign n4438 = n19988 & n4437 ;
  assign n20093 = ~n4437 ;
  assign n4439 = n4161 & n20093 ;
  assign n4440 = n4438 | n4439 ;
  assign n20094 = ~n4435 ;
  assign n4441 = n20094 & n4440 ;
  assign n20095 = ~n4441 ;
  assign n4442 = n4434 & n20095 ;
  assign n4443 = x77 | n4442 ;
  assign n4444 = x77 & n4442 ;
  assign n20096 = ~n4164 ;
  assign n4445 = n20096 & n4165 ;
  assign n4446 = n162 & n4445 ;
  assign n4447 = n4170 & n4446 ;
  assign n4448 = n4170 | n4446 ;
  assign n20097 = ~n4447 ;
  assign n4449 = n20097 & n4448 ;
  assign n20098 = ~n4444 ;
  assign n4450 = n20098 & n4449 ;
  assign n20099 = ~n4450 ;
  assign n4451 = n4443 & n20099 ;
  assign n4452 = x78 | n4451 ;
  assign n4453 = x78 & n4451 ;
  assign n20100 = ~n4173 ;
  assign n4454 = n20100 & n4174 ;
  assign n4455 = n162 & n4454 ;
  assign n4456 = n4179 & n4455 ;
  assign n4457 = n4179 | n4455 ;
  assign n20101 = ~n4456 ;
  assign n4458 = n20101 & n4457 ;
  assign n20102 = ~n4453 ;
  assign n4459 = n20102 & n4458 ;
  assign n20103 = ~n4459 ;
  assign n4460 = n4452 & n20103 ;
  assign n4461 = x79 | n4460 ;
  assign n4462 = x79 & n4460 ;
  assign n20104 = ~n4182 ;
  assign n4463 = n20104 & n4183 ;
  assign n4464 = n162 & n4463 ;
  assign n4465 = n4188 & n4464 ;
  assign n4466 = n4188 | n4464 ;
  assign n20105 = ~n4465 ;
  assign n4467 = n20105 & n4466 ;
  assign n20106 = ~n4462 ;
  assign n4468 = n20106 & n4467 ;
  assign n20107 = ~n4468 ;
  assign n4469 = n4461 & n20107 ;
  assign n4470 = x80 | n4469 ;
  assign n4471 = x80 & n4469 ;
  assign n20108 = ~n4191 ;
  assign n4472 = n20108 & n4192 ;
  assign n4473 = n162 & n4472 ;
  assign n4474 = n20000 & n4473 ;
  assign n20109 = ~n4473 ;
  assign n4475 = n4197 & n20109 ;
  assign n4476 = n4474 | n4475 ;
  assign n20110 = ~n4471 ;
  assign n4477 = n20110 & n4476 ;
  assign n20111 = ~n4477 ;
  assign n4478 = n4470 & n20111 ;
  assign n4479 = x81 | n4478 ;
  assign n4480 = x81 & n4478 ;
  assign n20112 = ~n4200 ;
  assign n4481 = n20112 & n4201 ;
  assign n4482 = n162 & n4481 ;
  assign n4483 = n20003 & n4482 ;
  assign n20113 = ~n4482 ;
  assign n4484 = n4206 & n20113 ;
  assign n4485 = n4483 | n4484 ;
  assign n20114 = ~n4480 ;
  assign n4486 = n20114 & n4485 ;
  assign n20115 = ~n4486 ;
  assign n4487 = n4479 & n20115 ;
  assign n4488 = x82 | n4487 ;
  assign n4489 = x82 & n4487 ;
  assign n20116 = ~n4209 ;
  assign n4490 = n20116 & n4210 ;
  assign n4491 = n162 & n4490 ;
  assign n4492 = n20006 & n4491 ;
  assign n20117 = ~n4491 ;
  assign n4493 = n4215 & n20117 ;
  assign n4494 = n4492 | n4493 ;
  assign n20118 = ~n4489 ;
  assign n4495 = n20118 & n4494 ;
  assign n20119 = ~n4495 ;
  assign n4496 = n4488 & n20119 ;
  assign n4497 = x83 | n4496 ;
  assign n4498 = x83 & n4496 ;
  assign n20120 = ~n4218 ;
  assign n4499 = n20120 & n4219 ;
  assign n4500 = n162 & n4499 ;
  assign n4501 = n20009 & n4500 ;
  assign n20121 = ~n4500 ;
  assign n4502 = n4224 & n20121 ;
  assign n4503 = n4501 | n4502 ;
  assign n20122 = ~n4498 ;
  assign n4504 = n20122 & n4503 ;
  assign n20123 = ~n4504 ;
  assign n4505 = n4497 & n20123 ;
  assign n4506 = x84 | n4505 ;
  assign n4507 = x84 & n4505 ;
  assign n20124 = ~n4227 ;
  assign n4508 = n20124 & n4228 ;
  assign n4509 = n162 & n4508 ;
  assign n4510 = n20012 & n4509 ;
  assign n20125 = ~n4509 ;
  assign n4511 = n4233 & n20125 ;
  assign n4512 = n4510 | n4511 ;
  assign n20126 = ~n4507 ;
  assign n4513 = n20126 & n4512 ;
  assign n20127 = ~n4513 ;
  assign n4514 = n4506 & n20127 ;
  assign n4515 = x85 | n4514 ;
  assign n4516 = x85 & n4514 ;
  assign n20128 = ~n4236 ;
  assign n4517 = n20128 & n4237 ;
  assign n4518 = n162 & n4517 ;
  assign n4519 = n20015 & n4518 ;
  assign n20129 = ~n4518 ;
  assign n4520 = n4242 & n20129 ;
  assign n4521 = n4519 | n4520 ;
  assign n20130 = ~n4516 ;
  assign n4522 = n20130 & n4521 ;
  assign n20131 = ~n4522 ;
  assign n4523 = n4515 & n20131 ;
  assign n4524 = x86 | n4523 ;
  assign n4525 = x86 & n4523 ;
  assign n20132 = ~n4245 ;
  assign n4526 = n20132 & n4246 ;
  assign n4527 = n162 & n4526 ;
  assign n4528 = n20018 & n4527 ;
  assign n20133 = ~n4527 ;
  assign n4529 = n4251 & n20133 ;
  assign n4530 = n4528 | n4529 ;
  assign n20134 = ~n4525 ;
  assign n4531 = n20134 & n4530 ;
  assign n20135 = ~n4531 ;
  assign n4532 = n4524 & n20135 ;
  assign n4533 = x87 | n4532 ;
  assign n4534 = x87 & n4532 ;
  assign n20136 = ~n4254 ;
  assign n4535 = n20136 & n4255 ;
  assign n4536 = n162 & n4535 ;
  assign n4537 = n20021 & n4536 ;
  assign n20137 = ~n4536 ;
  assign n4538 = n4260 & n20137 ;
  assign n4539 = n4537 | n4538 ;
  assign n20138 = ~n4534 ;
  assign n4540 = n20138 & n4539 ;
  assign n20139 = ~n4540 ;
  assign n4541 = n4533 & n20139 ;
  assign n4542 = x88 | n4541 ;
  assign n4543 = x88 & n4541 ;
  assign n20140 = ~n4263 ;
  assign n4544 = n20140 & n4264 ;
  assign n4545 = n162 & n4544 ;
  assign n4546 = n20024 & n4545 ;
  assign n20141 = ~n4545 ;
  assign n4547 = n4269 & n20141 ;
  assign n4548 = n4546 | n4547 ;
  assign n20142 = ~n4543 ;
  assign n4549 = n20142 & n4548 ;
  assign n20143 = ~n4549 ;
  assign n4550 = n4542 & n20143 ;
  assign n4551 = x89 | n4550 ;
  assign n4552 = x89 & n4550 ;
  assign n20144 = ~n4272 ;
  assign n4553 = n20144 & n4273 ;
  assign n4554 = n162 & n4553 ;
  assign n4555 = n20027 & n4554 ;
  assign n20145 = ~n4554 ;
  assign n4556 = n4278 & n20145 ;
  assign n4557 = n4555 | n4556 ;
  assign n20146 = ~n4552 ;
  assign n4558 = n20146 & n4557 ;
  assign n20147 = ~n4558 ;
  assign n4559 = n4551 & n20147 ;
  assign n4560 = x90 | n4559 ;
  assign n4561 = x90 & n4559 ;
  assign n20148 = ~n4281 ;
  assign n4562 = n20148 & n4282 ;
  assign n4563 = n162 & n4562 ;
  assign n4564 = n20030 & n4563 ;
  assign n20149 = ~n4563 ;
  assign n4565 = n4287 & n20149 ;
  assign n4566 = n4564 | n4565 ;
  assign n20150 = ~n4561 ;
  assign n4567 = n20150 & n4566 ;
  assign n20151 = ~n4567 ;
  assign n4568 = n4560 & n20151 ;
  assign n4569 = x91 | n4568 ;
  assign n4570 = x91 & n4568 ;
  assign n20152 = ~n4290 ;
  assign n4571 = n20152 & n4291 ;
  assign n4572 = n162 & n4571 ;
  assign n4573 = n20033 & n4572 ;
  assign n20153 = ~n4572 ;
  assign n4574 = n4296 & n20153 ;
  assign n4575 = n4573 | n4574 ;
  assign n20154 = ~n4570 ;
  assign n4576 = n20154 & n4575 ;
  assign n20155 = ~n4576 ;
  assign n4577 = n4569 & n20155 ;
  assign n4578 = x92 | n4577 ;
  assign n4579 = x92 & n4577 ;
  assign n20156 = ~n4299 ;
  assign n4580 = n20156 & n4300 ;
  assign n4581 = n162 & n4580 ;
  assign n4582 = n20036 & n4581 ;
  assign n20157 = ~n4581 ;
  assign n4583 = n4305 & n20157 ;
  assign n4584 = n4582 | n4583 ;
  assign n20158 = ~n4579 ;
  assign n4585 = n20158 & n4584 ;
  assign n20159 = ~n4585 ;
  assign n4586 = n4578 & n20159 ;
  assign n4587 = x93 | n4586 ;
  assign n4588 = x93 & n4586 ;
  assign n20160 = ~n4308 ;
  assign n4589 = n20160 & n4309 ;
  assign n4590 = n162 & n4589 ;
  assign n4591 = n20039 & n4590 ;
  assign n20161 = ~n4590 ;
  assign n4592 = n4314 & n20161 ;
  assign n4593 = n4591 | n4592 ;
  assign n20162 = ~n4588 ;
  assign n4594 = n20162 & n4593 ;
  assign n20163 = ~n4594 ;
  assign n4595 = n4587 & n20163 ;
  assign n4596 = x94 & n4595 ;
  assign n20164 = ~n4596 ;
  assign n4597 = n4330 & n20164 ;
  assign n20165 = ~x95 ;
  assign n4598 = n20165 & n4331 ;
  assign n4599 = x94 | n4595 ;
  assign n20166 = ~n4598 ;
  assign n4600 = n20166 & n4599 ;
  assign n20167 = ~n4597 ;
  assign n4602 = n20167 & n4600 ;
  assign n4603 = n4601 | n4602 ;
  assign n4604 = n20164 & n4599 ;
  assign n161 = ~n4603 ;
  assign n4605 = n161 & n4604 ;
  assign n4606 = n4330 & n4605 ;
  assign n4607 = n4330 | n4605 ;
  assign n20169 = ~n4606 ;
  assign n4608 = n20169 & n4607 ;
  assign n4609 = n21884 | n4602 ;
  assign n4610 = n4334 & n4609 ;
  assign n20170 = ~x31 ;
  assign n4611 = n20170 & x64 ;
  assign n4613 = x65 | n4611 ;
  assign n4612 = x65 & n4611 ;
  assign n4614 = x64 & n161 ;
  assign n4615 = x32 & n4614 ;
  assign n4616 = x32 | n4614 ;
  assign n20171 = ~n4615 ;
  assign n4617 = n20171 & n4616 ;
  assign n20172 = ~n4612 ;
  assign n4618 = n20172 & n4617 ;
  assign n20173 = ~n4618 ;
  assign n4619 = n4613 & n20173 ;
  assign n4620 = x66 & n4619 ;
  assign n4621 = x66 | n4619 ;
  assign n4622 = n20051 & n4337 ;
  assign n4623 = n161 & n4622 ;
  assign n4624 = n4341 & n4623 ;
  assign n4625 = n4341 | n4623 ;
  assign n20174 = ~n4624 ;
  assign n4626 = n20174 & n4625 ;
  assign n20175 = ~n4626 ;
  assign n4627 = n4621 & n20175 ;
  assign n4628 = n4620 | n4627 ;
  assign n4629 = x67 & n4628 ;
  assign n4630 = x67 | n4628 ;
  assign n4631 = n4344 & n20054 ;
  assign n4632 = n161 & n4631 ;
  assign n20176 = ~n4350 ;
  assign n4633 = n20176 & n4632 ;
  assign n20177 = ~n4632 ;
  assign n4634 = n4350 & n20177 ;
  assign n4635 = n4633 | n4634 ;
  assign n20178 = ~n4635 ;
  assign n4636 = n4630 & n20178 ;
  assign n4637 = n4629 | n4636 ;
  assign n4638 = x68 & n4637 ;
  assign n4639 = x68 | n4637 ;
  assign n4640 = n4353 & n20058 ;
  assign n4641 = n161 & n4640 ;
  assign n20179 = ~n4359 ;
  assign n4642 = n20179 & n4641 ;
  assign n20180 = ~n4641 ;
  assign n4643 = n4359 & n20180 ;
  assign n4644 = n4642 | n4643 ;
  assign n20181 = ~n4644 ;
  assign n4645 = n4639 & n20181 ;
  assign n4646 = n4638 | n4645 ;
  assign n4647 = x69 & n4646 ;
  assign n4648 = x69 | n4646 ;
  assign n4649 = n4362 & n20062 ;
  assign n4650 = n161 & n4649 ;
  assign n20182 = ~n4368 ;
  assign n4651 = n20182 & n4650 ;
  assign n20183 = ~n4650 ;
  assign n4652 = n4368 & n20183 ;
  assign n4653 = n4651 | n4652 ;
  assign n20184 = ~n4653 ;
  assign n4654 = n4648 & n20184 ;
  assign n4655 = n4647 | n4654 ;
  assign n4656 = x70 & n4655 ;
  assign n4657 = x70 | n4655 ;
  assign n4658 = n4371 & n20066 ;
  assign n4659 = n161 & n4658 ;
  assign n20185 = ~n4377 ;
  assign n4660 = n20185 & n4659 ;
  assign n20186 = ~n4659 ;
  assign n4661 = n4377 & n20186 ;
  assign n4662 = n4660 | n4661 ;
  assign n20187 = ~n4662 ;
  assign n4663 = n4657 & n20187 ;
  assign n4664 = n4656 | n4663 ;
  assign n4665 = x71 & n4664 ;
  assign n4666 = x71 | n4664 ;
  assign n4667 = n4380 & n20070 ;
  assign n4668 = n161 & n4667 ;
  assign n4669 = n4386 & n4668 ;
  assign n4670 = n4386 | n4668 ;
  assign n20188 = ~n4669 ;
  assign n4671 = n20188 & n4670 ;
  assign n20189 = ~n4671 ;
  assign n4672 = n4666 & n20189 ;
  assign n4673 = n4665 | n4672 ;
  assign n4674 = x72 & n4673 ;
  assign n4675 = x72 | n4673 ;
  assign n4676 = n4389 & n20074 ;
  assign n4677 = n161 & n4676 ;
  assign n20190 = ~n4395 ;
  assign n4678 = n20190 & n4677 ;
  assign n20191 = ~n4677 ;
  assign n4679 = n4395 & n20191 ;
  assign n4680 = n4678 | n4679 ;
  assign n20192 = ~n4680 ;
  assign n4681 = n4675 & n20192 ;
  assign n4682 = n4674 | n4681 ;
  assign n4683 = x73 & n4682 ;
  assign n4684 = x73 | n4682 ;
  assign n4685 = n4398 & n20078 ;
  assign n4686 = n161 & n4685 ;
  assign n20193 = ~n4404 ;
  assign n4687 = n20193 & n4686 ;
  assign n20194 = ~n4686 ;
  assign n4688 = n4404 & n20194 ;
  assign n4689 = n4687 | n4688 ;
  assign n20195 = ~n4689 ;
  assign n4690 = n4684 & n20195 ;
  assign n4691 = n4683 | n4690 ;
  assign n4692 = x74 & n4691 ;
  assign n4693 = x74 | n4691 ;
  assign n4694 = n4407 & n20082 ;
  assign n4695 = n161 & n4694 ;
  assign n4696 = n4413 & n4695 ;
  assign n4697 = n4413 | n4695 ;
  assign n20196 = ~n4696 ;
  assign n4698 = n20196 & n4697 ;
  assign n20197 = ~n4698 ;
  assign n4699 = n4693 & n20197 ;
  assign n4700 = n4692 | n4699 ;
  assign n4701 = x75 & n4700 ;
  assign n4702 = x75 | n4700 ;
  assign n4703 = n4416 & n20086 ;
  assign n4704 = n161 & n4703 ;
  assign n20198 = ~n4422 ;
  assign n4705 = n20198 & n4704 ;
  assign n20199 = ~n4704 ;
  assign n4706 = n4422 & n20199 ;
  assign n4707 = n4705 | n4706 ;
  assign n20200 = ~n4707 ;
  assign n4708 = n4702 & n20200 ;
  assign n4709 = n4701 | n4708 ;
  assign n4710 = x76 & n4709 ;
  assign n4711 = x76 | n4709 ;
  assign n4712 = n4425 & n20090 ;
  assign n4713 = n161 & n4712 ;
  assign n20201 = ~n4431 ;
  assign n4714 = n20201 & n4713 ;
  assign n20202 = ~n4713 ;
  assign n4715 = n4431 & n20202 ;
  assign n4716 = n4714 | n4715 ;
  assign n20203 = ~n4716 ;
  assign n4717 = n4711 & n20203 ;
  assign n4718 = n4710 | n4717 ;
  assign n4719 = x77 & n4718 ;
  assign n4720 = x77 | n4718 ;
  assign n4721 = n4434 & n20094 ;
  assign n4722 = n161 & n4721 ;
  assign n20204 = ~n4440 ;
  assign n4723 = n20204 & n4722 ;
  assign n20205 = ~n4722 ;
  assign n4724 = n4440 & n20205 ;
  assign n4725 = n4723 | n4724 ;
  assign n20206 = ~n4725 ;
  assign n4726 = n4720 & n20206 ;
  assign n4727 = n4719 | n4726 ;
  assign n4728 = x78 & n4727 ;
  assign n4729 = x78 | n4727 ;
  assign n4730 = n4443 & n20098 ;
  assign n4731 = n161 & n4730 ;
  assign n4732 = n4449 & n4731 ;
  assign n4733 = n4449 | n4731 ;
  assign n20207 = ~n4732 ;
  assign n4734 = n20207 & n4733 ;
  assign n20208 = ~n4734 ;
  assign n4735 = n4729 & n20208 ;
  assign n4736 = n4728 | n4735 ;
  assign n4737 = x79 & n4736 ;
  assign n4738 = x79 | n4736 ;
  assign n4739 = n4452 & n20102 ;
  assign n4740 = n161 & n4739 ;
  assign n4741 = n4458 & n4740 ;
  assign n4742 = n4458 | n4740 ;
  assign n20209 = ~n4741 ;
  assign n4743 = n20209 & n4742 ;
  assign n20210 = ~n4743 ;
  assign n4744 = n4738 & n20210 ;
  assign n4745 = n4737 | n4744 ;
  assign n4746 = x80 & n4745 ;
  assign n4747 = x80 | n4745 ;
  assign n4748 = n4461 & n20106 ;
  assign n4749 = n161 & n4748 ;
  assign n20211 = ~n4467 ;
  assign n4750 = n20211 & n4749 ;
  assign n20212 = ~n4749 ;
  assign n4751 = n4467 & n20212 ;
  assign n4752 = n4750 | n4751 ;
  assign n20213 = ~n4752 ;
  assign n4753 = n4747 & n20213 ;
  assign n4754 = n4746 | n4753 ;
  assign n4755 = x81 & n4754 ;
  assign n4756 = x81 | n4754 ;
  assign n4757 = n4470 & n20110 ;
  assign n4758 = n161 & n4757 ;
  assign n20214 = ~n4476 ;
  assign n4759 = n20214 & n4758 ;
  assign n20215 = ~n4758 ;
  assign n4760 = n4476 & n20215 ;
  assign n4761 = n4759 | n4760 ;
  assign n20216 = ~n4761 ;
  assign n4762 = n4756 & n20216 ;
  assign n4763 = n4755 | n4762 ;
  assign n4764 = x82 & n4763 ;
  assign n4765 = x82 | n4763 ;
  assign n4766 = n4479 & n20114 ;
  assign n4767 = n161 & n4766 ;
  assign n20217 = ~n4485 ;
  assign n4768 = n20217 & n4767 ;
  assign n20218 = ~n4767 ;
  assign n4769 = n4485 & n20218 ;
  assign n4770 = n4768 | n4769 ;
  assign n20219 = ~n4770 ;
  assign n4771 = n4765 & n20219 ;
  assign n4772 = n4764 | n4771 ;
  assign n4773 = x83 & n4772 ;
  assign n4774 = x83 | n4772 ;
  assign n4775 = n4488 & n20118 ;
  assign n4776 = n161 & n4775 ;
  assign n20220 = ~n4494 ;
  assign n4777 = n20220 & n4776 ;
  assign n20221 = ~n4776 ;
  assign n4778 = n4494 & n20221 ;
  assign n4779 = n4777 | n4778 ;
  assign n20222 = ~n4779 ;
  assign n4780 = n4774 & n20222 ;
  assign n4781 = n4773 | n4780 ;
  assign n4782 = x84 & n4781 ;
  assign n4783 = x84 | n4781 ;
  assign n4784 = n4497 & n20122 ;
  assign n4785 = n161 & n4784 ;
  assign n20223 = ~n4503 ;
  assign n4786 = n20223 & n4785 ;
  assign n20224 = ~n4785 ;
  assign n4787 = n4503 & n20224 ;
  assign n4788 = n4786 | n4787 ;
  assign n20225 = ~n4788 ;
  assign n4789 = n4783 & n20225 ;
  assign n4790 = n4782 | n4789 ;
  assign n4791 = x85 & n4790 ;
  assign n4792 = x85 | n4790 ;
  assign n4793 = n4506 & n20126 ;
  assign n4794 = n161 & n4793 ;
  assign n20226 = ~n4512 ;
  assign n4795 = n20226 & n4794 ;
  assign n20227 = ~n4794 ;
  assign n4796 = n4512 & n20227 ;
  assign n4797 = n4795 | n4796 ;
  assign n20228 = ~n4797 ;
  assign n4798 = n4792 & n20228 ;
  assign n4799 = n4791 | n4798 ;
  assign n4800 = x86 & n4799 ;
  assign n4801 = x86 | n4799 ;
  assign n4802 = n4515 & n20130 ;
  assign n4803 = n161 & n4802 ;
  assign n20229 = ~n4521 ;
  assign n4804 = n20229 & n4803 ;
  assign n20230 = ~n4803 ;
  assign n4805 = n4521 & n20230 ;
  assign n4806 = n4804 | n4805 ;
  assign n20231 = ~n4806 ;
  assign n4807 = n4801 & n20231 ;
  assign n4808 = n4800 | n4807 ;
  assign n4809 = x87 & n4808 ;
  assign n4810 = x87 | n4808 ;
  assign n4811 = n4524 & n20134 ;
  assign n4812 = n161 & n4811 ;
  assign n20232 = ~n4530 ;
  assign n4813 = n20232 & n4812 ;
  assign n20233 = ~n4812 ;
  assign n4814 = n4530 & n20233 ;
  assign n4815 = n4813 | n4814 ;
  assign n20234 = ~n4815 ;
  assign n4816 = n4810 & n20234 ;
  assign n4817 = n4809 | n4816 ;
  assign n4818 = x88 & n4817 ;
  assign n4819 = x88 | n4817 ;
  assign n4820 = n4533 & n20138 ;
  assign n4821 = n161 & n4820 ;
  assign n20235 = ~n4539 ;
  assign n4822 = n20235 & n4821 ;
  assign n20236 = ~n4821 ;
  assign n4823 = n4539 & n20236 ;
  assign n4824 = n4822 | n4823 ;
  assign n20237 = ~n4824 ;
  assign n4825 = n4819 & n20237 ;
  assign n4826 = n4818 | n4825 ;
  assign n4827 = x89 & n4826 ;
  assign n4828 = x89 | n4826 ;
  assign n4829 = n4542 & n20142 ;
  assign n4830 = n161 & n4829 ;
  assign n20238 = ~n4548 ;
  assign n4831 = n20238 & n4830 ;
  assign n20239 = ~n4830 ;
  assign n4832 = n4548 & n20239 ;
  assign n4833 = n4831 | n4832 ;
  assign n20240 = ~n4833 ;
  assign n4834 = n4828 & n20240 ;
  assign n4835 = n4827 | n4834 ;
  assign n4836 = x90 & n4835 ;
  assign n4837 = x90 | n4835 ;
  assign n4838 = n4551 & n20146 ;
  assign n4839 = n161 & n4838 ;
  assign n20241 = ~n4557 ;
  assign n4840 = n20241 & n4839 ;
  assign n20242 = ~n4839 ;
  assign n4841 = n4557 & n20242 ;
  assign n4842 = n4840 | n4841 ;
  assign n20243 = ~n4842 ;
  assign n4843 = n4837 & n20243 ;
  assign n4844 = n4836 | n4843 ;
  assign n4845 = x91 & n4844 ;
  assign n4846 = x91 | n4844 ;
  assign n4847 = n4560 & n20150 ;
  assign n4848 = n161 & n4847 ;
  assign n20244 = ~n4566 ;
  assign n4849 = n20244 & n4848 ;
  assign n20245 = ~n4848 ;
  assign n4850 = n4566 & n20245 ;
  assign n4851 = n4849 | n4850 ;
  assign n20246 = ~n4851 ;
  assign n4852 = n4846 & n20246 ;
  assign n4853 = n4845 | n4852 ;
  assign n4854 = x92 & n4853 ;
  assign n4855 = x92 | n4853 ;
  assign n4856 = n4569 & n20154 ;
  assign n4857 = n161 & n4856 ;
  assign n20247 = ~n4575 ;
  assign n4858 = n20247 & n4857 ;
  assign n20248 = ~n4857 ;
  assign n4859 = n4575 & n20248 ;
  assign n4860 = n4858 | n4859 ;
  assign n20249 = ~n4860 ;
  assign n4861 = n4855 & n20249 ;
  assign n4862 = n4854 | n4861 ;
  assign n4863 = x93 & n4862 ;
  assign n4864 = x93 | n4862 ;
  assign n4865 = n4578 & n20158 ;
  assign n4866 = n161 & n4865 ;
  assign n20250 = ~n4584 ;
  assign n4867 = n20250 & n4866 ;
  assign n20251 = ~n4866 ;
  assign n4868 = n4584 & n20251 ;
  assign n4869 = n4867 | n4868 ;
  assign n20252 = ~n4869 ;
  assign n4870 = n4864 & n20252 ;
  assign n4871 = n4863 | n4870 ;
  assign n4872 = x94 & n4871 ;
  assign n4873 = x94 | n4871 ;
  assign n4874 = n4587 & n20162 ;
  assign n4875 = n161 & n4874 ;
  assign n20253 = ~n4593 ;
  assign n4876 = n20253 & n4875 ;
  assign n20254 = ~n4875 ;
  assign n4877 = n4593 & n20254 ;
  assign n4878 = n4876 | n4877 ;
  assign n20255 = ~n4878 ;
  assign n4879 = n4873 & n20255 ;
  assign n4880 = n4872 | n4879 ;
  assign n4882 = x95 | n4880 ;
  assign n20256 = ~n4608 ;
  assign n4883 = n20256 & n4882 ;
  assign n4881 = x95 & n4880 ;
  assign n20257 = ~n4331 ;
  assign n4332 = x96 & n20257 ;
  assign n4884 = n18413 | n4332 ;
  assign n4885 = n4610 | n4884 ;
  assign n4886 = n4881 | n4885 ;
  assign n4887 = n4883 | n4886 ;
  assign n20258 = ~n4610 ;
  assign n4888 = n20258 & n4887 ;
  assign n20259 = ~n4881 ;
  assign n4889 = n20259 & n4882 ;
  assign n160 = ~n4888 ;
  assign n4890 = n160 & n4889 ;
  assign n4891 = n4608 & n4890 ;
  assign n4892 = n4608 | n4890 ;
  assign n20261 = ~n4891 ;
  assign n4893 = n20261 & n4892 ;
  assign n20262 = ~x30 ;
  assign n4894 = n20262 & x64 ;
  assign n4895 = x65 | n4894 ;
  assign n4896 = x64 & n160 ;
  assign n20263 = ~n4896 ;
  assign n4897 = x31 & n20263 ;
  assign n4898 = n4611 & n160 ;
  assign n4899 = n4897 | n4898 ;
  assign n4900 = x65 & n4894 ;
  assign n20264 = ~n4900 ;
  assign n4901 = n4899 & n20264 ;
  assign n20265 = ~n4901 ;
  assign n4902 = n4895 & n20265 ;
  assign n4903 = x66 | n4902 ;
  assign n4904 = x66 & n4902 ;
  assign n4905 = n20172 & n4613 ;
  assign n4906 = n160 & n4905 ;
  assign n4907 = n4617 & n4906 ;
  assign n4908 = n4617 | n4906 ;
  assign n20266 = ~n4907 ;
  assign n4909 = n20266 & n4908 ;
  assign n20267 = ~n4904 ;
  assign n4910 = n20267 & n4909 ;
  assign n20268 = ~n4910 ;
  assign n4911 = n4903 & n20268 ;
  assign n4913 = x67 | n4911 ;
  assign n4912 = x67 & n4911 ;
  assign n20269 = ~n4620 ;
  assign n4914 = n20269 & n4621 ;
  assign n4915 = n160 & n4914 ;
  assign n4916 = n4626 & n4915 ;
  assign n4917 = n4626 | n4915 ;
  assign n20270 = ~n4916 ;
  assign n4918 = n20270 & n4917 ;
  assign n20271 = ~n4912 ;
  assign n4919 = n20271 & n4918 ;
  assign n20272 = ~n4919 ;
  assign n4920 = n4913 & n20272 ;
  assign n4921 = x68 | n4920 ;
  assign n4922 = x68 & n4920 ;
  assign n20273 = ~n4629 ;
  assign n4923 = n20273 & n4630 ;
  assign n4924 = n160 & n4923 ;
  assign n4925 = n4635 & n4924 ;
  assign n4926 = n4635 | n4924 ;
  assign n20274 = ~n4925 ;
  assign n4927 = n20274 & n4926 ;
  assign n20275 = ~n4922 ;
  assign n4928 = n20275 & n4927 ;
  assign n20276 = ~n4928 ;
  assign n4929 = n4921 & n20276 ;
  assign n4930 = x69 | n4929 ;
  assign n4931 = x69 & n4929 ;
  assign n20277 = ~n4638 ;
  assign n4932 = n20277 & n4639 ;
  assign n4933 = n160 & n4932 ;
  assign n4934 = n4644 & n4933 ;
  assign n4935 = n4644 | n4933 ;
  assign n20278 = ~n4934 ;
  assign n4936 = n20278 & n4935 ;
  assign n20279 = ~n4931 ;
  assign n4937 = n20279 & n4936 ;
  assign n20280 = ~n4937 ;
  assign n4938 = n4930 & n20280 ;
  assign n4939 = x70 | n4938 ;
  assign n4940 = x70 & n4938 ;
  assign n20281 = ~n4647 ;
  assign n4941 = n20281 & n4648 ;
  assign n4942 = n160 & n4941 ;
  assign n4943 = n4653 & n4942 ;
  assign n4944 = n4653 | n4942 ;
  assign n20282 = ~n4943 ;
  assign n4945 = n20282 & n4944 ;
  assign n20283 = ~n4940 ;
  assign n4946 = n20283 & n4945 ;
  assign n20284 = ~n4946 ;
  assign n4947 = n4939 & n20284 ;
  assign n4948 = x71 | n4947 ;
  assign n4949 = x71 & n4947 ;
  assign n20285 = ~n4656 ;
  assign n4950 = n20285 & n4657 ;
  assign n4951 = n160 & n4950 ;
  assign n4952 = n20187 & n4951 ;
  assign n20286 = ~n4951 ;
  assign n4953 = n4662 & n20286 ;
  assign n4954 = n4952 | n4953 ;
  assign n20287 = ~n4949 ;
  assign n4955 = n20287 & n4954 ;
  assign n20288 = ~n4955 ;
  assign n4956 = n4948 & n20288 ;
  assign n4957 = x72 | n4956 ;
  assign n4958 = x72 & n4956 ;
  assign n20289 = ~n4665 ;
  assign n4959 = n20289 & n4666 ;
  assign n4960 = n160 & n4959 ;
  assign n4961 = n4671 & n4960 ;
  assign n4962 = n4671 | n4960 ;
  assign n20290 = ~n4961 ;
  assign n4963 = n20290 & n4962 ;
  assign n20291 = ~n4958 ;
  assign n4964 = n20291 & n4963 ;
  assign n20292 = ~n4964 ;
  assign n4965 = n4957 & n20292 ;
  assign n4966 = x73 | n4965 ;
  assign n4967 = x73 & n4965 ;
  assign n20293 = ~n4674 ;
  assign n4968 = n20293 & n4675 ;
  assign n4969 = n160 & n4968 ;
  assign n4970 = n20192 & n4969 ;
  assign n20294 = ~n4969 ;
  assign n4971 = n4680 & n20294 ;
  assign n4972 = n4970 | n4971 ;
  assign n20295 = ~n4967 ;
  assign n4973 = n20295 & n4972 ;
  assign n20296 = ~n4973 ;
  assign n4974 = n4966 & n20296 ;
  assign n4975 = x74 | n4974 ;
  assign n4976 = x74 & n4974 ;
  assign n20297 = ~n4683 ;
  assign n4977 = n20297 & n4684 ;
  assign n4978 = n160 & n4977 ;
  assign n4979 = n20195 & n4978 ;
  assign n20298 = ~n4978 ;
  assign n4980 = n4689 & n20298 ;
  assign n4981 = n4979 | n4980 ;
  assign n20299 = ~n4976 ;
  assign n4982 = n20299 & n4981 ;
  assign n20300 = ~n4982 ;
  assign n4983 = n4975 & n20300 ;
  assign n4984 = x75 | n4983 ;
  assign n4985 = x75 & n4983 ;
  assign n20301 = ~n4692 ;
  assign n4986 = n20301 & n4693 ;
  assign n4987 = n160 & n4986 ;
  assign n4988 = n4698 & n4987 ;
  assign n4989 = n4698 | n4987 ;
  assign n20302 = ~n4988 ;
  assign n4990 = n20302 & n4989 ;
  assign n20303 = ~n4985 ;
  assign n4991 = n20303 & n4990 ;
  assign n20304 = ~n4991 ;
  assign n4992 = n4984 & n20304 ;
  assign n4993 = x76 | n4992 ;
  assign n4994 = x76 & n4992 ;
  assign n20305 = ~n4701 ;
  assign n4995 = n20305 & n4702 ;
  assign n4996 = n160 & n4995 ;
  assign n4997 = n4707 & n4996 ;
  assign n4998 = n4707 | n4996 ;
  assign n20306 = ~n4997 ;
  assign n4999 = n20306 & n4998 ;
  assign n20307 = ~n4994 ;
  assign n5000 = n20307 & n4999 ;
  assign n20308 = ~n5000 ;
  assign n5001 = n4993 & n20308 ;
  assign n5002 = x77 | n5001 ;
  assign n5003 = x77 & n5001 ;
  assign n20309 = ~n4710 ;
  assign n5004 = n20309 & n4711 ;
  assign n5005 = n160 & n5004 ;
  assign n5006 = n4716 & n5005 ;
  assign n5007 = n4716 | n5005 ;
  assign n20310 = ~n5006 ;
  assign n5008 = n20310 & n5007 ;
  assign n20311 = ~n5003 ;
  assign n5009 = n20311 & n5008 ;
  assign n20312 = ~n5009 ;
  assign n5010 = n5002 & n20312 ;
  assign n5011 = x78 | n5010 ;
  assign n5012 = x78 & n5010 ;
  assign n20313 = ~n4719 ;
  assign n5013 = n20313 & n4720 ;
  assign n5014 = n160 & n5013 ;
  assign n5015 = n4725 & n5014 ;
  assign n5016 = n4725 | n5014 ;
  assign n20314 = ~n5015 ;
  assign n5017 = n20314 & n5016 ;
  assign n20315 = ~n5012 ;
  assign n5018 = n20315 & n5017 ;
  assign n20316 = ~n5018 ;
  assign n5019 = n5011 & n20316 ;
  assign n5020 = x79 | n5019 ;
  assign n5021 = x79 & n5019 ;
  assign n20317 = ~n4728 ;
  assign n5022 = n20317 & n4729 ;
  assign n5023 = n160 & n5022 ;
  assign n5024 = n4734 & n5023 ;
  assign n5025 = n4734 | n5023 ;
  assign n20318 = ~n5024 ;
  assign n5026 = n20318 & n5025 ;
  assign n20319 = ~n5021 ;
  assign n5027 = n20319 & n5026 ;
  assign n20320 = ~n5027 ;
  assign n5028 = n5020 & n20320 ;
  assign n5029 = x80 | n5028 ;
  assign n5030 = x80 & n5028 ;
  assign n20321 = ~n4737 ;
  assign n5031 = n20321 & n4738 ;
  assign n5032 = n160 & n5031 ;
  assign n5033 = n4743 & n5032 ;
  assign n5034 = n4743 | n5032 ;
  assign n20322 = ~n5033 ;
  assign n5035 = n20322 & n5034 ;
  assign n20323 = ~n5030 ;
  assign n5036 = n20323 & n5035 ;
  assign n20324 = ~n5036 ;
  assign n5037 = n5029 & n20324 ;
  assign n5038 = x81 | n5037 ;
  assign n5039 = x81 & n5037 ;
  assign n20325 = ~n4746 ;
  assign n5040 = n20325 & n4747 ;
  assign n5041 = n160 & n5040 ;
  assign n5042 = n20213 & n5041 ;
  assign n20326 = ~n5041 ;
  assign n5043 = n4752 & n20326 ;
  assign n5044 = n5042 | n5043 ;
  assign n20327 = ~n5039 ;
  assign n5045 = n20327 & n5044 ;
  assign n20328 = ~n5045 ;
  assign n5046 = n5038 & n20328 ;
  assign n5047 = x82 | n5046 ;
  assign n5048 = x82 & n5046 ;
  assign n20329 = ~n4755 ;
  assign n5049 = n20329 & n4756 ;
  assign n5050 = n160 & n5049 ;
  assign n5051 = n4761 & n5050 ;
  assign n5052 = n4761 | n5050 ;
  assign n20330 = ~n5051 ;
  assign n5053 = n20330 & n5052 ;
  assign n20331 = ~n5048 ;
  assign n5054 = n20331 & n5053 ;
  assign n20332 = ~n5054 ;
  assign n5055 = n5047 & n20332 ;
  assign n5056 = x83 | n5055 ;
  assign n5057 = x83 & n5055 ;
  assign n20333 = ~n4764 ;
  assign n5058 = n20333 & n4765 ;
  assign n5059 = n160 & n5058 ;
  assign n5060 = n4770 & n5059 ;
  assign n5061 = n4770 | n5059 ;
  assign n20334 = ~n5060 ;
  assign n5062 = n20334 & n5061 ;
  assign n20335 = ~n5057 ;
  assign n5063 = n20335 & n5062 ;
  assign n20336 = ~n5063 ;
  assign n5064 = n5056 & n20336 ;
  assign n5065 = x84 | n5064 ;
  assign n5066 = x84 & n5064 ;
  assign n20337 = ~n4773 ;
  assign n5067 = n20337 & n4774 ;
  assign n5068 = n160 & n5067 ;
  assign n5069 = n4779 & n5068 ;
  assign n5070 = n4779 | n5068 ;
  assign n20338 = ~n5069 ;
  assign n5071 = n20338 & n5070 ;
  assign n20339 = ~n5066 ;
  assign n5072 = n20339 & n5071 ;
  assign n20340 = ~n5072 ;
  assign n5073 = n5065 & n20340 ;
  assign n5074 = x85 | n5073 ;
  assign n5075 = x85 & n5073 ;
  assign n20341 = ~n4782 ;
  assign n5076 = n20341 & n4783 ;
  assign n5077 = n160 & n5076 ;
  assign n5078 = n4788 & n5077 ;
  assign n5079 = n4788 | n5077 ;
  assign n20342 = ~n5078 ;
  assign n5080 = n20342 & n5079 ;
  assign n20343 = ~n5075 ;
  assign n5081 = n20343 & n5080 ;
  assign n20344 = ~n5081 ;
  assign n5082 = n5074 & n20344 ;
  assign n5083 = x86 | n5082 ;
  assign n5084 = x86 & n5082 ;
  assign n20345 = ~n4791 ;
  assign n5085 = n20345 & n4792 ;
  assign n5086 = n160 & n5085 ;
  assign n5087 = n4797 & n5086 ;
  assign n5088 = n4797 | n5086 ;
  assign n20346 = ~n5087 ;
  assign n5089 = n20346 & n5088 ;
  assign n20347 = ~n5084 ;
  assign n5090 = n20347 & n5089 ;
  assign n20348 = ~n5090 ;
  assign n5091 = n5083 & n20348 ;
  assign n5092 = x87 | n5091 ;
  assign n5093 = x87 & n5091 ;
  assign n20349 = ~n4800 ;
  assign n5094 = n20349 & n4801 ;
  assign n5095 = n160 & n5094 ;
  assign n5096 = n4806 & n5095 ;
  assign n5097 = n4806 | n5095 ;
  assign n20350 = ~n5096 ;
  assign n5098 = n20350 & n5097 ;
  assign n20351 = ~n5093 ;
  assign n5099 = n20351 & n5098 ;
  assign n20352 = ~n5099 ;
  assign n5100 = n5092 & n20352 ;
  assign n5101 = x88 | n5100 ;
  assign n5102 = x88 & n5100 ;
  assign n20353 = ~n4809 ;
  assign n5103 = n20353 & n4810 ;
  assign n5104 = n160 & n5103 ;
  assign n5105 = n4815 & n5104 ;
  assign n5106 = n4815 | n5104 ;
  assign n20354 = ~n5105 ;
  assign n5107 = n20354 & n5106 ;
  assign n20355 = ~n5102 ;
  assign n5108 = n20355 & n5107 ;
  assign n20356 = ~n5108 ;
  assign n5109 = n5101 & n20356 ;
  assign n5110 = x89 | n5109 ;
  assign n5111 = x89 & n5109 ;
  assign n20357 = ~n4818 ;
  assign n5112 = n20357 & n4819 ;
  assign n5113 = n160 & n5112 ;
  assign n5114 = n20237 & n5113 ;
  assign n20358 = ~n5113 ;
  assign n5115 = n4824 & n20358 ;
  assign n5116 = n5114 | n5115 ;
  assign n20359 = ~n5111 ;
  assign n5117 = n20359 & n5116 ;
  assign n20360 = ~n5117 ;
  assign n5118 = n5110 & n20360 ;
  assign n5119 = x90 | n5118 ;
  assign n5120 = x90 & n5118 ;
  assign n20361 = ~n4827 ;
  assign n5121 = n20361 & n4828 ;
  assign n5122 = n160 & n5121 ;
  assign n5123 = n20240 & n5122 ;
  assign n20362 = ~n5122 ;
  assign n5124 = n4833 & n20362 ;
  assign n5125 = n5123 | n5124 ;
  assign n20363 = ~n5120 ;
  assign n5126 = n20363 & n5125 ;
  assign n20364 = ~n5126 ;
  assign n5127 = n5119 & n20364 ;
  assign n5128 = x91 | n5127 ;
  assign n5129 = x91 & n5127 ;
  assign n20365 = ~n4836 ;
  assign n5130 = n20365 & n4837 ;
  assign n5131 = n160 & n5130 ;
  assign n5132 = n4842 & n5131 ;
  assign n5133 = n4842 | n5131 ;
  assign n20366 = ~n5132 ;
  assign n5134 = n20366 & n5133 ;
  assign n20367 = ~n5129 ;
  assign n5135 = n20367 & n5134 ;
  assign n20368 = ~n5135 ;
  assign n5136 = n5128 & n20368 ;
  assign n5137 = x92 | n5136 ;
  assign n5138 = x92 & n5136 ;
  assign n20369 = ~n4845 ;
  assign n5139 = n20369 & n4846 ;
  assign n5140 = n160 & n5139 ;
  assign n5141 = n4851 & n5140 ;
  assign n5142 = n4851 | n5140 ;
  assign n20370 = ~n5141 ;
  assign n5143 = n20370 & n5142 ;
  assign n20371 = ~n5138 ;
  assign n5144 = n20371 & n5143 ;
  assign n20372 = ~n5144 ;
  assign n5145 = n5137 & n20372 ;
  assign n5146 = x93 | n5145 ;
  assign n5147 = x93 & n5145 ;
  assign n20373 = ~n4854 ;
  assign n5148 = n20373 & n4855 ;
  assign n5149 = n160 & n5148 ;
  assign n5150 = n4860 & n5149 ;
  assign n5151 = n4860 | n5149 ;
  assign n20374 = ~n5150 ;
  assign n5152 = n20374 & n5151 ;
  assign n20375 = ~n5147 ;
  assign n5153 = n20375 & n5152 ;
  assign n20376 = ~n5153 ;
  assign n5154 = n5146 & n20376 ;
  assign n5155 = x94 | n5154 ;
  assign n5156 = x94 & n5154 ;
  assign n20377 = ~n4863 ;
  assign n5157 = n20377 & n4864 ;
  assign n5158 = n160 & n5157 ;
  assign n5159 = n4869 & n5158 ;
  assign n5160 = n4869 | n5158 ;
  assign n20378 = ~n5159 ;
  assign n5161 = n20378 & n5160 ;
  assign n20379 = ~n5156 ;
  assign n5162 = n20379 & n5161 ;
  assign n20380 = ~n5162 ;
  assign n5163 = n5155 & n20380 ;
  assign n5164 = x95 | n5163 ;
  assign n5165 = x95 & n5163 ;
  assign n20381 = ~n4872 ;
  assign n5166 = n20381 & n4873 ;
  assign n5167 = n160 & n5166 ;
  assign n5168 = n4878 & n5167 ;
  assign n5169 = n4878 | n5167 ;
  assign n20382 = ~n5168 ;
  assign n5170 = n20382 & n5169 ;
  assign n20383 = ~n5165 ;
  assign n5171 = n20383 & n5170 ;
  assign n20384 = ~n5171 ;
  assign n5172 = n5164 & n20384 ;
  assign n5173 = x96 | n5172 ;
  assign n5174 = x96 & n5172 ;
  assign n20385 = ~n5174 ;
  assign n5175 = n4893 & n20385 ;
  assign n20386 = ~n5175 ;
  assign n5176 = n5173 & n20386 ;
  assign n5178 = x97 & n5176 ;
  assign n5179 = n18408 | n5178 ;
  assign n5177 = x97 | n5176 ;
  assign n4333 = n18418 & n4331 ;
  assign n5180 = n4333 & n4887 ;
  assign n5181 = n21884 | n5180 ;
  assign n20387 = ~n5181 ;
  assign n5185 = n5177 & n20387 ;
  assign n5186 = n5179 | n5185 ;
  assign n5188 = n5173 & n20385 ;
  assign n159 = ~n5186 ;
  assign n5189 = n159 & n5188 ;
  assign n20389 = ~n4893 ;
  assign n5190 = n20389 & n5189 ;
  assign n20390 = ~n5189 ;
  assign n5191 = n4893 & n20390 ;
  assign n5192 = n5190 | n5191 ;
  assign n20391 = ~x29 ;
  assign n5193 = n20391 & x64 ;
  assign n5195 = x65 | n5193 ;
  assign n5194 = x65 & n5193 ;
  assign n5196 = x64 & n159 ;
  assign n5197 = x30 & n5196 ;
  assign n5198 = x30 | n5196 ;
  assign n20392 = ~n5197 ;
  assign n5199 = n20392 & n5198 ;
  assign n20393 = ~n5194 ;
  assign n5200 = n20393 & n5199 ;
  assign n20394 = ~n5200 ;
  assign n5201 = n5195 & n20394 ;
  assign n5202 = x66 & n5201 ;
  assign n5203 = x66 | n5201 ;
  assign n5204 = n4895 & n159 ;
  assign n5205 = n4901 & n5204 ;
  assign n5206 = n20264 & n5204 ;
  assign n5207 = n4899 | n5206 ;
  assign n20395 = ~n5205 ;
  assign n5208 = n20395 & n5207 ;
  assign n20396 = ~n5208 ;
  assign n5209 = n5203 & n20396 ;
  assign n5210 = n5202 | n5209 ;
  assign n5211 = x67 & n5210 ;
  assign n5187 = n4903 & n159 ;
  assign n5212 = n20267 & n5187 ;
  assign n5213 = n4909 | n5212 ;
  assign n5214 = n4910 & n5187 ;
  assign n20397 = ~n5214 ;
  assign n5215 = n5213 & n20397 ;
  assign n5216 = x67 | n5210 ;
  assign n20398 = ~n5215 ;
  assign n5217 = n20398 & n5216 ;
  assign n5218 = n5211 | n5217 ;
  assign n5219 = x68 & n5218 ;
  assign n5220 = x68 | n5218 ;
  assign n5221 = n4913 & n159 ;
  assign n5222 = n4919 & n5221 ;
  assign n5223 = n20271 & n5221 ;
  assign n5224 = n4918 | n5223 ;
  assign n20399 = ~n5222 ;
  assign n5225 = n20399 & n5224 ;
  assign n20400 = ~n5225 ;
  assign n5226 = n5220 & n20400 ;
  assign n5227 = n5219 | n5226 ;
  assign n5228 = x69 & n5227 ;
  assign n5229 = x69 | n5227 ;
  assign n5230 = n4921 & n20275 ;
  assign n5231 = n159 & n5230 ;
  assign n20401 = ~n4927 ;
  assign n5232 = n20401 & n5231 ;
  assign n20402 = ~n5231 ;
  assign n5233 = n4927 & n20402 ;
  assign n5234 = n5232 | n5233 ;
  assign n20403 = ~n5234 ;
  assign n5235 = n5229 & n20403 ;
  assign n5236 = n5228 | n5235 ;
  assign n5237 = x70 & n5236 ;
  assign n5238 = x70 | n5236 ;
  assign n5239 = n4930 & n20279 ;
  assign n5240 = n159 & n5239 ;
  assign n5241 = n4936 & n5240 ;
  assign n5242 = n4936 | n5240 ;
  assign n20404 = ~n5241 ;
  assign n5243 = n20404 & n5242 ;
  assign n20405 = ~n5243 ;
  assign n5244 = n5238 & n20405 ;
  assign n5245 = n5237 | n5244 ;
  assign n5246 = x71 & n5245 ;
  assign n5247 = x71 | n5245 ;
  assign n5248 = n4939 & n20283 ;
  assign n5249 = n159 & n5248 ;
  assign n5250 = n4945 & n5249 ;
  assign n5251 = n4945 | n5249 ;
  assign n20406 = ~n5250 ;
  assign n5252 = n20406 & n5251 ;
  assign n20407 = ~n5252 ;
  assign n5253 = n5247 & n20407 ;
  assign n5254 = n5246 | n5253 ;
  assign n5255 = x72 & n5254 ;
  assign n5256 = x72 | n5254 ;
  assign n5257 = n4948 & n20287 ;
  assign n5258 = n159 & n5257 ;
  assign n20408 = ~n4954 ;
  assign n5259 = n20408 & n5258 ;
  assign n20409 = ~n5258 ;
  assign n5260 = n4954 & n20409 ;
  assign n5261 = n5259 | n5260 ;
  assign n20410 = ~n5261 ;
  assign n5262 = n5256 & n20410 ;
  assign n5263 = n5255 | n5262 ;
  assign n5264 = x73 & n5263 ;
  assign n5265 = x73 | n5263 ;
  assign n5266 = n4957 & n20291 ;
  assign n5267 = n159 & n5266 ;
  assign n20411 = ~n4963 ;
  assign n5268 = n20411 & n5267 ;
  assign n20412 = ~n5267 ;
  assign n5269 = n4963 & n20412 ;
  assign n5270 = n5268 | n5269 ;
  assign n20413 = ~n5270 ;
  assign n5271 = n5265 & n20413 ;
  assign n5272 = n5264 | n5271 ;
  assign n5273 = x74 & n5272 ;
  assign n5274 = x74 | n5272 ;
  assign n5275 = n4966 & n20295 ;
  assign n5276 = n159 & n5275 ;
  assign n20414 = ~n4972 ;
  assign n5277 = n20414 & n5276 ;
  assign n20415 = ~n5276 ;
  assign n5278 = n4972 & n20415 ;
  assign n5279 = n5277 | n5278 ;
  assign n20416 = ~n5279 ;
  assign n5280 = n5274 & n20416 ;
  assign n5281 = n5273 | n5280 ;
  assign n5282 = x75 & n5281 ;
  assign n5283 = x75 | n5281 ;
  assign n5284 = n4975 & n20299 ;
  assign n5285 = n159 & n5284 ;
  assign n20417 = ~n4981 ;
  assign n5286 = n20417 & n5285 ;
  assign n20418 = ~n5285 ;
  assign n5287 = n4981 & n20418 ;
  assign n5288 = n5286 | n5287 ;
  assign n20419 = ~n5288 ;
  assign n5289 = n5283 & n20419 ;
  assign n5290 = n5282 | n5289 ;
  assign n5291 = x76 & n5290 ;
  assign n5292 = x76 | n5290 ;
  assign n5293 = n4984 & n20303 ;
  assign n5294 = n159 & n5293 ;
  assign n20420 = ~n4990 ;
  assign n5295 = n20420 & n5294 ;
  assign n20421 = ~n5294 ;
  assign n5296 = n4990 & n20421 ;
  assign n5297 = n5295 | n5296 ;
  assign n20422 = ~n5297 ;
  assign n5298 = n5292 & n20422 ;
  assign n5299 = n5291 | n5298 ;
  assign n5300 = x77 & n5299 ;
  assign n5301 = x77 | n5299 ;
  assign n5302 = n4993 & n20307 ;
  assign n5303 = n159 & n5302 ;
  assign n5304 = n4999 & n5303 ;
  assign n5305 = n4999 | n5303 ;
  assign n20423 = ~n5304 ;
  assign n5306 = n20423 & n5305 ;
  assign n20424 = ~n5306 ;
  assign n5307 = n5301 & n20424 ;
  assign n5308 = n5300 | n5307 ;
  assign n5309 = x78 & n5308 ;
  assign n5310 = x78 | n5308 ;
  assign n5311 = n5002 & n20311 ;
  assign n5312 = n159 & n5311 ;
  assign n5313 = n5008 & n5312 ;
  assign n5314 = n5008 | n5312 ;
  assign n20425 = ~n5313 ;
  assign n5315 = n20425 & n5314 ;
  assign n20426 = ~n5315 ;
  assign n5316 = n5310 & n20426 ;
  assign n5317 = n5309 | n5316 ;
  assign n5318 = x79 & n5317 ;
  assign n5319 = x79 | n5317 ;
  assign n5320 = n5011 & n20315 ;
  assign n5321 = n159 & n5320 ;
  assign n5322 = n5017 & n5321 ;
  assign n5323 = n5017 | n5321 ;
  assign n20427 = ~n5322 ;
  assign n5324 = n20427 & n5323 ;
  assign n20428 = ~n5324 ;
  assign n5325 = n5319 & n20428 ;
  assign n5326 = n5318 | n5325 ;
  assign n5327 = x80 & n5326 ;
  assign n5328 = x80 | n5326 ;
  assign n5329 = n5020 & n20319 ;
  assign n5330 = n159 & n5329 ;
  assign n20429 = ~n5026 ;
  assign n5331 = n20429 & n5330 ;
  assign n20430 = ~n5330 ;
  assign n5332 = n5026 & n20430 ;
  assign n5333 = n5331 | n5332 ;
  assign n20431 = ~n5333 ;
  assign n5334 = n5328 & n20431 ;
  assign n5335 = n5327 | n5334 ;
  assign n5336 = x81 & n5335 ;
  assign n5337 = x81 | n5335 ;
  assign n5338 = n5029 & n20323 ;
  assign n5339 = n159 & n5338 ;
  assign n20432 = ~n5035 ;
  assign n5340 = n20432 & n5339 ;
  assign n20433 = ~n5339 ;
  assign n5341 = n5035 & n20433 ;
  assign n5342 = n5340 | n5341 ;
  assign n20434 = ~n5342 ;
  assign n5343 = n5337 & n20434 ;
  assign n5344 = n5336 | n5343 ;
  assign n5345 = x82 & n5344 ;
  assign n5346 = x82 | n5344 ;
  assign n5347 = n5038 & n20327 ;
  assign n5348 = n159 & n5347 ;
  assign n20435 = ~n5044 ;
  assign n5349 = n20435 & n5348 ;
  assign n20436 = ~n5348 ;
  assign n5350 = n5044 & n20436 ;
  assign n5351 = n5349 | n5350 ;
  assign n20437 = ~n5351 ;
  assign n5352 = n5346 & n20437 ;
  assign n5353 = n5345 | n5352 ;
  assign n5354 = x83 & n5353 ;
  assign n5355 = x83 | n5353 ;
  assign n5356 = n5047 & n20331 ;
  assign n5357 = n159 & n5356 ;
  assign n5358 = n5053 & n5357 ;
  assign n5359 = n5053 | n5357 ;
  assign n20438 = ~n5358 ;
  assign n5360 = n20438 & n5359 ;
  assign n20439 = ~n5360 ;
  assign n5361 = n5355 & n20439 ;
  assign n5362 = n5354 | n5361 ;
  assign n5363 = x84 & n5362 ;
  assign n5364 = x84 | n5362 ;
  assign n5365 = n5056 & n20335 ;
  assign n5366 = n159 & n5365 ;
  assign n5367 = n5062 & n5366 ;
  assign n5368 = n5062 | n5366 ;
  assign n20440 = ~n5367 ;
  assign n5369 = n20440 & n5368 ;
  assign n20441 = ~n5369 ;
  assign n5370 = n5364 & n20441 ;
  assign n5371 = n5363 | n5370 ;
  assign n5372 = x85 & n5371 ;
  assign n5373 = x85 | n5371 ;
  assign n5374 = n5065 & n20339 ;
  assign n5375 = n159 & n5374 ;
  assign n5376 = n5071 & n5375 ;
  assign n5377 = n5071 | n5375 ;
  assign n20442 = ~n5376 ;
  assign n5378 = n20442 & n5377 ;
  assign n20443 = ~n5378 ;
  assign n5379 = n5373 & n20443 ;
  assign n5380 = n5372 | n5379 ;
  assign n5381 = x86 & n5380 ;
  assign n5382 = x86 | n5380 ;
  assign n5383 = n5074 & n20343 ;
  assign n5384 = n159 & n5383 ;
  assign n5385 = n5080 & n5384 ;
  assign n5386 = n5080 | n5384 ;
  assign n20444 = ~n5385 ;
  assign n5387 = n20444 & n5386 ;
  assign n20445 = ~n5387 ;
  assign n5388 = n5382 & n20445 ;
  assign n5389 = n5381 | n5388 ;
  assign n5390 = x87 & n5389 ;
  assign n5391 = x87 | n5389 ;
  assign n5392 = n5083 & n20347 ;
  assign n5393 = n159 & n5392 ;
  assign n5394 = n5089 & n5393 ;
  assign n5395 = n5089 | n5393 ;
  assign n20446 = ~n5394 ;
  assign n5396 = n20446 & n5395 ;
  assign n20447 = ~n5396 ;
  assign n5397 = n5391 & n20447 ;
  assign n5398 = n5390 | n5397 ;
  assign n5399 = x88 & n5398 ;
  assign n5400 = x88 | n5398 ;
  assign n5401 = n5092 & n20351 ;
  assign n5402 = n159 & n5401 ;
  assign n5403 = n5098 & n5402 ;
  assign n5404 = n5098 | n5402 ;
  assign n20448 = ~n5403 ;
  assign n5405 = n20448 & n5404 ;
  assign n20449 = ~n5405 ;
  assign n5406 = n5400 & n20449 ;
  assign n5407 = n5399 | n5406 ;
  assign n5408 = x89 & n5407 ;
  assign n5409 = x89 | n5407 ;
  assign n5410 = n5101 & n20355 ;
  assign n5411 = n159 & n5410 ;
  assign n5412 = n5107 & n5411 ;
  assign n5413 = n5107 | n5411 ;
  assign n20450 = ~n5412 ;
  assign n5414 = n20450 & n5413 ;
  assign n20451 = ~n5414 ;
  assign n5415 = n5409 & n20451 ;
  assign n5416 = n5408 | n5415 ;
  assign n5417 = x90 & n5416 ;
  assign n5418 = x90 | n5416 ;
  assign n5419 = n5110 & n20359 ;
  assign n5420 = n159 & n5419 ;
  assign n20452 = ~n5116 ;
  assign n5421 = n20452 & n5420 ;
  assign n20453 = ~n5420 ;
  assign n5422 = n5116 & n20453 ;
  assign n5423 = n5421 | n5422 ;
  assign n20454 = ~n5423 ;
  assign n5424 = n5418 & n20454 ;
  assign n5425 = n5417 | n5424 ;
  assign n5426 = x91 & n5425 ;
  assign n5427 = x91 | n5425 ;
  assign n5428 = n5119 & n20363 ;
  assign n5429 = n159 & n5428 ;
  assign n20455 = ~n5125 ;
  assign n5430 = n20455 & n5429 ;
  assign n20456 = ~n5429 ;
  assign n5431 = n5125 & n20456 ;
  assign n5432 = n5430 | n5431 ;
  assign n20457 = ~n5432 ;
  assign n5433 = n5427 & n20457 ;
  assign n5434 = n5426 | n5433 ;
  assign n5435 = x92 & n5434 ;
  assign n5436 = x92 | n5434 ;
  assign n5437 = n5128 & n20367 ;
  assign n5438 = n159 & n5437 ;
  assign n5439 = n5134 & n5438 ;
  assign n5440 = n5134 | n5438 ;
  assign n20458 = ~n5439 ;
  assign n5441 = n20458 & n5440 ;
  assign n20459 = ~n5441 ;
  assign n5442 = n5436 & n20459 ;
  assign n5443 = n5435 | n5442 ;
  assign n5444 = x93 & n5443 ;
  assign n5445 = x93 | n5443 ;
  assign n5446 = n5137 & n20371 ;
  assign n5447 = n159 & n5446 ;
  assign n5448 = n5143 & n5447 ;
  assign n5449 = n5143 | n5447 ;
  assign n20460 = ~n5448 ;
  assign n5450 = n20460 & n5449 ;
  assign n20461 = ~n5450 ;
  assign n5451 = n5445 & n20461 ;
  assign n5452 = n5444 | n5451 ;
  assign n5453 = x94 & n5452 ;
  assign n5454 = x94 | n5452 ;
  assign n5455 = n5146 & n20375 ;
  assign n5456 = n159 & n5455 ;
  assign n5457 = n5152 & n5456 ;
  assign n5458 = n5152 | n5456 ;
  assign n20462 = ~n5457 ;
  assign n5459 = n20462 & n5458 ;
  assign n20463 = ~n5459 ;
  assign n5460 = n5454 & n20463 ;
  assign n5461 = n5453 | n5460 ;
  assign n5462 = x95 & n5461 ;
  assign n5463 = x95 | n5461 ;
  assign n5464 = n5155 & n20379 ;
  assign n5465 = n159 & n5464 ;
  assign n5466 = n5161 & n5465 ;
  assign n5467 = n5161 | n5465 ;
  assign n20464 = ~n5466 ;
  assign n5468 = n20464 & n5467 ;
  assign n20465 = ~n5468 ;
  assign n5469 = n5463 & n20465 ;
  assign n5470 = n5462 | n5469 ;
  assign n5471 = x96 & n5470 ;
  assign n5472 = x96 | n5470 ;
  assign n5473 = n5164 & n20383 ;
  assign n5474 = n159 & n5473 ;
  assign n5475 = n5170 & n5474 ;
  assign n5476 = n5170 | n5474 ;
  assign n20466 = ~n5475 ;
  assign n5477 = n20466 & n5476 ;
  assign n20467 = ~n5477 ;
  assign n5478 = n5472 & n20467 ;
  assign n5479 = n5471 | n5478 ;
  assign n5481 = x97 & n5479 ;
  assign n20468 = ~n5481 ;
  assign n5482 = n5192 & n20468 ;
  assign n5182 = n21884 | n5179 ;
  assign n5183 = n5181 & n5182 ;
  assign n20469 = ~x98 ;
  assign n5184 = n20469 & n5183 ;
  assign n5480 = x97 | n5479 ;
  assign n20470 = ~n5184 ;
  assign n5483 = n20470 & n5480 ;
  assign n20471 = ~n5482 ;
  assign n5484 = n20471 & n5483 ;
  assign n5485 = n18403 | n5484 ;
  assign n20472 = ~n5183 ;
  assign n5487 = x98 & n20472 ;
  assign n5488 = n5485 | n5487 ;
  assign n5502 = n5480 & n20468 ;
  assign n158 = ~n5488 ;
  assign n5503 = n158 & n5502 ;
  assign n20474 = ~n5192 ;
  assign n5504 = n20474 & n5503 ;
  assign n20475 = ~n5503 ;
  assign n5505 = n5192 & n20475 ;
  assign n5506 = n5504 | n5505 ;
  assign n5486 = n21884 | n5485 ;
  assign n5507 = n5183 & n5486 ;
  assign n20476 = ~n5507 ;
  assign n5509 = x99 & n20476 ;
  assign n20477 = ~x28 ;
  assign n5510 = n20477 & x64 ;
  assign n5512 = x65 | n5510 ;
  assign n5511 = x65 & n5510 ;
  assign n5513 = x64 & n158 ;
  assign n5514 = x29 & n5513 ;
  assign n5515 = x29 | n5513 ;
  assign n20478 = ~n5514 ;
  assign n5516 = n20478 & n5515 ;
  assign n20479 = ~n5511 ;
  assign n5517 = n20479 & n5516 ;
  assign n20480 = ~n5517 ;
  assign n5518 = n5512 & n20480 ;
  assign n5519 = x66 & n5518 ;
  assign n5520 = x66 | n5518 ;
  assign n5521 = n20393 & n5195 ;
  assign n5522 = n158 & n5521 ;
  assign n5523 = n5199 & n5522 ;
  assign n5524 = n5199 | n5522 ;
  assign n20481 = ~n5523 ;
  assign n5525 = n20481 & n5524 ;
  assign n20482 = ~n5525 ;
  assign n5526 = n5520 & n20482 ;
  assign n5527 = n5519 | n5526 ;
  assign n5528 = x67 & n5527 ;
  assign n5529 = x67 | n5527 ;
  assign n20483 = ~n5202 ;
  assign n5530 = n20483 & n5203 ;
  assign n5531 = n158 & n5530 ;
  assign n5532 = n5208 & n5531 ;
  assign n5533 = n5208 | n5531 ;
  assign n20484 = ~n5532 ;
  assign n5534 = n20484 & n5533 ;
  assign n20485 = ~n5534 ;
  assign n5535 = n5529 & n20485 ;
  assign n5536 = n5528 | n5535 ;
  assign n5537 = x68 & n5536 ;
  assign n5538 = x68 | n5536 ;
  assign n5539 = n5211 | n5488 ;
  assign n20486 = ~n5539 ;
  assign n5540 = n5216 & n20486 ;
  assign n20487 = ~n5540 ;
  assign n5541 = n5215 & n20487 ;
  assign n5542 = n5217 & n20486 ;
  assign n5543 = n5541 | n5542 ;
  assign n20488 = ~n5543 ;
  assign n5544 = n5538 & n20488 ;
  assign n5545 = n5537 | n5544 ;
  assign n5546 = x69 & n5545 ;
  assign n5547 = x69 | n5545 ;
  assign n20489 = ~n5219 ;
  assign n5548 = n20489 & n5220 ;
  assign n5549 = n158 & n5548 ;
  assign n5550 = n20400 & n5549 ;
  assign n20490 = ~n5549 ;
  assign n5551 = n5225 & n20490 ;
  assign n5552 = n5550 | n5551 ;
  assign n20491 = ~n5552 ;
  assign n5553 = n5547 & n20491 ;
  assign n5554 = n5546 | n5553 ;
  assign n5555 = x70 & n5554 ;
  assign n5556 = x70 | n5554 ;
  assign n20492 = ~n5228 ;
  assign n5557 = n20492 & n5229 ;
  assign n5558 = n158 & n5557 ;
  assign n5559 = n20403 & n5558 ;
  assign n20493 = ~n5558 ;
  assign n5560 = n5234 & n20493 ;
  assign n5561 = n5559 | n5560 ;
  assign n20494 = ~n5561 ;
  assign n5562 = n5556 & n20494 ;
  assign n5563 = n5555 | n5562 ;
  assign n5564 = x71 & n5563 ;
  assign n5565 = x71 | n5563 ;
  assign n20495 = ~n5237 ;
  assign n5566 = n20495 & n5238 ;
  assign n5567 = n158 & n5566 ;
  assign n5568 = n5243 & n5567 ;
  assign n5569 = n5243 | n5567 ;
  assign n20496 = ~n5568 ;
  assign n5570 = n20496 & n5569 ;
  assign n20497 = ~n5570 ;
  assign n5571 = n5565 & n20497 ;
  assign n5572 = n5564 | n5571 ;
  assign n5573 = x72 & n5572 ;
  assign n5574 = x72 | n5572 ;
  assign n20498 = ~n5246 ;
  assign n5575 = n20498 & n5247 ;
  assign n5576 = n158 & n5575 ;
  assign n5577 = n5252 & n5576 ;
  assign n5578 = n5252 | n5576 ;
  assign n20499 = ~n5577 ;
  assign n5579 = n20499 & n5578 ;
  assign n20500 = ~n5579 ;
  assign n5580 = n5574 & n20500 ;
  assign n5581 = n5573 | n5580 ;
  assign n5582 = x73 & n5581 ;
  assign n5583 = x73 | n5581 ;
  assign n20501 = ~n5255 ;
  assign n5584 = n20501 & n5256 ;
  assign n5585 = n158 & n5584 ;
  assign n5586 = n20410 & n5585 ;
  assign n20502 = ~n5585 ;
  assign n5587 = n5261 & n20502 ;
  assign n5588 = n5586 | n5587 ;
  assign n20503 = ~n5588 ;
  assign n5589 = n5583 & n20503 ;
  assign n5590 = n5582 | n5589 ;
  assign n5591 = x74 & n5590 ;
  assign n5592 = x74 | n5590 ;
  assign n20504 = ~n5264 ;
  assign n5593 = n20504 & n5265 ;
  assign n5594 = n158 & n5593 ;
  assign n5595 = n20413 & n5594 ;
  assign n20505 = ~n5594 ;
  assign n5596 = n5270 & n20505 ;
  assign n5597 = n5595 | n5596 ;
  assign n20506 = ~n5597 ;
  assign n5598 = n5592 & n20506 ;
  assign n5599 = n5591 | n5598 ;
  assign n5600 = x75 & n5599 ;
  assign n5601 = x75 | n5599 ;
  assign n20507 = ~n5273 ;
  assign n5602 = n20507 & n5274 ;
  assign n5603 = n158 & n5602 ;
  assign n5604 = n20416 & n5603 ;
  assign n20508 = ~n5603 ;
  assign n5605 = n5279 & n20508 ;
  assign n5606 = n5604 | n5605 ;
  assign n20509 = ~n5606 ;
  assign n5607 = n5601 & n20509 ;
  assign n5608 = n5600 | n5607 ;
  assign n5609 = x76 & n5608 ;
  assign n5610 = x76 | n5608 ;
  assign n20510 = ~n5282 ;
  assign n5611 = n20510 & n5283 ;
  assign n5612 = n158 & n5611 ;
  assign n5613 = n5288 & n5612 ;
  assign n5614 = n5288 | n5612 ;
  assign n20511 = ~n5613 ;
  assign n5615 = n20511 & n5614 ;
  assign n20512 = ~n5615 ;
  assign n5616 = n5610 & n20512 ;
  assign n5617 = n5609 | n5616 ;
  assign n5618 = x77 & n5617 ;
  assign n5619 = x77 | n5617 ;
  assign n20513 = ~n5291 ;
  assign n5620 = n20513 & n5292 ;
  assign n5621 = n158 & n5620 ;
  assign n5622 = n20422 & n5621 ;
  assign n20514 = ~n5621 ;
  assign n5623 = n5297 & n20514 ;
  assign n5624 = n5622 | n5623 ;
  assign n20515 = ~n5624 ;
  assign n5625 = n5619 & n20515 ;
  assign n5626 = n5618 | n5625 ;
  assign n5627 = x78 & n5626 ;
  assign n5628 = x78 | n5626 ;
  assign n20516 = ~n5300 ;
  assign n5629 = n20516 & n5301 ;
  assign n5630 = n158 & n5629 ;
  assign n5631 = n5306 & n5630 ;
  assign n5632 = n5306 | n5630 ;
  assign n20517 = ~n5631 ;
  assign n5633 = n20517 & n5632 ;
  assign n20518 = ~n5633 ;
  assign n5634 = n5628 & n20518 ;
  assign n5635 = n5627 | n5634 ;
  assign n5636 = x79 & n5635 ;
  assign n5637 = x79 | n5635 ;
  assign n20519 = ~n5309 ;
  assign n5638 = n20519 & n5310 ;
  assign n5639 = n158 & n5638 ;
  assign n5640 = n5315 & n5639 ;
  assign n5641 = n5315 | n5639 ;
  assign n20520 = ~n5640 ;
  assign n5642 = n20520 & n5641 ;
  assign n20521 = ~n5642 ;
  assign n5643 = n5637 & n20521 ;
  assign n5644 = n5636 | n5643 ;
  assign n5645 = x80 & n5644 ;
  assign n5646 = x80 | n5644 ;
  assign n20522 = ~n5318 ;
  assign n5647 = n20522 & n5319 ;
  assign n5648 = n158 & n5647 ;
  assign n5649 = n5324 & n5648 ;
  assign n5650 = n5324 | n5648 ;
  assign n20523 = ~n5649 ;
  assign n5651 = n20523 & n5650 ;
  assign n20524 = ~n5651 ;
  assign n5652 = n5646 & n20524 ;
  assign n5653 = n5645 | n5652 ;
  assign n5654 = x81 & n5653 ;
  assign n5655 = x81 | n5653 ;
  assign n20525 = ~n5327 ;
  assign n5656 = n20525 & n5328 ;
  assign n5657 = n158 & n5656 ;
  assign n5658 = n20431 & n5657 ;
  assign n20526 = ~n5657 ;
  assign n5659 = n5333 & n20526 ;
  assign n5660 = n5658 | n5659 ;
  assign n20527 = ~n5660 ;
  assign n5661 = n5655 & n20527 ;
  assign n5662 = n5654 | n5661 ;
  assign n5663 = x82 & n5662 ;
  assign n5664 = x82 | n5662 ;
  assign n20528 = ~n5336 ;
  assign n5665 = n20528 & n5337 ;
  assign n5666 = n158 & n5665 ;
  assign n5667 = n20434 & n5666 ;
  assign n20529 = ~n5666 ;
  assign n5668 = n5342 & n20529 ;
  assign n5669 = n5667 | n5668 ;
  assign n20530 = ~n5669 ;
  assign n5670 = n5664 & n20530 ;
  assign n5671 = n5663 | n5670 ;
  assign n5672 = x83 & n5671 ;
  assign n5673 = x83 | n5671 ;
  assign n20531 = ~n5345 ;
  assign n5674 = n20531 & n5346 ;
  assign n5675 = n158 & n5674 ;
  assign n5676 = n5351 & n5675 ;
  assign n5677 = n5351 | n5675 ;
  assign n20532 = ~n5676 ;
  assign n5678 = n20532 & n5677 ;
  assign n20533 = ~n5678 ;
  assign n5679 = n5673 & n20533 ;
  assign n5680 = n5672 | n5679 ;
  assign n5681 = x84 & n5680 ;
  assign n5682 = x84 | n5680 ;
  assign n20534 = ~n5354 ;
  assign n5683 = n20534 & n5355 ;
  assign n5684 = n158 & n5683 ;
  assign n5685 = n5360 & n5684 ;
  assign n5686 = n5360 | n5684 ;
  assign n20535 = ~n5685 ;
  assign n5687 = n20535 & n5686 ;
  assign n20536 = ~n5687 ;
  assign n5688 = n5682 & n20536 ;
  assign n5689 = n5681 | n5688 ;
  assign n5690 = x85 & n5689 ;
  assign n5691 = x85 | n5689 ;
  assign n20537 = ~n5363 ;
  assign n5692 = n20537 & n5364 ;
  assign n5693 = n158 & n5692 ;
  assign n5694 = n5369 & n5693 ;
  assign n5695 = n5369 | n5693 ;
  assign n20538 = ~n5694 ;
  assign n5696 = n20538 & n5695 ;
  assign n20539 = ~n5696 ;
  assign n5697 = n5691 & n20539 ;
  assign n5698 = n5690 | n5697 ;
  assign n5699 = x86 & n5698 ;
  assign n5700 = x86 | n5698 ;
  assign n20540 = ~n5372 ;
  assign n5701 = n20540 & n5373 ;
  assign n5702 = n158 & n5701 ;
  assign n5703 = n5378 & n5702 ;
  assign n5704 = n5378 | n5702 ;
  assign n20541 = ~n5703 ;
  assign n5705 = n20541 & n5704 ;
  assign n20542 = ~n5705 ;
  assign n5706 = n5700 & n20542 ;
  assign n5707 = n5699 | n5706 ;
  assign n5708 = x87 & n5707 ;
  assign n5709 = x87 | n5707 ;
  assign n20543 = ~n5381 ;
  assign n5710 = n20543 & n5382 ;
  assign n5711 = n158 & n5710 ;
  assign n5712 = n5387 & n5711 ;
  assign n5713 = n5387 | n5711 ;
  assign n20544 = ~n5712 ;
  assign n5714 = n20544 & n5713 ;
  assign n20545 = ~n5714 ;
  assign n5715 = n5709 & n20545 ;
  assign n5716 = n5708 | n5715 ;
  assign n5717 = x88 & n5716 ;
  assign n5718 = x88 | n5716 ;
  assign n20546 = ~n5390 ;
  assign n5719 = n20546 & n5391 ;
  assign n5720 = n158 & n5719 ;
  assign n5721 = n5396 & n5720 ;
  assign n5722 = n5396 | n5720 ;
  assign n20547 = ~n5721 ;
  assign n5723 = n20547 & n5722 ;
  assign n20548 = ~n5723 ;
  assign n5724 = n5718 & n20548 ;
  assign n5725 = n5717 | n5724 ;
  assign n5726 = x89 & n5725 ;
  assign n5727 = x89 | n5725 ;
  assign n20549 = ~n5399 ;
  assign n5728 = n20549 & n5400 ;
  assign n5729 = n158 & n5728 ;
  assign n5730 = n5405 & n5729 ;
  assign n5731 = n5405 | n5729 ;
  assign n20550 = ~n5730 ;
  assign n5732 = n20550 & n5731 ;
  assign n20551 = ~n5732 ;
  assign n5733 = n5727 & n20551 ;
  assign n5734 = n5726 | n5733 ;
  assign n5735 = x90 & n5734 ;
  assign n5736 = x90 | n5734 ;
  assign n20552 = ~n5408 ;
  assign n5737 = n20552 & n5409 ;
  assign n5738 = n158 & n5737 ;
  assign n5739 = n5414 & n5738 ;
  assign n5740 = n5414 | n5738 ;
  assign n20553 = ~n5739 ;
  assign n5741 = n20553 & n5740 ;
  assign n20554 = ~n5741 ;
  assign n5742 = n5736 & n20554 ;
  assign n5743 = n5735 | n5742 ;
  assign n5744 = x91 & n5743 ;
  assign n5745 = x91 | n5743 ;
  assign n20555 = ~n5417 ;
  assign n5746 = n20555 & n5418 ;
  assign n5747 = n158 & n5746 ;
  assign n5748 = n20454 & n5747 ;
  assign n20556 = ~n5747 ;
  assign n5749 = n5423 & n20556 ;
  assign n5750 = n5748 | n5749 ;
  assign n20557 = ~n5750 ;
  assign n5751 = n5745 & n20557 ;
  assign n5752 = n5744 | n5751 ;
  assign n5753 = x92 & n5752 ;
  assign n5754 = x92 | n5752 ;
  assign n20558 = ~n5426 ;
  assign n5755 = n20558 & n5427 ;
  assign n5756 = n158 & n5755 ;
  assign n5757 = n20457 & n5756 ;
  assign n20559 = ~n5756 ;
  assign n5758 = n5432 & n20559 ;
  assign n5759 = n5757 | n5758 ;
  assign n20560 = ~n5759 ;
  assign n5760 = n5754 & n20560 ;
  assign n5761 = n5753 | n5760 ;
  assign n5762 = x93 & n5761 ;
  assign n5763 = x93 | n5761 ;
  assign n20561 = ~n5435 ;
  assign n5764 = n20561 & n5436 ;
  assign n5765 = n158 & n5764 ;
  assign n5766 = n5441 & n5765 ;
  assign n5767 = n5441 | n5765 ;
  assign n20562 = ~n5766 ;
  assign n5768 = n20562 & n5767 ;
  assign n20563 = ~n5768 ;
  assign n5769 = n5763 & n20563 ;
  assign n5770 = n5762 | n5769 ;
  assign n5771 = x94 & n5770 ;
  assign n5772 = x94 | n5770 ;
  assign n20564 = ~n5444 ;
  assign n5773 = n20564 & n5445 ;
  assign n5774 = n158 & n5773 ;
  assign n5775 = n5450 & n5774 ;
  assign n5776 = n5450 | n5774 ;
  assign n20565 = ~n5775 ;
  assign n5777 = n20565 & n5776 ;
  assign n20566 = ~n5777 ;
  assign n5778 = n5772 & n20566 ;
  assign n5779 = n5771 | n5778 ;
  assign n5780 = x95 & n5779 ;
  assign n5781 = x95 | n5779 ;
  assign n20567 = ~n5453 ;
  assign n5782 = n20567 & n5454 ;
  assign n5783 = n158 & n5782 ;
  assign n5784 = n5459 & n5783 ;
  assign n5785 = n5459 | n5783 ;
  assign n20568 = ~n5784 ;
  assign n5786 = n20568 & n5785 ;
  assign n20569 = ~n5786 ;
  assign n5787 = n5781 & n20569 ;
  assign n5788 = n5780 | n5787 ;
  assign n5789 = x96 & n5788 ;
  assign n5790 = x96 | n5788 ;
  assign n20570 = ~n5462 ;
  assign n5791 = n20570 & n5463 ;
  assign n5792 = n158 & n5791 ;
  assign n5793 = n5468 & n5792 ;
  assign n5794 = n5468 | n5792 ;
  assign n20571 = ~n5793 ;
  assign n5795 = n20571 & n5794 ;
  assign n20572 = ~n5795 ;
  assign n5796 = n5790 & n20572 ;
  assign n5797 = n5789 | n5796 ;
  assign n5798 = x97 & n5797 ;
  assign n5799 = x97 | n5797 ;
  assign n20573 = ~n5471 ;
  assign n5800 = n20573 & n5472 ;
  assign n5801 = n158 & n5800 ;
  assign n5802 = n5477 & n5801 ;
  assign n5803 = n5477 | n5801 ;
  assign n20574 = ~n5802 ;
  assign n5804 = n20574 & n5803 ;
  assign n20575 = ~n5804 ;
  assign n5805 = n5799 & n20575 ;
  assign n5806 = n5798 | n5805 ;
  assign n5809 = x98 & n5806 ;
  assign n20576 = ~n5809 ;
  assign n5810 = n5506 & n20576 ;
  assign n20577 = ~x99 ;
  assign n5508 = n20577 & n5507 ;
  assign n5807 = x98 | n5806 ;
  assign n20578 = ~n5508 ;
  assign n5811 = n20578 & n5807 ;
  assign n20579 = ~n5810 ;
  assign n5812 = n20579 & n5811 ;
  assign n5813 = n18398 | n5812 ;
  assign n5814 = n5509 | n5813 ;
  assign n20580 = ~n5806 ;
  assign n5808 = x98 & n20580 ;
  assign n5815 = n20469 & n5806 ;
  assign n5816 = n5808 | n5815 ;
  assign n157 = ~n5814 ;
  assign n5817 = n157 & n5816 ;
  assign n20582 = ~n5506 ;
  assign n5818 = n20582 & n5817 ;
  assign n20583 = ~n5817 ;
  assign n5819 = n5506 & n20583 ;
  assign n5820 = n5818 | n5819 ;
  assign n20584 = ~x27 ;
  assign n5821 = n20584 & x64 ;
  assign n5823 = x65 | n5821 ;
  assign n5822 = x65 & n5821 ;
  assign n5824 = x64 & n157 ;
  assign n5825 = x28 & n5824 ;
  assign n5826 = x28 | n5824 ;
  assign n20585 = ~n5825 ;
  assign n5827 = n20585 & n5826 ;
  assign n20586 = ~n5822 ;
  assign n5828 = n20586 & n5827 ;
  assign n20587 = ~n5828 ;
  assign n5829 = n5823 & n20587 ;
  assign n5830 = x66 & n5829 ;
  assign n5831 = x66 | n5829 ;
  assign n5832 = n20479 & n5512 ;
  assign n5833 = n157 & n5832 ;
  assign n5834 = n5516 & n5833 ;
  assign n5835 = n5516 | n5833 ;
  assign n20588 = ~n5834 ;
  assign n5836 = n20588 & n5835 ;
  assign n20589 = ~n5836 ;
  assign n5837 = n5831 & n20589 ;
  assign n5838 = n5830 | n5837 ;
  assign n5839 = x67 & n5838 ;
  assign n5840 = x67 | n5838 ;
  assign n20590 = ~n5519 ;
  assign n5841 = n20590 & n5520 ;
  assign n5842 = n157 & n5841 ;
  assign n5843 = n5525 & n5842 ;
  assign n5844 = n5525 | n5842 ;
  assign n20591 = ~n5843 ;
  assign n5845 = n20591 & n5844 ;
  assign n20592 = ~n5845 ;
  assign n5846 = n5840 & n20592 ;
  assign n5847 = n5839 | n5846 ;
  assign n5848 = x68 & n5847 ;
  assign n5849 = x68 | n5847 ;
  assign n20593 = ~n5528 ;
  assign n5850 = n20593 & n5529 ;
  assign n5851 = n157 & n5850 ;
  assign n5852 = n5534 & n5851 ;
  assign n5853 = n5534 | n5851 ;
  assign n20594 = ~n5852 ;
  assign n5854 = n20594 & n5853 ;
  assign n20595 = ~n5854 ;
  assign n5855 = n5849 & n20595 ;
  assign n5856 = n5848 | n5855 ;
  assign n5857 = x69 & n5856 ;
  assign n5858 = x69 | n5856 ;
  assign n20596 = ~n5537 ;
  assign n5859 = n20596 & n5538 ;
  assign n5860 = n157 & n5859 ;
  assign n5861 = n5543 & n5860 ;
  assign n5862 = n5543 | n5860 ;
  assign n20597 = ~n5861 ;
  assign n5863 = n20597 & n5862 ;
  assign n20598 = ~n5863 ;
  assign n5864 = n5858 & n20598 ;
  assign n5865 = n5857 | n5864 ;
  assign n5866 = x70 & n5865 ;
  assign n5867 = x70 | n5865 ;
  assign n20599 = ~n5546 ;
  assign n5868 = n20599 & n5547 ;
  assign n5869 = n157 & n5868 ;
  assign n5870 = n20491 & n5869 ;
  assign n20600 = ~n5869 ;
  assign n5871 = n5552 & n20600 ;
  assign n5872 = n5870 | n5871 ;
  assign n20601 = ~n5872 ;
  assign n5873 = n5867 & n20601 ;
  assign n5874 = n5866 | n5873 ;
  assign n5875 = x71 & n5874 ;
  assign n5876 = x71 | n5874 ;
  assign n20602 = ~n5555 ;
  assign n5877 = n20602 & n5556 ;
  assign n5878 = n157 & n5877 ;
  assign n5879 = n20494 & n5878 ;
  assign n20603 = ~n5878 ;
  assign n5880 = n5561 & n20603 ;
  assign n5881 = n5879 | n5880 ;
  assign n20604 = ~n5881 ;
  assign n5882 = n5876 & n20604 ;
  assign n5883 = n5875 | n5882 ;
  assign n5884 = x72 & n5883 ;
  assign n5885 = x72 | n5883 ;
  assign n20605 = ~n5564 ;
  assign n5886 = n20605 & n5565 ;
  assign n5887 = n157 & n5886 ;
  assign n5888 = n5570 & n5887 ;
  assign n5889 = n5570 | n5887 ;
  assign n20606 = ~n5888 ;
  assign n5890 = n20606 & n5889 ;
  assign n20607 = ~n5890 ;
  assign n5891 = n5885 & n20607 ;
  assign n5892 = n5884 | n5891 ;
  assign n5893 = x73 & n5892 ;
  assign n5894 = x73 | n5892 ;
  assign n20608 = ~n5573 ;
  assign n5895 = n20608 & n5574 ;
  assign n5896 = n157 & n5895 ;
  assign n5897 = n20500 & n5896 ;
  assign n20609 = ~n5896 ;
  assign n5898 = n5579 & n20609 ;
  assign n5899 = n5897 | n5898 ;
  assign n20610 = ~n5899 ;
  assign n5900 = n5894 & n20610 ;
  assign n5901 = n5893 | n5900 ;
  assign n5902 = x74 & n5901 ;
  assign n5903 = x74 | n5901 ;
  assign n20611 = ~n5582 ;
  assign n5904 = n20611 & n5583 ;
  assign n5905 = n157 & n5904 ;
  assign n5906 = n20503 & n5905 ;
  assign n20612 = ~n5905 ;
  assign n5907 = n5588 & n20612 ;
  assign n5908 = n5906 | n5907 ;
  assign n20613 = ~n5908 ;
  assign n5909 = n5903 & n20613 ;
  assign n5910 = n5902 | n5909 ;
  assign n5911 = x75 & n5910 ;
  assign n5912 = x75 | n5910 ;
  assign n20614 = ~n5591 ;
  assign n5913 = n20614 & n5592 ;
  assign n5914 = n157 & n5913 ;
  assign n5915 = n20506 & n5914 ;
  assign n20615 = ~n5914 ;
  assign n5916 = n5597 & n20615 ;
  assign n5917 = n5915 | n5916 ;
  assign n20616 = ~n5917 ;
  assign n5918 = n5912 & n20616 ;
  assign n5919 = n5911 | n5918 ;
  assign n5920 = x76 & n5919 ;
  assign n5921 = x76 | n5919 ;
  assign n20617 = ~n5600 ;
  assign n5922 = n20617 & n5601 ;
  assign n5923 = n157 & n5922 ;
  assign n5924 = n20509 & n5923 ;
  assign n20618 = ~n5923 ;
  assign n5925 = n5606 & n20618 ;
  assign n5926 = n5924 | n5925 ;
  assign n20619 = ~n5926 ;
  assign n5927 = n5921 & n20619 ;
  assign n5928 = n5920 | n5927 ;
  assign n5929 = x77 & n5928 ;
  assign n5930 = x77 | n5928 ;
  assign n20620 = ~n5609 ;
  assign n5931 = n20620 & n5610 ;
  assign n5932 = n157 & n5931 ;
  assign n5933 = n5615 & n5932 ;
  assign n5934 = n5615 | n5932 ;
  assign n20621 = ~n5933 ;
  assign n5935 = n20621 & n5934 ;
  assign n20622 = ~n5935 ;
  assign n5936 = n5930 & n20622 ;
  assign n5937 = n5929 | n5936 ;
  assign n5938 = x78 & n5937 ;
  assign n5939 = x78 | n5937 ;
  assign n20623 = ~n5618 ;
  assign n5940 = n20623 & n5619 ;
  assign n5941 = n157 & n5940 ;
  assign n5942 = n5624 & n5941 ;
  assign n5943 = n5624 | n5941 ;
  assign n20624 = ~n5942 ;
  assign n5944 = n20624 & n5943 ;
  assign n20625 = ~n5944 ;
  assign n5945 = n5939 & n20625 ;
  assign n5946 = n5938 | n5945 ;
  assign n5947 = x79 & n5946 ;
  assign n5948 = x79 | n5946 ;
  assign n20626 = ~n5627 ;
  assign n5949 = n20626 & n5628 ;
  assign n5950 = n157 & n5949 ;
  assign n5951 = n5633 & n5950 ;
  assign n5952 = n5633 | n5950 ;
  assign n20627 = ~n5951 ;
  assign n5953 = n20627 & n5952 ;
  assign n20628 = ~n5953 ;
  assign n5954 = n5948 & n20628 ;
  assign n5955 = n5947 | n5954 ;
  assign n5956 = x80 & n5955 ;
  assign n5957 = x80 | n5955 ;
  assign n20629 = ~n5636 ;
  assign n5958 = n20629 & n5637 ;
  assign n5959 = n157 & n5958 ;
  assign n5960 = n20521 & n5959 ;
  assign n20630 = ~n5959 ;
  assign n5961 = n5642 & n20630 ;
  assign n5962 = n5960 | n5961 ;
  assign n20631 = ~n5962 ;
  assign n5963 = n5957 & n20631 ;
  assign n5964 = n5956 | n5963 ;
  assign n5965 = x81 & n5964 ;
  assign n5966 = x81 | n5964 ;
  assign n20632 = ~n5645 ;
  assign n5967 = n20632 & n5646 ;
  assign n5968 = n157 & n5967 ;
  assign n5969 = n20524 & n5968 ;
  assign n20633 = ~n5968 ;
  assign n5970 = n5651 & n20633 ;
  assign n5971 = n5969 | n5970 ;
  assign n20634 = ~n5971 ;
  assign n5972 = n5966 & n20634 ;
  assign n5973 = n5965 | n5972 ;
  assign n5974 = x82 & n5973 ;
  assign n5975 = x82 | n5973 ;
  assign n20635 = ~n5654 ;
  assign n5976 = n20635 & n5655 ;
  assign n5977 = n157 & n5976 ;
  assign n5978 = n20527 & n5977 ;
  assign n20636 = ~n5977 ;
  assign n5979 = n5660 & n20636 ;
  assign n5980 = n5978 | n5979 ;
  assign n20637 = ~n5980 ;
  assign n5981 = n5975 & n20637 ;
  assign n5982 = n5974 | n5981 ;
  assign n5983 = x83 & n5982 ;
  assign n5984 = x83 | n5982 ;
  assign n20638 = ~n5663 ;
  assign n5985 = n20638 & n5664 ;
  assign n5986 = n157 & n5985 ;
  assign n5987 = n5669 & n5986 ;
  assign n5988 = n5669 | n5986 ;
  assign n20639 = ~n5987 ;
  assign n5989 = n20639 & n5988 ;
  assign n20640 = ~n5989 ;
  assign n5990 = n5984 & n20640 ;
  assign n5991 = n5983 | n5990 ;
  assign n5992 = x84 & n5991 ;
  assign n5993 = x84 | n5991 ;
  assign n20641 = ~n5672 ;
  assign n5994 = n20641 & n5673 ;
  assign n5995 = n157 & n5994 ;
  assign n5996 = n5678 & n5995 ;
  assign n5997 = n5678 | n5995 ;
  assign n20642 = ~n5996 ;
  assign n5998 = n20642 & n5997 ;
  assign n20643 = ~n5998 ;
  assign n5999 = n5993 & n20643 ;
  assign n6000 = n5992 | n5999 ;
  assign n6001 = x85 & n6000 ;
  assign n6002 = x85 | n6000 ;
  assign n20644 = ~n5681 ;
  assign n6003 = n20644 & n5682 ;
  assign n6004 = n157 & n6003 ;
  assign n6005 = n5687 & n6004 ;
  assign n6006 = n5687 | n6004 ;
  assign n20645 = ~n6005 ;
  assign n6007 = n20645 & n6006 ;
  assign n20646 = ~n6007 ;
  assign n6008 = n6002 & n20646 ;
  assign n6009 = n6001 | n6008 ;
  assign n6010 = x86 & n6009 ;
  assign n6011 = x86 | n6009 ;
  assign n20647 = ~n5690 ;
  assign n6012 = n20647 & n5691 ;
  assign n6013 = n157 & n6012 ;
  assign n6014 = n5696 & n6013 ;
  assign n6015 = n5696 | n6013 ;
  assign n20648 = ~n6014 ;
  assign n6016 = n20648 & n6015 ;
  assign n20649 = ~n6016 ;
  assign n6017 = n6011 & n20649 ;
  assign n6018 = n6010 | n6017 ;
  assign n6019 = x87 & n6018 ;
  assign n6020 = x87 | n6018 ;
  assign n20650 = ~n5699 ;
  assign n6021 = n20650 & n5700 ;
  assign n6022 = n157 & n6021 ;
  assign n6023 = n5705 & n6022 ;
  assign n6024 = n5705 | n6022 ;
  assign n20651 = ~n6023 ;
  assign n6025 = n20651 & n6024 ;
  assign n20652 = ~n6025 ;
  assign n6026 = n6020 & n20652 ;
  assign n6027 = n6019 | n6026 ;
  assign n6028 = x88 & n6027 ;
  assign n6029 = x88 | n6027 ;
  assign n20653 = ~n5708 ;
  assign n6030 = n20653 & n5709 ;
  assign n6031 = n157 & n6030 ;
  assign n6032 = n5714 & n6031 ;
  assign n6033 = n5714 | n6031 ;
  assign n20654 = ~n6032 ;
  assign n6034 = n20654 & n6033 ;
  assign n20655 = ~n6034 ;
  assign n6035 = n6029 & n20655 ;
  assign n6036 = n6028 | n6035 ;
  assign n6037 = x89 & n6036 ;
  assign n6038 = x89 | n6036 ;
  assign n20656 = ~n5717 ;
  assign n6039 = n20656 & n5718 ;
  assign n6040 = n157 & n6039 ;
  assign n6041 = n5723 & n6040 ;
  assign n6042 = n5723 | n6040 ;
  assign n20657 = ~n6041 ;
  assign n6043 = n20657 & n6042 ;
  assign n20658 = ~n6043 ;
  assign n6044 = n6038 & n20658 ;
  assign n6045 = n6037 | n6044 ;
  assign n6046 = x90 & n6045 ;
  assign n6047 = x90 | n6045 ;
  assign n20659 = ~n5726 ;
  assign n6048 = n20659 & n5727 ;
  assign n6049 = n157 & n6048 ;
  assign n6050 = n5732 & n6049 ;
  assign n6051 = n5732 | n6049 ;
  assign n20660 = ~n6050 ;
  assign n6052 = n20660 & n6051 ;
  assign n20661 = ~n6052 ;
  assign n6053 = n6047 & n20661 ;
  assign n6054 = n6046 | n6053 ;
  assign n6055 = x91 & n6054 ;
  assign n6056 = x91 | n6054 ;
  assign n20662 = ~n5735 ;
  assign n6057 = n20662 & n5736 ;
  assign n6058 = n157 & n6057 ;
  assign n6059 = n5741 & n6058 ;
  assign n6060 = n5741 | n6058 ;
  assign n20663 = ~n6059 ;
  assign n6061 = n20663 & n6060 ;
  assign n20664 = ~n6061 ;
  assign n6062 = n6056 & n20664 ;
  assign n6063 = n6055 | n6062 ;
  assign n6064 = x92 & n6063 ;
  assign n6065 = x92 | n6063 ;
  assign n20665 = ~n5744 ;
  assign n6066 = n20665 & n5745 ;
  assign n6067 = n157 & n6066 ;
  assign n6068 = n20557 & n6067 ;
  assign n20666 = ~n6067 ;
  assign n6069 = n5750 & n20666 ;
  assign n6070 = n6068 | n6069 ;
  assign n20667 = ~n6070 ;
  assign n6071 = n6065 & n20667 ;
  assign n6072 = n6064 | n6071 ;
  assign n6073 = x93 & n6072 ;
  assign n6074 = x93 | n6072 ;
  assign n20668 = ~n5753 ;
  assign n6075 = n20668 & n5754 ;
  assign n6076 = n157 & n6075 ;
  assign n6077 = n20560 & n6076 ;
  assign n20669 = ~n6076 ;
  assign n6078 = n5759 & n20669 ;
  assign n6079 = n6077 | n6078 ;
  assign n20670 = ~n6079 ;
  assign n6080 = n6074 & n20670 ;
  assign n6081 = n6073 | n6080 ;
  assign n6082 = x94 & n6081 ;
  assign n6083 = x94 | n6081 ;
  assign n20671 = ~n5762 ;
  assign n6084 = n20671 & n5763 ;
  assign n6085 = n157 & n6084 ;
  assign n6086 = n5768 & n6085 ;
  assign n6087 = n5768 | n6085 ;
  assign n20672 = ~n6086 ;
  assign n6088 = n20672 & n6087 ;
  assign n20673 = ~n6088 ;
  assign n6089 = n6083 & n20673 ;
  assign n6090 = n6082 | n6089 ;
  assign n6091 = x95 & n6090 ;
  assign n6092 = x95 | n6090 ;
  assign n20674 = ~n5771 ;
  assign n6093 = n20674 & n5772 ;
  assign n6094 = n157 & n6093 ;
  assign n6095 = n5777 & n6094 ;
  assign n6096 = n5777 | n6094 ;
  assign n20675 = ~n6095 ;
  assign n6097 = n20675 & n6096 ;
  assign n20676 = ~n6097 ;
  assign n6098 = n6092 & n20676 ;
  assign n6099 = n6091 | n6098 ;
  assign n6100 = x96 & n6099 ;
  assign n6101 = x96 | n6099 ;
  assign n20677 = ~n5780 ;
  assign n6102 = n20677 & n5781 ;
  assign n6103 = n157 & n6102 ;
  assign n6104 = n5786 & n6103 ;
  assign n6105 = n5786 | n6103 ;
  assign n20678 = ~n6104 ;
  assign n6106 = n20678 & n6105 ;
  assign n20679 = ~n6106 ;
  assign n6107 = n6101 & n20679 ;
  assign n6108 = n6100 | n6107 ;
  assign n6109 = x97 & n6108 ;
  assign n6110 = x97 | n6108 ;
  assign n20680 = ~n5789 ;
  assign n6111 = n20680 & n5790 ;
  assign n6112 = n157 & n6111 ;
  assign n6113 = n5795 & n6112 ;
  assign n6114 = n5795 | n6112 ;
  assign n20681 = ~n6113 ;
  assign n6115 = n20681 & n6114 ;
  assign n20682 = ~n6115 ;
  assign n6116 = n6110 & n20682 ;
  assign n6117 = n6109 | n6116 ;
  assign n6118 = x98 & n6117 ;
  assign n6119 = x98 | n6117 ;
  assign n20683 = ~n5798 ;
  assign n6120 = n20683 & n5799 ;
  assign n6121 = n157 & n6120 ;
  assign n6122 = n20575 & n6121 ;
  assign n20684 = ~n6121 ;
  assign n6123 = n5804 & n20684 ;
  assign n6124 = n6122 | n6123 ;
  assign n20685 = ~n6124 ;
  assign n6125 = n6119 & n20685 ;
  assign n6126 = n6118 | n6125 ;
  assign n6127 = x99 & n6126 ;
  assign n20686 = ~n6127 ;
  assign n6129 = n5820 & n20686 ;
  assign n6128 = x99 | n6126 ;
  assign n20687 = ~n6129 ;
  assign n6130 = n6128 & n20687 ;
  assign n6132 = x100 & n6130 ;
  assign n6133 = n18393 | n6132 ;
  assign n6131 = x100 | n6130 ;
  assign n6134 = n5507 & n5813 ;
  assign n6135 = n21884 | n6134 ;
  assign n20688 = ~n6135 ;
  assign n6136 = n6131 & n20688 ;
  assign n6137 = n6133 | n6136 ;
  assign n156 = ~n6137 ;
  assign n6139 = n6128 & n156 ;
  assign n6140 = n6129 & n6139 ;
  assign n6141 = n20686 & n6139 ;
  assign n6142 = n5820 | n6141 ;
  assign n20690 = ~n6140 ;
  assign n6143 = n20690 & n6142 ;
  assign n6144 = n6133 & n6134 ;
  assign n6145 = n21884 | n6144 ;
  assign n20691 = ~x26 ;
  assign n6146 = n20691 & x64 ;
  assign n6147 = x65 | n6146 ;
  assign n6138 = n5821 & n156 ;
  assign n6148 = x64 & n156 ;
  assign n20692 = ~n6148 ;
  assign n6149 = x27 & n20692 ;
  assign n6150 = n6138 | n6149 ;
  assign n6151 = x65 & n6146 ;
  assign n20693 = ~n6151 ;
  assign n6152 = n6150 & n20693 ;
  assign n20694 = ~n6152 ;
  assign n6153 = n6147 & n20694 ;
  assign n6154 = x66 & n6153 ;
  assign n6155 = n20586 & n5823 ;
  assign n6156 = n156 & n6155 ;
  assign n6157 = n5827 & n6156 ;
  assign n6158 = n5827 | n6156 ;
  assign n20695 = ~n6157 ;
  assign n6159 = n20695 & n6158 ;
  assign n6160 = x66 | n6153 ;
  assign n20696 = ~n6159 ;
  assign n6161 = n20696 & n6160 ;
  assign n6162 = n6154 | n6161 ;
  assign n6163 = x67 & n6162 ;
  assign n6164 = x67 | n6162 ;
  assign n20697 = ~n5830 ;
  assign n6165 = n20697 & n5831 ;
  assign n6166 = n156 & n6165 ;
  assign n6167 = n5836 & n6166 ;
  assign n6168 = n5836 | n6166 ;
  assign n20698 = ~n6167 ;
  assign n6169 = n20698 & n6168 ;
  assign n20699 = ~n6169 ;
  assign n6170 = n6164 & n20699 ;
  assign n6171 = n6163 | n6170 ;
  assign n6172 = x68 & n6171 ;
  assign n6173 = x68 | n6171 ;
  assign n20700 = ~n5839 ;
  assign n6174 = n20700 & n5840 ;
  assign n6175 = n156 & n6174 ;
  assign n6176 = n5845 & n6175 ;
  assign n6177 = n5845 | n6175 ;
  assign n20701 = ~n6176 ;
  assign n6178 = n20701 & n6177 ;
  assign n20702 = ~n6178 ;
  assign n6179 = n6173 & n20702 ;
  assign n6180 = n6172 | n6179 ;
  assign n6181 = x69 & n6180 ;
  assign n6182 = x69 | n6180 ;
  assign n20703 = ~n5848 ;
  assign n6183 = n20703 & n5849 ;
  assign n6184 = n156 & n6183 ;
  assign n6185 = n20595 & n6184 ;
  assign n20704 = ~n6184 ;
  assign n6186 = n5854 & n20704 ;
  assign n6187 = n6185 | n6186 ;
  assign n20705 = ~n6187 ;
  assign n6188 = n6182 & n20705 ;
  assign n6189 = n6181 | n6188 ;
  assign n6190 = x70 & n6189 ;
  assign n6191 = x70 | n6189 ;
  assign n20706 = ~n5857 ;
  assign n6192 = n20706 & n5858 ;
  assign n6193 = n156 & n6192 ;
  assign n6194 = n5863 & n6193 ;
  assign n6195 = n5863 | n6193 ;
  assign n20707 = ~n6194 ;
  assign n6196 = n20707 & n6195 ;
  assign n20708 = ~n6196 ;
  assign n6197 = n6191 & n20708 ;
  assign n6198 = n6190 | n6197 ;
  assign n6199 = x71 & n6198 ;
  assign n6200 = x71 | n6198 ;
  assign n20709 = ~n5866 ;
  assign n6201 = n20709 & n5867 ;
  assign n6202 = n156 & n6201 ;
  assign n6203 = n20601 & n6202 ;
  assign n20710 = ~n6202 ;
  assign n6204 = n5872 & n20710 ;
  assign n6205 = n6203 | n6204 ;
  assign n20711 = ~n6205 ;
  assign n6206 = n6200 & n20711 ;
  assign n6207 = n6199 | n6206 ;
  assign n6208 = x72 & n6207 ;
  assign n6209 = x72 | n6207 ;
  assign n20712 = ~n5875 ;
  assign n6210 = n20712 & n5876 ;
  assign n6211 = n156 & n6210 ;
  assign n6212 = n20604 & n6211 ;
  assign n20713 = ~n6211 ;
  assign n6213 = n5881 & n20713 ;
  assign n6214 = n6212 | n6213 ;
  assign n20714 = ~n6214 ;
  assign n6215 = n6209 & n20714 ;
  assign n6216 = n6208 | n6215 ;
  assign n6217 = x73 & n6216 ;
  assign n6218 = x73 | n6216 ;
  assign n20715 = ~n5884 ;
  assign n6219 = n20715 & n5885 ;
  assign n6220 = n156 & n6219 ;
  assign n6221 = n20607 & n6220 ;
  assign n20716 = ~n6220 ;
  assign n6222 = n5890 & n20716 ;
  assign n6223 = n6221 | n6222 ;
  assign n20717 = ~n6223 ;
  assign n6224 = n6218 & n20717 ;
  assign n6225 = n6217 | n6224 ;
  assign n6226 = x74 & n6225 ;
  assign n6227 = x74 | n6225 ;
  assign n20718 = ~n5893 ;
  assign n6228 = n20718 & n5894 ;
  assign n6229 = n156 & n6228 ;
  assign n6230 = n20610 & n6229 ;
  assign n20719 = ~n6229 ;
  assign n6231 = n5899 & n20719 ;
  assign n6232 = n6230 | n6231 ;
  assign n20720 = ~n6232 ;
  assign n6233 = n6227 & n20720 ;
  assign n6234 = n6226 | n6233 ;
  assign n6235 = x75 & n6234 ;
  assign n6236 = x75 | n6234 ;
  assign n20721 = ~n5902 ;
  assign n6237 = n20721 & n5903 ;
  assign n6238 = n156 & n6237 ;
  assign n6239 = n20613 & n6238 ;
  assign n20722 = ~n6238 ;
  assign n6240 = n5908 & n20722 ;
  assign n6241 = n6239 | n6240 ;
  assign n20723 = ~n6241 ;
  assign n6242 = n6236 & n20723 ;
  assign n6243 = n6235 | n6242 ;
  assign n6244 = x76 & n6243 ;
  assign n6245 = x76 | n6243 ;
  assign n20724 = ~n5911 ;
  assign n6246 = n20724 & n5912 ;
  assign n6247 = n156 & n6246 ;
  assign n6248 = n5917 & n6247 ;
  assign n6249 = n5917 | n6247 ;
  assign n20725 = ~n6248 ;
  assign n6250 = n20725 & n6249 ;
  assign n20726 = ~n6250 ;
  assign n6251 = n6245 & n20726 ;
  assign n6252 = n6244 | n6251 ;
  assign n6253 = x77 & n6252 ;
  assign n6254 = x77 | n6252 ;
  assign n20727 = ~n5920 ;
  assign n6255 = n20727 & n5921 ;
  assign n6256 = n156 & n6255 ;
  assign n6257 = n20619 & n6256 ;
  assign n20728 = ~n6256 ;
  assign n6258 = n5926 & n20728 ;
  assign n6259 = n6257 | n6258 ;
  assign n20729 = ~n6259 ;
  assign n6260 = n6254 & n20729 ;
  assign n6261 = n6253 | n6260 ;
  assign n6262 = x78 & n6261 ;
  assign n6263 = x78 | n6261 ;
  assign n20730 = ~n5929 ;
  assign n6264 = n20730 & n5930 ;
  assign n6265 = n156 & n6264 ;
  assign n6266 = n5935 & n6265 ;
  assign n6267 = n5935 | n6265 ;
  assign n20731 = ~n6266 ;
  assign n6268 = n20731 & n6267 ;
  assign n20732 = ~n6268 ;
  assign n6269 = n6263 & n20732 ;
  assign n6270 = n6262 | n6269 ;
  assign n6271 = x79 & n6270 ;
  assign n6272 = x79 | n6270 ;
  assign n20733 = ~n5938 ;
  assign n6273 = n20733 & n5939 ;
  assign n6274 = n156 & n6273 ;
  assign n6275 = n5944 & n6274 ;
  assign n6276 = n5944 | n6274 ;
  assign n20734 = ~n6275 ;
  assign n6277 = n20734 & n6276 ;
  assign n20735 = ~n6277 ;
  assign n6278 = n6272 & n20735 ;
  assign n6279 = n6271 | n6278 ;
  assign n6280 = x80 & n6279 ;
  assign n6281 = x80 | n6279 ;
  assign n20736 = ~n5947 ;
  assign n6282 = n20736 & n5948 ;
  assign n6283 = n156 & n6282 ;
  assign n6284 = n20628 & n6283 ;
  assign n20737 = ~n6283 ;
  assign n6285 = n5953 & n20737 ;
  assign n6286 = n6284 | n6285 ;
  assign n20738 = ~n6286 ;
  assign n6287 = n6281 & n20738 ;
  assign n6288 = n6280 | n6287 ;
  assign n6289 = x81 & n6288 ;
  assign n6290 = x81 | n6288 ;
  assign n20739 = ~n5956 ;
  assign n6291 = n20739 & n5957 ;
  assign n6292 = n156 & n6291 ;
  assign n6293 = n20631 & n6292 ;
  assign n20740 = ~n6292 ;
  assign n6294 = n5962 & n20740 ;
  assign n6295 = n6293 | n6294 ;
  assign n20741 = ~n6295 ;
  assign n6296 = n6290 & n20741 ;
  assign n6297 = n6289 | n6296 ;
  assign n6298 = x82 & n6297 ;
  assign n6299 = x82 | n6297 ;
  assign n20742 = ~n5965 ;
  assign n6300 = n20742 & n5966 ;
  assign n6301 = n156 & n6300 ;
  assign n6302 = n20634 & n6301 ;
  assign n20743 = ~n6301 ;
  assign n6303 = n5971 & n20743 ;
  assign n6304 = n6302 | n6303 ;
  assign n20744 = ~n6304 ;
  assign n6305 = n6299 & n20744 ;
  assign n6306 = n6298 | n6305 ;
  assign n6307 = x83 & n6306 ;
  assign n6308 = x83 | n6306 ;
  assign n20745 = ~n5974 ;
  assign n6309 = n20745 & n5975 ;
  assign n6310 = n156 & n6309 ;
  assign n6311 = n5980 & n6310 ;
  assign n6312 = n5980 | n6310 ;
  assign n20746 = ~n6311 ;
  assign n6313 = n20746 & n6312 ;
  assign n20747 = ~n6313 ;
  assign n6314 = n6308 & n20747 ;
  assign n6315 = n6307 | n6314 ;
  assign n6316 = x84 & n6315 ;
  assign n6317 = x84 | n6315 ;
  assign n20748 = ~n5983 ;
  assign n6318 = n20748 & n5984 ;
  assign n6319 = n156 & n6318 ;
  assign n6320 = n5989 & n6319 ;
  assign n6321 = n5989 | n6319 ;
  assign n20749 = ~n6320 ;
  assign n6322 = n20749 & n6321 ;
  assign n20750 = ~n6322 ;
  assign n6323 = n6317 & n20750 ;
  assign n6324 = n6316 | n6323 ;
  assign n6325 = x85 & n6324 ;
  assign n6326 = x85 | n6324 ;
  assign n20751 = ~n5992 ;
  assign n6327 = n20751 & n5993 ;
  assign n6328 = n156 & n6327 ;
  assign n6329 = n5998 & n6328 ;
  assign n6330 = n5998 | n6328 ;
  assign n20752 = ~n6329 ;
  assign n6331 = n20752 & n6330 ;
  assign n20753 = ~n6331 ;
  assign n6332 = n6326 & n20753 ;
  assign n6333 = n6325 | n6332 ;
  assign n6334 = x86 & n6333 ;
  assign n6335 = x86 | n6333 ;
  assign n20754 = ~n6001 ;
  assign n6336 = n20754 & n6002 ;
  assign n6337 = n156 & n6336 ;
  assign n6338 = n20646 & n6337 ;
  assign n20755 = ~n6337 ;
  assign n6339 = n6007 & n20755 ;
  assign n6340 = n6338 | n6339 ;
  assign n20756 = ~n6340 ;
  assign n6341 = n6335 & n20756 ;
  assign n6342 = n6334 | n6341 ;
  assign n6343 = x87 & n6342 ;
  assign n6344 = x87 | n6342 ;
  assign n20757 = ~n6010 ;
  assign n6345 = n20757 & n6011 ;
  assign n6346 = n156 & n6345 ;
  assign n6347 = n20649 & n6346 ;
  assign n20758 = ~n6346 ;
  assign n6348 = n6016 & n20758 ;
  assign n6349 = n6347 | n6348 ;
  assign n20759 = ~n6349 ;
  assign n6350 = n6344 & n20759 ;
  assign n6351 = n6343 | n6350 ;
  assign n6352 = x88 & n6351 ;
  assign n6353 = x88 | n6351 ;
  assign n20760 = ~n6019 ;
  assign n6354 = n20760 & n6020 ;
  assign n6355 = n156 & n6354 ;
  assign n6356 = n20652 & n6355 ;
  assign n20761 = ~n6355 ;
  assign n6357 = n6025 & n20761 ;
  assign n6358 = n6356 | n6357 ;
  assign n20762 = ~n6358 ;
  assign n6359 = n6353 & n20762 ;
  assign n6360 = n6352 | n6359 ;
  assign n6361 = x89 & n6360 ;
  assign n6362 = x89 | n6360 ;
  assign n20763 = ~n6028 ;
  assign n6363 = n20763 & n6029 ;
  assign n6364 = n156 & n6363 ;
  assign n6365 = n20655 & n6364 ;
  assign n20764 = ~n6364 ;
  assign n6366 = n6034 & n20764 ;
  assign n6367 = n6365 | n6366 ;
  assign n20765 = ~n6367 ;
  assign n6368 = n6362 & n20765 ;
  assign n6369 = n6361 | n6368 ;
  assign n6370 = x90 & n6369 ;
  assign n6371 = x90 | n6369 ;
  assign n20766 = ~n6037 ;
  assign n6372 = n20766 & n6038 ;
  assign n6373 = n156 & n6372 ;
  assign n6374 = n20658 & n6373 ;
  assign n20767 = ~n6373 ;
  assign n6375 = n6043 & n20767 ;
  assign n6376 = n6374 | n6375 ;
  assign n20768 = ~n6376 ;
  assign n6377 = n6371 & n20768 ;
  assign n6378 = n6370 | n6377 ;
  assign n6379 = x91 & n6378 ;
  assign n6380 = x91 | n6378 ;
  assign n20769 = ~n6046 ;
  assign n6381 = n20769 & n6047 ;
  assign n6382 = n156 & n6381 ;
  assign n6383 = n20661 & n6382 ;
  assign n20770 = ~n6382 ;
  assign n6384 = n6052 & n20770 ;
  assign n6385 = n6383 | n6384 ;
  assign n20771 = ~n6385 ;
  assign n6386 = n6380 & n20771 ;
  assign n6387 = n6379 | n6386 ;
  assign n6388 = x92 & n6387 ;
  assign n6389 = x92 | n6387 ;
  assign n20772 = ~n6055 ;
  assign n6390 = n20772 & n6056 ;
  assign n6391 = n156 & n6390 ;
  assign n6392 = n20664 & n6391 ;
  assign n20773 = ~n6391 ;
  assign n6393 = n6061 & n20773 ;
  assign n6394 = n6392 | n6393 ;
  assign n20774 = ~n6394 ;
  assign n6395 = n6389 & n20774 ;
  assign n6396 = n6388 | n6395 ;
  assign n6397 = x93 & n6396 ;
  assign n6398 = x93 | n6396 ;
  assign n20775 = ~n6064 ;
  assign n6399 = n20775 & n6065 ;
  assign n6400 = n156 & n6399 ;
  assign n6401 = n20667 & n6400 ;
  assign n20776 = ~n6400 ;
  assign n6402 = n6070 & n20776 ;
  assign n6403 = n6401 | n6402 ;
  assign n20777 = ~n6403 ;
  assign n6404 = n6398 & n20777 ;
  assign n6405 = n6397 | n6404 ;
  assign n6406 = x94 & n6405 ;
  assign n6407 = x94 | n6405 ;
  assign n20778 = ~n6073 ;
  assign n6408 = n20778 & n6074 ;
  assign n6409 = n156 & n6408 ;
  assign n6410 = n20670 & n6409 ;
  assign n20779 = ~n6409 ;
  assign n6411 = n6079 & n20779 ;
  assign n6412 = n6410 | n6411 ;
  assign n20780 = ~n6412 ;
  assign n6413 = n6407 & n20780 ;
  assign n6414 = n6406 | n6413 ;
  assign n6415 = x95 & n6414 ;
  assign n6416 = x95 | n6414 ;
  assign n20781 = ~n6082 ;
  assign n6417 = n20781 & n6083 ;
  assign n6418 = n156 & n6417 ;
  assign n6419 = n20673 & n6418 ;
  assign n20782 = ~n6418 ;
  assign n6420 = n6088 & n20782 ;
  assign n6421 = n6419 | n6420 ;
  assign n20783 = ~n6421 ;
  assign n6422 = n6416 & n20783 ;
  assign n6423 = n6415 | n6422 ;
  assign n6424 = x96 & n6423 ;
  assign n6425 = x96 | n6423 ;
  assign n20784 = ~n6091 ;
  assign n6426 = n20784 & n6092 ;
  assign n6427 = n156 & n6426 ;
  assign n6428 = n20676 & n6427 ;
  assign n20785 = ~n6427 ;
  assign n6429 = n6097 & n20785 ;
  assign n6430 = n6428 | n6429 ;
  assign n20786 = ~n6430 ;
  assign n6431 = n6425 & n20786 ;
  assign n6432 = n6424 | n6431 ;
  assign n6433 = x97 & n6432 ;
  assign n6434 = x97 | n6432 ;
  assign n20787 = ~n6100 ;
  assign n6435 = n20787 & n6101 ;
  assign n6436 = n156 & n6435 ;
  assign n6437 = n20679 & n6436 ;
  assign n20788 = ~n6436 ;
  assign n6438 = n6106 & n20788 ;
  assign n6439 = n6437 | n6438 ;
  assign n20789 = ~n6439 ;
  assign n6440 = n6434 & n20789 ;
  assign n6441 = n6433 | n6440 ;
  assign n6442 = x98 & n6441 ;
  assign n6443 = x98 | n6441 ;
  assign n20790 = ~n6109 ;
  assign n6444 = n20790 & n6110 ;
  assign n6445 = n156 & n6444 ;
  assign n6446 = n20682 & n6445 ;
  assign n20791 = ~n6445 ;
  assign n6447 = n6115 & n20791 ;
  assign n6448 = n6446 | n6447 ;
  assign n20792 = ~n6448 ;
  assign n6449 = n6443 & n20792 ;
  assign n6450 = n6442 | n6449 ;
  assign n6451 = x99 & n6450 ;
  assign n6452 = x99 | n6450 ;
  assign n20793 = ~n6118 ;
  assign n6453 = n20793 & n6119 ;
  assign n6454 = n156 & n6453 ;
  assign n6455 = n20685 & n6454 ;
  assign n20794 = ~n6454 ;
  assign n6456 = n6124 & n20794 ;
  assign n6457 = n6455 | n6456 ;
  assign n20795 = ~n6457 ;
  assign n6458 = n6452 & n20795 ;
  assign n6459 = n6451 | n6458 ;
  assign n6460 = x100 & n6459 ;
  assign n6461 = x100 | n6459 ;
  assign n20796 = ~n6143 ;
  assign n6462 = n20796 & n6461 ;
  assign n6463 = n6460 | n6462 ;
  assign n6464 = x101 | n6463 ;
  assign n20797 = ~n6145 ;
  assign n6465 = n20797 & n6464 ;
  assign n6466 = x101 & n6463 ;
  assign n6467 = n18388 | n6466 ;
  assign n6469 = n6465 | n6467 ;
  assign n20798 = ~n6460 ;
  assign n6470 = n20798 & n6461 ;
  assign n155 = ~n6469 ;
  assign n6471 = n155 & n6470 ;
  assign n6472 = n6143 & n6471 ;
  assign n6473 = n6143 | n6471 ;
  assign n20800 = ~n6472 ;
  assign n6474 = n20800 & n6473 ;
  assign n6468 = n6144 & n6467 ;
  assign n6475 = n21884 | n6468 ;
  assign n20801 = ~n18388 ;
  assign n6477 = n20801 & n6475 ;
  assign n20802 = ~x25 ;
  assign n6478 = n20802 & x64 ;
  assign n6480 = x65 | n6478 ;
  assign n6479 = x65 & n6478 ;
  assign n6481 = x64 & n155 ;
  assign n6482 = x26 & n6481 ;
  assign n6483 = x26 | n6481 ;
  assign n20803 = ~n6482 ;
  assign n6484 = n20803 & n6483 ;
  assign n20804 = ~n6479 ;
  assign n6485 = n20804 & n6484 ;
  assign n20805 = ~n6485 ;
  assign n6486 = n6480 & n20805 ;
  assign n6487 = x66 | n6486 ;
  assign n6488 = x66 & n6486 ;
  assign n6489 = n6147 & n155 ;
  assign n6490 = n20693 & n6489 ;
  assign n6491 = n6150 | n6490 ;
  assign n6492 = n6152 & n6489 ;
  assign n20806 = ~n6492 ;
  assign n6493 = n6491 & n20806 ;
  assign n20807 = ~n6488 ;
  assign n6494 = n20807 & n6493 ;
  assign n20808 = ~n6494 ;
  assign n6495 = n6487 & n20808 ;
  assign n6496 = x67 | n6495 ;
  assign n6497 = x67 & n6495 ;
  assign n20809 = ~n6154 ;
  assign n6498 = n20809 & n6160 ;
  assign n6499 = n155 & n6498 ;
  assign n6500 = n6159 & n6499 ;
  assign n6501 = n6159 | n6499 ;
  assign n20810 = ~n6500 ;
  assign n6502 = n20810 & n6501 ;
  assign n20811 = ~n6497 ;
  assign n6503 = n20811 & n6502 ;
  assign n20812 = ~n6503 ;
  assign n6504 = n6496 & n20812 ;
  assign n6505 = x68 | n6504 ;
  assign n6506 = x68 & n6504 ;
  assign n20813 = ~n6163 ;
  assign n6507 = n20813 & n6164 ;
  assign n6508 = n155 & n6507 ;
  assign n6509 = n6169 & n6508 ;
  assign n6510 = n6169 | n6508 ;
  assign n20814 = ~n6509 ;
  assign n6511 = n20814 & n6510 ;
  assign n20815 = ~n6506 ;
  assign n6512 = n20815 & n6511 ;
  assign n20816 = ~n6512 ;
  assign n6513 = n6505 & n20816 ;
  assign n6514 = x69 | n6513 ;
  assign n6515 = x69 & n6513 ;
  assign n20817 = ~n6172 ;
  assign n6516 = n20817 & n6173 ;
  assign n6517 = n155 & n6516 ;
  assign n6518 = n6178 & n6517 ;
  assign n6519 = n6178 | n6517 ;
  assign n20818 = ~n6518 ;
  assign n6520 = n20818 & n6519 ;
  assign n20819 = ~n6515 ;
  assign n6521 = n20819 & n6520 ;
  assign n20820 = ~n6521 ;
  assign n6522 = n6514 & n20820 ;
  assign n6523 = x70 | n6522 ;
  assign n6524 = x70 & n6522 ;
  assign n20821 = ~n6181 ;
  assign n6525 = n20821 & n6182 ;
  assign n6526 = n155 & n6525 ;
  assign n6527 = n6187 & n6526 ;
  assign n6528 = n6187 | n6526 ;
  assign n20822 = ~n6527 ;
  assign n6529 = n20822 & n6528 ;
  assign n20823 = ~n6524 ;
  assign n6530 = n20823 & n6529 ;
  assign n20824 = ~n6530 ;
  assign n6531 = n6523 & n20824 ;
  assign n6532 = x71 | n6531 ;
  assign n6533 = x71 & n6531 ;
  assign n20825 = ~n6190 ;
  assign n6534 = n20825 & n6191 ;
  assign n6535 = n155 & n6534 ;
  assign n6536 = n6196 & n6535 ;
  assign n6537 = n6196 | n6535 ;
  assign n20826 = ~n6536 ;
  assign n6538 = n20826 & n6537 ;
  assign n20827 = ~n6533 ;
  assign n6539 = n20827 & n6538 ;
  assign n20828 = ~n6539 ;
  assign n6540 = n6532 & n20828 ;
  assign n6541 = x72 | n6540 ;
  assign n6542 = x72 & n6540 ;
  assign n20829 = ~n6199 ;
  assign n6543 = n20829 & n6200 ;
  assign n6544 = n155 & n6543 ;
  assign n6545 = n6205 & n6544 ;
  assign n6546 = n6205 | n6544 ;
  assign n20830 = ~n6545 ;
  assign n6547 = n20830 & n6546 ;
  assign n20831 = ~n6542 ;
  assign n6548 = n20831 & n6547 ;
  assign n20832 = ~n6548 ;
  assign n6549 = n6541 & n20832 ;
  assign n6550 = x73 | n6549 ;
  assign n6551 = x73 & n6549 ;
  assign n20833 = ~n6208 ;
  assign n6552 = n20833 & n6209 ;
  assign n6553 = n155 & n6552 ;
  assign n6554 = n20714 & n6553 ;
  assign n20834 = ~n6553 ;
  assign n6555 = n6214 & n20834 ;
  assign n6556 = n6554 | n6555 ;
  assign n20835 = ~n6551 ;
  assign n6557 = n20835 & n6556 ;
  assign n20836 = ~n6557 ;
  assign n6558 = n6550 & n20836 ;
  assign n6559 = x74 | n6558 ;
  assign n6560 = x74 & n6558 ;
  assign n20837 = ~n6217 ;
  assign n6561 = n20837 & n6218 ;
  assign n6562 = n155 & n6561 ;
  assign n6563 = n20717 & n6562 ;
  assign n20838 = ~n6562 ;
  assign n6564 = n6223 & n20838 ;
  assign n6565 = n6563 | n6564 ;
  assign n20839 = ~n6560 ;
  assign n6566 = n20839 & n6565 ;
  assign n20840 = ~n6566 ;
  assign n6567 = n6559 & n20840 ;
  assign n6568 = x75 | n6567 ;
  assign n6569 = x75 & n6567 ;
  assign n20841 = ~n6226 ;
  assign n6570 = n20841 & n6227 ;
  assign n6571 = n155 & n6570 ;
  assign n6572 = n6232 & n6571 ;
  assign n6573 = n6232 | n6571 ;
  assign n20842 = ~n6572 ;
  assign n6574 = n20842 & n6573 ;
  assign n20843 = ~n6569 ;
  assign n6575 = n20843 & n6574 ;
  assign n20844 = ~n6575 ;
  assign n6576 = n6568 & n20844 ;
  assign n6577 = x76 | n6576 ;
  assign n6578 = x76 & n6576 ;
  assign n20845 = ~n6235 ;
  assign n6579 = n20845 & n6236 ;
  assign n6580 = n155 & n6579 ;
  assign n6581 = n6241 & n6580 ;
  assign n6582 = n6241 | n6580 ;
  assign n20846 = ~n6581 ;
  assign n6583 = n20846 & n6582 ;
  assign n20847 = ~n6578 ;
  assign n6584 = n20847 & n6583 ;
  assign n20848 = ~n6584 ;
  assign n6585 = n6577 & n20848 ;
  assign n6586 = x77 | n6585 ;
  assign n6587 = x77 & n6585 ;
  assign n20849 = ~n6244 ;
  assign n6588 = n20849 & n6245 ;
  assign n6589 = n155 & n6588 ;
  assign n6590 = n6250 & n6589 ;
  assign n6591 = n6250 | n6589 ;
  assign n20850 = ~n6590 ;
  assign n6592 = n20850 & n6591 ;
  assign n20851 = ~n6587 ;
  assign n6593 = n20851 & n6592 ;
  assign n20852 = ~n6593 ;
  assign n6594 = n6586 & n20852 ;
  assign n6595 = x78 | n6594 ;
  assign n6596 = x78 & n6594 ;
  assign n20853 = ~n6253 ;
  assign n6597 = n20853 & n6254 ;
  assign n6598 = n155 & n6597 ;
  assign n6599 = n6259 & n6598 ;
  assign n6600 = n6259 | n6598 ;
  assign n20854 = ~n6599 ;
  assign n6601 = n20854 & n6600 ;
  assign n20855 = ~n6596 ;
  assign n6602 = n20855 & n6601 ;
  assign n20856 = ~n6602 ;
  assign n6603 = n6595 & n20856 ;
  assign n6604 = x79 | n6603 ;
  assign n6605 = x79 & n6603 ;
  assign n20857 = ~n6262 ;
  assign n6606 = n20857 & n6263 ;
  assign n6607 = n155 & n6606 ;
  assign n6608 = n20732 & n6607 ;
  assign n20858 = ~n6607 ;
  assign n6609 = n6268 & n20858 ;
  assign n6610 = n6608 | n6609 ;
  assign n20859 = ~n6605 ;
  assign n6611 = n20859 & n6610 ;
  assign n20860 = ~n6611 ;
  assign n6612 = n6604 & n20860 ;
  assign n6613 = x80 | n6612 ;
  assign n6614 = x80 & n6612 ;
  assign n20861 = ~n6271 ;
  assign n6615 = n20861 & n6272 ;
  assign n6616 = n155 & n6615 ;
  assign n6617 = n6277 & n6616 ;
  assign n6618 = n6277 | n6616 ;
  assign n20862 = ~n6617 ;
  assign n6619 = n20862 & n6618 ;
  assign n20863 = ~n6614 ;
  assign n6620 = n20863 & n6619 ;
  assign n20864 = ~n6620 ;
  assign n6621 = n6613 & n20864 ;
  assign n6622 = x81 | n6621 ;
  assign n6623 = x81 & n6621 ;
  assign n20865 = ~n6280 ;
  assign n6624 = n20865 & n6281 ;
  assign n6625 = n155 & n6624 ;
  assign n6626 = n20738 & n6625 ;
  assign n20866 = ~n6625 ;
  assign n6627 = n6286 & n20866 ;
  assign n6628 = n6626 | n6627 ;
  assign n20867 = ~n6623 ;
  assign n6629 = n20867 & n6628 ;
  assign n20868 = ~n6629 ;
  assign n6630 = n6622 & n20868 ;
  assign n6631 = x82 | n6630 ;
  assign n6632 = x82 & n6630 ;
  assign n20869 = ~n6289 ;
  assign n6633 = n20869 & n6290 ;
  assign n6634 = n155 & n6633 ;
  assign n6635 = n6295 & n6634 ;
  assign n6636 = n6295 | n6634 ;
  assign n20870 = ~n6635 ;
  assign n6637 = n20870 & n6636 ;
  assign n20871 = ~n6632 ;
  assign n6638 = n20871 & n6637 ;
  assign n20872 = ~n6638 ;
  assign n6639 = n6631 & n20872 ;
  assign n6640 = x83 | n6639 ;
  assign n6641 = x83 & n6639 ;
  assign n20873 = ~n6298 ;
  assign n6642 = n20873 & n6299 ;
  assign n6643 = n155 & n6642 ;
  assign n6644 = n6304 & n6643 ;
  assign n6645 = n6304 | n6643 ;
  assign n20874 = ~n6644 ;
  assign n6646 = n20874 & n6645 ;
  assign n20875 = ~n6641 ;
  assign n6647 = n20875 & n6646 ;
  assign n20876 = ~n6647 ;
  assign n6648 = n6640 & n20876 ;
  assign n6649 = x84 | n6648 ;
  assign n6650 = x84 & n6648 ;
  assign n20877 = ~n6307 ;
  assign n6651 = n20877 & n6308 ;
  assign n6652 = n155 & n6651 ;
  assign n6653 = n6313 & n6652 ;
  assign n6654 = n6313 | n6652 ;
  assign n20878 = ~n6653 ;
  assign n6655 = n20878 & n6654 ;
  assign n20879 = ~n6650 ;
  assign n6656 = n20879 & n6655 ;
  assign n20880 = ~n6656 ;
  assign n6657 = n6649 & n20880 ;
  assign n6658 = x85 | n6657 ;
  assign n6659 = x85 & n6657 ;
  assign n20881 = ~n6316 ;
  assign n6660 = n20881 & n6317 ;
  assign n6661 = n155 & n6660 ;
  assign n6662 = n6322 & n6661 ;
  assign n6663 = n6322 | n6661 ;
  assign n20882 = ~n6662 ;
  assign n6664 = n20882 & n6663 ;
  assign n20883 = ~n6659 ;
  assign n6665 = n20883 & n6664 ;
  assign n20884 = ~n6665 ;
  assign n6666 = n6658 & n20884 ;
  assign n6667 = x86 | n6666 ;
  assign n6668 = x86 & n6666 ;
  assign n20885 = ~n6325 ;
  assign n6669 = n20885 & n6326 ;
  assign n6670 = n155 & n6669 ;
  assign n6671 = n6331 & n6670 ;
  assign n6672 = n6331 | n6670 ;
  assign n20886 = ~n6671 ;
  assign n6673 = n20886 & n6672 ;
  assign n20887 = ~n6668 ;
  assign n6674 = n20887 & n6673 ;
  assign n20888 = ~n6674 ;
  assign n6675 = n6667 & n20888 ;
  assign n6676 = x87 | n6675 ;
  assign n6677 = x87 & n6675 ;
  assign n20889 = ~n6334 ;
  assign n6678 = n20889 & n6335 ;
  assign n6679 = n155 & n6678 ;
  assign n6680 = n20756 & n6679 ;
  assign n20890 = ~n6679 ;
  assign n6681 = n6340 & n20890 ;
  assign n6682 = n6680 | n6681 ;
  assign n20891 = ~n6677 ;
  assign n6683 = n20891 & n6682 ;
  assign n20892 = ~n6683 ;
  assign n6684 = n6676 & n20892 ;
  assign n6685 = x88 | n6684 ;
  assign n6686 = x88 & n6684 ;
  assign n20893 = ~n6343 ;
  assign n6687 = n20893 & n6344 ;
  assign n6688 = n155 & n6687 ;
  assign n6689 = n20759 & n6688 ;
  assign n20894 = ~n6688 ;
  assign n6690 = n6349 & n20894 ;
  assign n6691 = n6689 | n6690 ;
  assign n20895 = ~n6686 ;
  assign n6692 = n20895 & n6691 ;
  assign n20896 = ~n6692 ;
  assign n6693 = n6685 & n20896 ;
  assign n6694 = x89 | n6693 ;
  assign n6695 = x89 & n6693 ;
  assign n20897 = ~n6352 ;
  assign n6696 = n20897 & n6353 ;
  assign n6697 = n155 & n6696 ;
  assign n6698 = n20762 & n6697 ;
  assign n20898 = ~n6697 ;
  assign n6699 = n6358 & n20898 ;
  assign n6700 = n6698 | n6699 ;
  assign n20899 = ~n6695 ;
  assign n6701 = n20899 & n6700 ;
  assign n20900 = ~n6701 ;
  assign n6702 = n6694 & n20900 ;
  assign n6703 = x90 | n6702 ;
  assign n6704 = x90 & n6702 ;
  assign n20901 = ~n6361 ;
  assign n6705 = n20901 & n6362 ;
  assign n6706 = n155 & n6705 ;
  assign n6707 = n20765 & n6706 ;
  assign n20902 = ~n6706 ;
  assign n6708 = n6367 & n20902 ;
  assign n6709 = n6707 | n6708 ;
  assign n20903 = ~n6704 ;
  assign n6710 = n20903 & n6709 ;
  assign n20904 = ~n6710 ;
  assign n6711 = n6703 & n20904 ;
  assign n6712 = x91 | n6711 ;
  assign n6713 = x91 & n6711 ;
  assign n20905 = ~n6370 ;
  assign n6714 = n20905 & n6371 ;
  assign n6715 = n155 & n6714 ;
  assign n6716 = n20768 & n6715 ;
  assign n20906 = ~n6715 ;
  assign n6717 = n6376 & n20906 ;
  assign n6718 = n6716 | n6717 ;
  assign n20907 = ~n6713 ;
  assign n6719 = n20907 & n6718 ;
  assign n20908 = ~n6719 ;
  assign n6720 = n6712 & n20908 ;
  assign n6721 = x92 | n6720 ;
  assign n6722 = x92 & n6720 ;
  assign n20909 = ~n6379 ;
  assign n6723 = n20909 & n6380 ;
  assign n6724 = n155 & n6723 ;
  assign n6725 = n20771 & n6724 ;
  assign n20910 = ~n6724 ;
  assign n6726 = n6385 & n20910 ;
  assign n6727 = n6725 | n6726 ;
  assign n20911 = ~n6722 ;
  assign n6728 = n20911 & n6727 ;
  assign n20912 = ~n6728 ;
  assign n6729 = n6721 & n20912 ;
  assign n6730 = x93 | n6729 ;
  assign n6731 = x93 & n6729 ;
  assign n20913 = ~n6388 ;
  assign n6732 = n20913 & n6389 ;
  assign n6733 = n155 & n6732 ;
  assign n6734 = n20774 & n6733 ;
  assign n20914 = ~n6733 ;
  assign n6735 = n6394 & n20914 ;
  assign n6736 = n6734 | n6735 ;
  assign n20915 = ~n6731 ;
  assign n6737 = n20915 & n6736 ;
  assign n20916 = ~n6737 ;
  assign n6738 = n6730 & n20916 ;
  assign n6739 = x94 | n6738 ;
  assign n6740 = x94 & n6738 ;
  assign n20917 = ~n6397 ;
  assign n6741 = n20917 & n6398 ;
  assign n6742 = n155 & n6741 ;
  assign n6743 = n20777 & n6742 ;
  assign n20918 = ~n6742 ;
  assign n6744 = n6403 & n20918 ;
  assign n6745 = n6743 | n6744 ;
  assign n20919 = ~n6740 ;
  assign n6746 = n20919 & n6745 ;
  assign n20920 = ~n6746 ;
  assign n6747 = n6739 & n20920 ;
  assign n6748 = x95 | n6747 ;
  assign n6749 = x95 & n6747 ;
  assign n20921 = ~n6406 ;
  assign n6750 = n20921 & n6407 ;
  assign n6751 = n155 & n6750 ;
  assign n6752 = n20780 & n6751 ;
  assign n20922 = ~n6751 ;
  assign n6753 = n6412 & n20922 ;
  assign n6754 = n6752 | n6753 ;
  assign n20923 = ~n6749 ;
  assign n6755 = n20923 & n6754 ;
  assign n20924 = ~n6755 ;
  assign n6756 = n6748 & n20924 ;
  assign n6757 = x96 | n6756 ;
  assign n6758 = x96 & n6756 ;
  assign n20925 = ~n6415 ;
  assign n6759 = n20925 & n6416 ;
  assign n6760 = n155 & n6759 ;
  assign n6761 = n20783 & n6760 ;
  assign n20926 = ~n6760 ;
  assign n6762 = n6421 & n20926 ;
  assign n6763 = n6761 | n6762 ;
  assign n20927 = ~n6758 ;
  assign n6764 = n20927 & n6763 ;
  assign n20928 = ~n6764 ;
  assign n6765 = n6757 & n20928 ;
  assign n6766 = x97 | n6765 ;
  assign n6767 = x97 & n6765 ;
  assign n20929 = ~n6424 ;
  assign n6768 = n20929 & n6425 ;
  assign n6769 = n155 & n6768 ;
  assign n6770 = n20786 & n6769 ;
  assign n20930 = ~n6769 ;
  assign n6771 = n6430 & n20930 ;
  assign n6772 = n6770 | n6771 ;
  assign n20931 = ~n6767 ;
  assign n6773 = n20931 & n6772 ;
  assign n20932 = ~n6773 ;
  assign n6774 = n6766 & n20932 ;
  assign n6775 = x98 | n6774 ;
  assign n6776 = x98 & n6774 ;
  assign n20933 = ~n6433 ;
  assign n6777 = n20933 & n6434 ;
  assign n6778 = n155 & n6777 ;
  assign n6779 = n20789 & n6778 ;
  assign n20934 = ~n6778 ;
  assign n6780 = n6439 & n20934 ;
  assign n6781 = n6779 | n6780 ;
  assign n20935 = ~n6776 ;
  assign n6782 = n20935 & n6781 ;
  assign n20936 = ~n6782 ;
  assign n6783 = n6775 & n20936 ;
  assign n6784 = x99 | n6783 ;
  assign n6785 = x99 & n6783 ;
  assign n20937 = ~n6442 ;
  assign n6786 = n20937 & n6443 ;
  assign n6787 = n155 & n6786 ;
  assign n6788 = n20792 & n6787 ;
  assign n20938 = ~n6787 ;
  assign n6789 = n6448 & n20938 ;
  assign n6790 = n6788 | n6789 ;
  assign n20939 = ~n6785 ;
  assign n6791 = n20939 & n6790 ;
  assign n20940 = ~n6791 ;
  assign n6792 = n6784 & n20940 ;
  assign n6793 = x100 | n6792 ;
  assign n6794 = x100 & n6792 ;
  assign n20941 = ~n6451 ;
  assign n6795 = n20941 & n6452 ;
  assign n6796 = n155 & n6795 ;
  assign n6797 = n20795 & n6796 ;
  assign n20942 = ~n6796 ;
  assign n6798 = n6457 & n20942 ;
  assign n6799 = n6797 | n6798 ;
  assign n20943 = ~n6794 ;
  assign n6800 = n20943 & n6799 ;
  assign n20944 = ~n6800 ;
  assign n6801 = n6793 & n20944 ;
  assign n6803 = x101 | n6801 ;
  assign n20945 = ~n6474 ;
  assign n6804 = n20945 & n6803 ;
  assign n6802 = x101 & n6801 ;
  assign n20946 = ~x102 ;
  assign n6476 = n20946 & n6475 ;
  assign n6805 = n18383 | n6476 ;
  assign n20947 = ~n6475 ;
  assign n6806 = x102 & n20947 ;
  assign n6807 = n6805 | n6806 ;
  assign n6808 = n6802 | n6807 ;
  assign n6809 = n6804 | n6808 ;
  assign n20948 = ~n6477 ;
  assign n6810 = n20948 & n6809 ;
  assign n20949 = ~n6802 ;
  assign n6811 = n20949 & n6803 ;
  assign n154 = ~n6810 ;
  assign n6812 = n154 & n6811 ;
  assign n6813 = n6474 & n6812 ;
  assign n6814 = n6474 | n6812 ;
  assign n20951 = ~n6813 ;
  assign n6815 = n20951 & n6814 ;
  assign n6816 = n6145 & n6809 ;
  assign n6817 = n18388 & n6816 ;
  assign n6818 = n21884 | n6817 ;
  assign n20952 = ~x24 ;
  assign n6819 = n20952 & x64 ;
  assign n6820 = x65 | n6819 ;
  assign n6821 = x64 & n154 ;
  assign n20953 = ~n6821 ;
  assign n6822 = x25 & n20953 ;
  assign n6823 = n6478 & n154 ;
  assign n6824 = n6822 | n6823 ;
  assign n6825 = x65 & n6819 ;
  assign n20954 = ~n6825 ;
  assign n6826 = n6824 & n20954 ;
  assign n20955 = ~n6826 ;
  assign n6827 = n6820 & n20955 ;
  assign n6828 = x66 & n6827 ;
  assign n6829 = n20804 & n6480 ;
  assign n6830 = n154 & n6829 ;
  assign n6831 = n6484 & n6830 ;
  assign n6832 = n6484 | n6830 ;
  assign n20956 = ~n6831 ;
  assign n6833 = n20956 & n6832 ;
  assign n6834 = x66 | n6827 ;
  assign n20957 = ~n6833 ;
  assign n6835 = n20957 & n6834 ;
  assign n6836 = n6828 | n6835 ;
  assign n6837 = x67 & n6836 ;
  assign n6838 = x67 | n6836 ;
  assign n6839 = n6487 & n20807 ;
  assign n6840 = n154 & n6839 ;
  assign n20958 = ~n6493 ;
  assign n6841 = n20958 & n6840 ;
  assign n20959 = ~n6840 ;
  assign n6842 = n6493 & n20959 ;
  assign n6843 = n6841 | n6842 ;
  assign n20960 = ~n6843 ;
  assign n6844 = n6838 & n20960 ;
  assign n6845 = n6837 | n6844 ;
  assign n6846 = x68 & n6845 ;
  assign n6847 = x68 | n6845 ;
  assign n6848 = n6496 & n20811 ;
  assign n6849 = n154 & n6848 ;
  assign n20961 = ~n6502 ;
  assign n6850 = n20961 & n6849 ;
  assign n20962 = ~n6849 ;
  assign n6851 = n6502 & n20962 ;
  assign n6852 = n6850 | n6851 ;
  assign n20963 = ~n6852 ;
  assign n6853 = n6847 & n20963 ;
  assign n6854 = n6846 | n6853 ;
  assign n6855 = x69 & n6854 ;
  assign n6856 = x69 | n6854 ;
  assign n6857 = n6505 & n20815 ;
  assign n6858 = n154 & n6857 ;
  assign n20964 = ~n6511 ;
  assign n6859 = n20964 & n6858 ;
  assign n20965 = ~n6858 ;
  assign n6860 = n6511 & n20965 ;
  assign n6861 = n6859 | n6860 ;
  assign n20966 = ~n6861 ;
  assign n6862 = n6856 & n20966 ;
  assign n6863 = n6855 | n6862 ;
  assign n6864 = x70 & n6863 ;
  assign n6865 = x70 | n6863 ;
  assign n6866 = n6514 & n20819 ;
  assign n6867 = n154 & n6866 ;
  assign n6868 = n6520 & n6867 ;
  assign n6869 = n6520 | n6867 ;
  assign n20967 = ~n6868 ;
  assign n6870 = n20967 & n6869 ;
  assign n20968 = ~n6870 ;
  assign n6871 = n6865 & n20968 ;
  assign n6872 = n6864 | n6871 ;
  assign n6873 = x71 & n6872 ;
  assign n6874 = x71 | n6872 ;
  assign n6875 = n6523 & n20823 ;
  assign n6876 = n154 & n6875 ;
  assign n6877 = n6529 & n6876 ;
  assign n6878 = n6529 | n6876 ;
  assign n20969 = ~n6877 ;
  assign n6879 = n20969 & n6878 ;
  assign n20970 = ~n6879 ;
  assign n6880 = n6874 & n20970 ;
  assign n6881 = n6873 | n6880 ;
  assign n6882 = x72 & n6881 ;
  assign n6883 = x72 | n6881 ;
  assign n6884 = n6532 & n20827 ;
  assign n6885 = n154 & n6884 ;
  assign n20971 = ~n6538 ;
  assign n6886 = n20971 & n6885 ;
  assign n20972 = ~n6885 ;
  assign n6887 = n6538 & n20972 ;
  assign n6888 = n6886 | n6887 ;
  assign n20973 = ~n6888 ;
  assign n6889 = n6883 & n20973 ;
  assign n6890 = n6882 | n6889 ;
  assign n6891 = x73 & n6890 ;
  assign n6892 = x73 | n6890 ;
  assign n6893 = n6541 & n20831 ;
  assign n6894 = n154 & n6893 ;
  assign n6895 = n6547 & n6894 ;
  assign n6896 = n6547 | n6894 ;
  assign n20974 = ~n6895 ;
  assign n6897 = n20974 & n6896 ;
  assign n20975 = ~n6897 ;
  assign n6898 = n6892 & n20975 ;
  assign n6899 = n6891 | n6898 ;
  assign n6900 = x74 & n6899 ;
  assign n6901 = x74 | n6899 ;
  assign n6902 = n6550 & n20835 ;
  assign n6903 = n154 & n6902 ;
  assign n20976 = ~n6556 ;
  assign n6904 = n20976 & n6903 ;
  assign n20977 = ~n6903 ;
  assign n6905 = n6556 & n20977 ;
  assign n6906 = n6904 | n6905 ;
  assign n20978 = ~n6906 ;
  assign n6907 = n6901 & n20978 ;
  assign n6908 = n6900 | n6907 ;
  assign n6909 = x75 & n6908 ;
  assign n6910 = x75 | n6908 ;
  assign n6911 = n6559 & n20839 ;
  assign n6912 = n154 & n6911 ;
  assign n20979 = ~n6565 ;
  assign n6913 = n20979 & n6912 ;
  assign n20980 = ~n6912 ;
  assign n6914 = n6565 & n20980 ;
  assign n6915 = n6913 | n6914 ;
  assign n20981 = ~n6915 ;
  assign n6916 = n6910 & n20981 ;
  assign n6917 = n6909 | n6916 ;
  assign n6918 = x76 & n6917 ;
  assign n6919 = x76 | n6917 ;
  assign n6920 = n6568 & n20843 ;
  assign n6921 = n154 & n6920 ;
  assign n6922 = n6574 & n6921 ;
  assign n6923 = n6574 | n6921 ;
  assign n20982 = ~n6922 ;
  assign n6924 = n20982 & n6923 ;
  assign n20983 = ~n6924 ;
  assign n6925 = n6919 & n20983 ;
  assign n6926 = n6918 | n6925 ;
  assign n6927 = x77 & n6926 ;
  assign n6928 = x77 | n6926 ;
  assign n6929 = n6577 & n20847 ;
  assign n6930 = n154 & n6929 ;
  assign n6931 = n6583 & n6930 ;
  assign n6932 = n6583 | n6930 ;
  assign n20984 = ~n6931 ;
  assign n6933 = n20984 & n6932 ;
  assign n20985 = ~n6933 ;
  assign n6934 = n6928 & n20985 ;
  assign n6935 = n6927 | n6934 ;
  assign n6936 = x78 & n6935 ;
  assign n6937 = x78 | n6935 ;
  assign n6938 = n6586 & n20851 ;
  assign n6939 = n154 & n6938 ;
  assign n6940 = n6592 & n6939 ;
  assign n6941 = n6592 | n6939 ;
  assign n20986 = ~n6940 ;
  assign n6942 = n20986 & n6941 ;
  assign n20987 = ~n6942 ;
  assign n6943 = n6937 & n20987 ;
  assign n6944 = n6936 | n6943 ;
  assign n6945 = x79 & n6944 ;
  assign n6946 = x79 | n6944 ;
  assign n6947 = n6595 & n20855 ;
  assign n6948 = n154 & n6947 ;
  assign n6949 = n6601 & n6948 ;
  assign n6950 = n6601 | n6948 ;
  assign n20988 = ~n6949 ;
  assign n6951 = n20988 & n6950 ;
  assign n20989 = ~n6951 ;
  assign n6952 = n6946 & n20989 ;
  assign n6953 = n6945 | n6952 ;
  assign n6954 = x80 & n6953 ;
  assign n6955 = x80 | n6953 ;
  assign n6956 = n6604 & n20859 ;
  assign n6957 = n154 & n6956 ;
  assign n20990 = ~n6610 ;
  assign n6958 = n20990 & n6957 ;
  assign n20991 = ~n6957 ;
  assign n6959 = n6610 & n20991 ;
  assign n6960 = n6958 | n6959 ;
  assign n20992 = ~n6960 ;
  assign n6961 = n6955 & n20992 ;
  assign n6962 = n6954 | n6961 ;
  assign n6963 = x81 & n6962 ;
  assign n6964 = x81 | n6962 ;
  assign n6965 = n6613 & n20863 ;
  assign n6966 = n154 & n6965 ;
  assign n20993 = ~n6619 ;
  assign n6967 = n20993 & n6966 ;
  assign n20994 = ~n6966 ;
  assign n6968 = n6619 & n20994 ;
  assign n6969 = n6967 | n6968 ;
  assign n20995 = ~n6969 ;
  assign n6970 = n6964 & n20995 ;
  assign n6971 = n6963 | n6970 ;
  assign n6972 = x82 & n6971 ;
  assign n6973 = x82 | n6971 ;
  assign n6974 = n6622 & n20867 ;
  assign n6975 = n154 & n6974 ;
  assign n20996 = ~n6628 ;
  assign n6976 = n20996 & n6975 ;
  assign n20997 = ~n6975 ;
  assign n6977 = n6628 & n20997 ;
  assign n6978 = n6976 | n6977 ;
  assign n20998 = ~n6978 ;
  assign n6979 = n6973 & n20998 ;
  assign n6980 = n6972 | n6979 ;
  assign n6981 = x83 & n6980 ;
  assign n6982 = x83 | n6980 ;
  assign n6983 = n6631 & n20871 ;
  assign n6984 = n154 & n6983 ;
  assign n6985 = n6637 & n6984 ;
  assign n6986 = n6637 | n6984 ;
  assign n20999 = ~n6985 ;
  assign n6987 = n20999 & n6986 ;
  assign n21000 = ~n6987 ;
  assign n6988 = n6982 & n21000 ;
  assign n6989 = n6981 | n6988 ;
  assign n6990 = x84 & n6989 ;
  assign n6991 = x84 | n6989 ;
  assign n6992 = n6640 & n20875 ;
  assign n6993 = n154 & n6992 ;
  assign n6994 = n6646 & n6993 ;
  assign n6995 = n6646 | n6993 ;
  assign n21001 = ~n6994 ;
  assign n6996 = n21001 & n6995 ;
  assign n21002 = ~n6996 ;
  assign n6997 = n6991 & n21002 ;
  assign n6998 = n6990 | n6997 ;
  assign n6999 = x85 & n6998 ;
  assign n7000 = x85 | n6998 ;
  assign n7001 = n6649 & n20879 ;
  assign n7002 = n154 & n7001 ;
  assign n7003 = n6655 & n7002 ;
  assign n7004 = n6655 | n7002 ;
  assign n21003 = ~n7003 ;
  assign n7005 = n21003 & n7004 ;
  assign n21004 = ~n7005 ;
  assign n7006 = n7000 & n21004 ;
  assign n7007 = n6999 | n7006 ;
  assign n7008 = x86 & n7007 ;
  assign n7009 = x86 | n7007 ;
  assign n7010 = n6658 & n20883 ;
  assign n7011 = n154 & n7010 ;
  assign n21005 = ~n6664 ;
  assign n7012 = n21005 & n7011 ;
  assign n21006 = ~n7011 ;
  assign n7013 = n6664 & n21006 ;
  assign n7014 = n7012 | n7013 ;
  assign n21007 = ~n7014 ;
  assign n7015 = n7009 & n21007 ;
  assign n7016 = n7008 | n7015 ;
  assign n7017 = x87 & n7016 ;
  assign n7018 = x87 | n7016 ;
  assign n7019 = n6667 & n20887 ;
  assign n7020 = n154 & n7019 ;
  assign n21008 = ~n6673 ;
  assign n7021 = n21008 & n7020 ;
  assign n21009 = ~n7020 ;
  assign n7022 = n6673 & n21009 ;
  assign n7023 = n7021 | n7022 ;
  assign n21010 = ~n7023 ;
  assign n7024 = n7018 & n21010 ;
  assign n7025 = n7017 | n7024 ;
  assign n7026 = x88 & n7025 ;
  assign n7027 = x88 | n7025 ;
  assign n7028 = n6676 & n20891 ;
  assign n7029 = n154 & n7028 ;
  assign n21011 = ~n6682 ;
  assign n7030 = n21011 & n7029 ;
  assign n21012 = ~n7029 ;
  assign n7031 = n6682 & n21012 ;
  assign n7032 = n7030 | n7031 ;
  assign n21013 = ~n7032 ;
  assign n7033 = n7027 & n21013 ;
  assign n7034 = n7026 | n7033 ;
  assign n7035 = x89 & n7034 ;
  assign n7036 = x89 | n7034 ;
  assign n7037 = n6685 & n20895 ;
  assign n7038 = n154 & n7037 ;
  assign n21014 = ~n6691 ;
  assign n7039 = n21014 & n7038 ;
  assign n21015 = ~n7038 ;
  assign n7040 = n6691 & n21015 ;
  assign n7041 = n7039 | n7040 ;
  assign n21016 = ~n7041 ;
  assign n7042 = n7036 & n21016 ;
  assign n7043 = n7035 | n7042 ;
  assign n7044 = x90 & n7043 ;
  assign n7045 = x90 | n7043 ;
  assign n7046 = n6694 & n20899 ;
  assign n7047 = n154 & n7046 ;
  assign n21017 = ~n6700 ;
  assign n7048 = n21017 & n7047 ;
  assign n21018 = ~n7047 ;
  assign n7049 = n6700 & n21018 ;
  assign n7050 = n7048 | n7049 ;
  assign n21019 = ~n7050 ;
  assign n7051 = n7045 & n21019 ;
  assign n7052 = n7044 | n7051 ;
  assign n7053 = x91 & n7052 ;
  assign n7054 = x91 | n7052 ;
  assign n7055 = n6703 & n20903 ;
  assign n7056 = n154 & n7055 ;
  assign n21020 = ~n6709 ;
  assign n7057 = n21020 & n7056 ;
  assign n21021 = ~n7056 ;
  assign n7058 = n6709 & n21021 ;
  assign n7059 = n7057 | n7058 ;
  assign n21022 = ~n7059 ;
  assign n7060 = n7054 & n21022 ;
  assign n7061 = n7053 | n7060 ;
  assign n7062 = x92 & n7061 ;
  assign n7063 = x92 | n7061 ;
  assign n7064 = n6712 & n20907 ;
  assign n7065 = n154 & n7064 ;
  assign n21023 = ~n6718 ;
  assign n7066 = n21023 & n7065 ;
  assign n21024 = ~n7065 ;
  assign n7067 = n6718 & n21024 ;
  assign n7068 = n7066 | n7067 ;
  assign n21025 = ~n7068 ;
  assign n7069 = n7063 & n21025 ;
  assign n7070 = n7062 | n7069 ;
  assign n7071 = x93 & n7070 ;
  assign n7072 = x93 | n7070 ;
  assign n7073 = n6721 & n20911 ;
  assign n7074 = n154 & n7073 ;
  assign n21026 = ~n6727 ;
  assign n7075 = n21026 & n7074 ;
  assign n21027 = ~n7074 ;
  assign n7076 = n6727 & n21027 ;
  assign n7077 = n7075 | n7076 ;
  assign n21028 = ~n7077 ;
  assign n7078 = n7072 & n21028 ;
  assign n7079 = n7071 | n7078 ;
  assign n7080 = x94 & n7079 ;
  assign n7081 = x94 | n7079 ;
  assign n7082 = n6730 & n20915 ;
  assign n7083 = n154 & n7082 ;
  assign n21029 = ~n6736 ;
  assign n7084 = n21029 & n7083 ;
  assign n21030 = ~n7083 ;
  assign n7085 = n6736 & n21030 ;
  assign n7086 = n7084 | n7085 ;
  assign n21031 = ~n7086 ;
  assign n7087 = n7081 & n21031 ;
  assign n7088 = n7080 | n7087 ;
  assign n7089 = x95 & n7088 ;
  assign n7090 = x95 | n7088 ;
  assign n7091 = n6739 & n20919 ;
  assign n7092 = n154 & n7091 ;
  assign n21032 = ~n6745 ;
  assign n7093 = n21032 & n7092 ;
  assign n21033 = ~n7092 ;
  assign n7094 = n6745 & n21033 ;
  assign n7095 = n7093 | n7094 ;
  assign n21034 = ~n7095 ;
  assign n7096 = n7090 & n21034 ;
  assign n7097 = n7089 | n7096 ;
  assign n7098 = x96 & n7097 ;
  assign n7099 = x96 | n7097 ;
  assign n7100 = n6748 & n20923 ;
  assign n7101 = n154 & n7100 ;
  assign n21035 = ~n6754 ;
  assign n7102 = n21035 & n7101 ;
  assign n21036 = ~n7101 ;
  assign n7103 = n6754 & n21036 ;
  assign n7104 = n7102 | n7103 ;
  assign n21037 = ~n7104 ;
  assign n7105 = n7099 & n21037 ;
  assign n7106 = n7098 | n7105 ;
  assign n7107 = x97 & n7106 ;
  assign n7108 = x97 | n7106 ;
  assign n7109 = n6757 & n20927 ;
  assign n7110 = n154 & n7109 ;
  assign n21038 = ~n6763 ;
  assign n7111 = n21038 & n7110 ;
  assign n21039 = ~n7110 ;
  assign n7112 = n6763 & n21039 ;
  assign n7113 = n7111 | n7112 ;
  assign n21040 = ~n7113 ;
  assign n7114 = n7108 & n21040 ;
  assign n7115 = n7107 | n7114 ;
  assign n7116 = x98 & n7115 ;
  assign n7117 = x98 | n7115 ;
  assign n7118 = n6766 & n20931 ;
  assign n7119 = n154 & n7118 ;
  assign n21041 = ~n6772 ;
  assign n7120 = n21041 & n7119 ;
  assign n21042 = ~n7119 ;
  assign n7121 = n6772 & n21042 ;
  assign n7122 = n7120 | n7121 ;
  assign n21043 = ~n7122 ;
  assign n7123 = n7117 & n21043 ;
  assign n7124 = n7116 | n7123 ;
  assign n7125 = x99 & n7124 ;
  assign n7126 = x99 | n7124 ;
  assign n7127 = n6775 & n20935 ;
  assign n7128 = n154 & n7127 ;
  assign n21044 = ~n6781 ;
  assign n7129 = n21044 & n7128 ;
  assign n21045 = ~n7128 ;
  assign n7130 = n6781 & n21045 ;
  assign n7131 = n7129 | n7130 ;
  assign n21046 = ~n7131 ;
  assign n7132 = n7126 & n21046 ;
  assign n7133 = n7125 | n7132 ;
  assign n7134 = x100 & n7133 ;
  assign n7135 = x100 | n7133 ;
  assign n7136 = n6784 & n20939 ;
  assign n7137 = n154 & n7136 ;
  assign n21047 = ~n6790 ;
  assign n7138 = n21047 & n7137 ;
  assign n21048 = ~n7137 ;
  assign n7139 = n6790 & n21048 ;
  assign n7140 = n7138 | n7139 ;
  assign n21049 = ~n7140 ;
  assign n7141 = n7135 & n21049 ;
  assign n7142 = n7134 | n7141 ;
  assign n7143 = x101 & n7142 ;
  assign n7144 = x101 | n7142 ;
  assign n7145 = n6793 & n20943 ;
  assign n7146 = n154 & n7145 ;
  assign n7147 = n6799 & n7146 ;
  assign n7148 = n6799 | n7146 ;
  assign n21050 = ~n7147 ;
  assign n7149 = n21050 & n7148 ;
  assign n21051 = ~n7149 ;
  assign n7150 = n7144 & n21051 ;
  assign n7151 = n7143 | n7150 ;
  assign n7152 = x102 & n7151 ;
  assign n7153 = x102 | n7151 ;
  assign n21052 = ~n6815 ;
  assign n7154 = n21052 & n7153 ;
  assign n7155 = n7152 | n7154 ;
  assign n21053 = ~n7155 ;
  assign n7156 = n6818 & n21053 ;
  assign n21054 = ~n7156 ;
  assign n7157 = x103 & n21054 ;
  assign n7158 = n18378 | n7157 ;
  assign n21055 = ~n6818 ;
  assign n7160 = n21055 & n7155 ;
  assign n7161 = n7158 | n7160 ;
  assign n21056 = ~n7152 ;
  assign n7162 = n21056 & n7153 ;
  assign n153 = ~n7161 ;
  assign n7163 = n153 & n7162 ;
  assign n7164 = n6815 & n7163 ;
  assign n7165 = n6815 | n7163 ;
  assign n21058 = ~n7164 ;
  assign n7166 = n21058 & n7165 ;
  assign n7159 = n6816 & n7158 ;
  assign n7167 = n21884 | n7159 ;
  assign n21059 = ~x23 ;
  assign n7168 = n21059 & x64 ;
  assign n7170 = x65 | n7168 ;
  assign n7169 = x65 & n7168 ;
  assign n7171 = x64 & n153 ;
  assign n7172 = x24 & n7171 ;
  assign n7173 = x24 | n7171 ;
  assign n21060 = ~n7172 ;
  assign n7174 = n21060 & n7173 ;
  assign n21061 = ~n7169 ;
  assign n7175 = n21061 & n7174 ;
  assign n21062 = ~n7175 ;
  assign n7176 = n7170 & n21062 ;
  assign n7177 = x66 | n7176 ;
  assign n7178 = x66 & n7176 ;
  assign n7179 = n6820 & n153 ;
  assign n7180 = n20954 & n7179 ;
  assign n7181 = n6824 | n7180 ;
  assign n7182 = n6826 & n7179 ;
  assign n21063 = ~n7182 ;
  assign n7183 = n7181 & n21063 ;
  assign n21064 = ~n7178 ;
  assign n7184 = n21064 & n7183 ;
  assign n21065 = ~n7184 ;
  assign n7185 = n7177 & n21065 ;
  assign n7186 = x67 | n7185 ;
  assign n7187 = x67 & n7185 ;
  assign n21066 = ~n6828 ;
  assign n7188 = n21066 & n6834 ;
  assign n7189 = n153 & n7188 ;
  assign n7190 = n6833 & n7189 ;
  assign n7191 = n6833 | n7189 ;
  assign n21067 = ~n7190 ;
  assign n7192 = n21067 & n7191 ;
  assign n21068 = ~n7187 ;
  assign n7193 = n21068 & n7192 ;
  assign n21069 = ~n7193 ;
  assign n7194 = n7186 & n21069 ;
  assign n7195 = x68 | n7194 ;
  assign n7196 = x68 & n7194 ;
  assign n21070 = ~n6837 ;
  assign n7197 = n21070 & n6838 ;
  assign n7198 = n153 & n7197 ;
  assign n7199 = n6843 & n7198 ;
  assign n7200 = n6843 | n7198 ;
  assign n21071 = ~n7199 ;
  assign n7201 = n21071 & n7200 ;
  assign n21072 = ~n7196 ;
  assign n7202 = n21072 & n7201 ;
  assign n21073 = ~n7202 ;
  assign n7203 = n7195 & n21073 ;
  assign n7204 = x69 | n7203 ;
  assign n7205 = x69 & n7203 ;
  assign n21074 = ~n6846 ;
  assign n7206 = n21074 & n6847 ;
  assign n7207 = n153 & n7206 ;
  assign n7208 = n6852 & n7207 ;
  assign n7209 = n6852 | n7207 ;
  assign n21075 = ~n7208 ;
  assign n7210 = n21075 & n7209 ;
  assign n21076 = ~n7205 ;
  assign n7211 = n21076 & n7210 ;
  assign n21077 = ~n7211 ;
  assign n7212 = n7204 & n21077 ;
  assign n7213 = x70 | n7212 ;
  assign n7214 = x70 & n7212 ;
  assign n21078 = ~n6855 ;
  assign n7215 = n21078 & n6856 ;
  assign n7216 = n153 & n7215 ;
  assign n7217 = n6861 & n7216 ;
  assign n7218 = n6861 | n7216 ;
  assign n21079 = ~n7217 ;
  assign n7219 = n21079 & n7218 ;
  assign n21080 = ~n7214 ;
  assign n7220 = n21080 & n7219 ;
  assign n21081 = ~n7220 ;
  assign n7221 = n7213 & n21081 ;
  assign n7222 = x71 | n7221 ;
  assign n7223 = x71 & n7221 ;
  assign n21082 = ~n6864 ;
  assign n7224 = n21082 & n6865 ;
  assign n7225 = n153 & n7224 ;
  assign n7226 = n6870 & n7225 ;
  assign n7227 = n6870 | n7225 ;
  assign n21083 = ~n7226 ;
  assign n7228 = n21083 & n7227 ;
  assign n21084 = ~n7223 ;
  assign n7229 = n21084 & n7228 ;
  assign n21085 = ~n7229 ;
  assign n7230 = n7222 & n21085 ;
  assign n7231 = x72 | n7230 ;
  assign n7232 = x72 & n7230 ;
  assign n21086 = ~n6873 ;
  assign n7233 = n21086 & n6874 ;
  assign n7234 = n153 & n7233 ;
  assign n7235 = n6879 & n7234 ;
  assign n7236 = n6879 | n7234 ;
  assign n21087 = ~n7235 ;
  assign n7237 = n21087 & n7236 ;
  assign n21088 = ~n7232 ;
  assign n7238 = n21088 & n7237 ;
  assign n21089 = ~n7238 ;
  assign n7239 = n7231 & n21089 ;
  assign n7240 = x73 | n7239 ;
  assign n7241 = x73 & n7239 ;
  assign n21090 = ~n6882 ;
  assign n7242 = n21090 & n6883 ;
  assign n7243 = n153 & n7242 ;
  assign n7244 = n20973 & n7243 ;
  assign n21091 = ~n7243 ;
  assign n7245 = n6888 & n21091 ;
  assign n7246 = n7244 | n7245 ;
  assign n21092 = ~n7241 ;
  assign n7247 = n21092 & n7246 ;
  assign n21093 = ~n7247 ;
  assign n7248 = n7240 & n21093 ;
  assign n7249 = x74 | n7248 ;
  assign n7250 = x74 & n7248 ;
  assign n21094 = ~n6891 ;
  assign n7251 = n21094 & n6892 ;
  assign n7252 = n153 & n7251 ;
  assign n7253 = n6897 & n7252 ;
  assign n7254 = n6897 | n7252 ;
  assign n21095 = ~n7253 ;
  assign n7255 = n21095 & n7254 ;
  assign n21096 = ~n7250 ;
  assign n7256 = n21096 & n7255 ;
  assign n21097 = ~n7256 ;
  assign n7257 = n7249 & n21097 ;
  assign n7258 = x75 | n7257 ;
  assign n7259 = x75 & n7257 ;
  assign n21098 = ~n6900 ;
  assign n7260 = n21098 & n6901 ;
  assign n7261 = n153 & n7260 ;
  assign n7262 = n6906 & n7261 ;
  assign n7263 = n6906 | n7261 ;
  assign n21099 = ~n7262 ;
  assign n7264 = n21099 & n7263 ;
  assign n21100 = ~n7259 ;
  assign n7265 = n21100 & n7264 ;
  assign n21101 = ~n7265 ;
  assign n7266 = n7258 & n21101 ;
  assign n7267 = x76 | n7266 ;
  assign n7268 = x76 & n7266 ;
  assign n21102 = ~n6909 ;
  assign n7269 = n21102 & n6910 ;
  assign n7270 = n153 & n7269 ;
  assign n7271 = n6915 & n7270 ;
  assign n7272 = n6915 | n7270 ;
  assign n21103 = ~n7271 ;
  assign n7273 = n21103 & n7272 ;
  assign n21104 = ~n7268 ;
  assign n7274 = n21104 & n7273 ;
  assign n21105 = ~n7274 ;
  assign n7275 = n7267 & n21105 ;
  assign n7276 = x77 | n7275 ;
  assign n7277 = x77 & n7275 ;
  assign n21106 = ~n6918 ;
  assign n7278 = n21106 & n6919 ;
  assign n7279 = n153 & n7278 ;
  assign n7280 = n6924 & n7279 ;
  assign n7281 = n6924 | n7279 ;
  assign n21107 = ~n7280 ;
  assign n7282 = n21107 & n7281 ;
  assign n21108 = ~n7277 ;
  assign n7283 = n21108 & n7282 ;
  assign n21109 = ~n7283 ;
  assign n7284 = n7276 & n21109 ;
  assign n7285 = x78 | n7284 ;
  assign n7286 = x78 & n7284 ;
  assign n21110 = ~n6927 ;
  assign n7287 = n21110 & n6928 ;
  assign n7288 = n153 & n7287 ;
  assign n7289 = n6933 & n7288 ;
  assign n7290 = n6933 | n7288 ;
  assign n21111 = ~n7289 ;
  assign n7291 = n21111 & n7290 ;
  assign n21112 = ~n7286 ;
  assign n7292 = n21112 & n7291 ;
  assign n21113 = ~n7292 ;
  assign n7293 = n7285 & n21113 ;
  assign n7294 = x79 | n7293 ;
  assign n7295 = x79 & n7293 ;
  assign n21114 = ~n6936 ;
  assign n7296 = n21114 & n6937 ;
  assign n7297 = n153 & n7296 ;
  assign n7298 = n6942 & n7297 ;
  assign n7299 = n6942 | n7297 ;
  assign n21115 = ~n7298 ;
  assign n7300 = n21115 & n7299 ;
  assign n21116 = ~n7295 ;
  assign n7301 = n21116 & n7300 ;
  assign n21117 = ~n7301 ;
  assign n7302 = n7294 & n21117 ;
  assign n7303 = x80 | n7302 ;
  assign n7304 = x80 & n7302 ;
  assign n21118 = ~n6945 ;
  assign n7305 = n21118 & n6946 ;
  assign n7306 = n153 & n7305 ;
  assign n7307 = n6951 & n7306 ;
  assign n7308 = n6951 | n7306 ;
  assign n21119 = ~n7307 ;
  assign n7309 = n21119 & n7308 ;
  assign n21120 = ~n7304 ;
  assign n7310 = n21120 & n7309 ;
  assign n21121 = ~n7310 ;
  assign n7311 = n7303 & n21121 ;
  assign n7312 = x81 | n7311 ;
  assign n7313 = x81 & n7311 ;
  assign n21122 = ~n6954 ;
  assign n7314 = n21122 & n6955 ;
  assign n7315 = n153 & n7314 ;
  assign n7316 = n6960 & n7315 ;
  assign n7317 = n6960 | n7315 ;
  assign n21123 = ~n7316 ;
  assign n7318 = n21123 & n7317 ;
  assign n21124 = ~n7313 ;
  assign n7319 = n21124 & n7318 ;
  assign n21125 = ~n7319 ;
  assign n7320 = n7312 & n21125 ;
  assign n7321 = x82 | n7320 ;
  assign n7322 = x82 & n7320 ;
  assign n21126 = ~n6963 ;
  assign n7323 = n21126 & n6964 ;
  assign n7324 = n153 & n7323 ;
  assign n7325 = n20995 & n7324 ;
  assign n21127 = ~n7324 ;
  assign n7326 = n6969 & n21127 ;
  assign n7327 = n7325 | n7326 ;
  assign n21128 = ~n7322 ;
  assign n7328 = n21128 & n7327 ;
  assign n21129 = ~n7328 ;
  assign n7329 = n7321 & n21129 ;
  assign n7330 = x83 | n7329 ;
  assign n7331 = x83 & n7329 ;
  assign n21130 = ~n6972 ;
  assign n7332 = n21130 & n6973 ;
  assign n7333 = n153 & n7332 ;
  assign n7334 = n6978 & n7333 ;
  assign n7335 = n6978 | n7333 ;
  assign n21131 = ~n7334 ;
  assign n7336 = n21131 & n7335 ;
  assign n21132 = ~n7331 ;
  assign n7337 = n21132 & n7336 ;
  assign n21133 = ~n7337 ;
  assign n7338 = n7330 & n21133 ;
  assign n7339 = x84 | n7338 ;
  assign n7340 = x84 & n7338 ;
  assign n21134 = ~n6981 ;
  assign n7341 = n21134 & n6982 ;
  assign n7342 = n153 & n7341 ;
  assign n7343 = n6987 & n7342 ;
  assign n7344 = n6987 | n7342 ;
  assign n21135 = ~n7343 ;
  assign n7345 = n21135 & n7344 ;
  assign n21136 = ~n7340 ;
  assign n7346 = n21136 & n7345 ;
  assign n21137 = ~n7346 ;
  assign n7347 = n7339 & n21137 ;
  assign n7348 = x85 | n7347 ;
  assign n7349 = x85 & n7347 ;
  assign n21138 = ~n6990 ;
  assign n7350 = n21138 & n6991 ;
  assign n7351 = n153 & n7350 ;
  assign n7352 = n6996 & n7351 ;
  assign n7353 = n6996 | n7351 ;
  assign n21139 = ~n7352 ;
  assign n7354 = n21139 & n7353 ;
  assign n21140 = ~n7349 ;
  assign n7355 = n21140 & n7354 ;
  assign n21141 = ~n7355 ;
  assign n7356 = n7348 & n21141 ;
  assign n7357 = x86 | n7356 ;
  assign n7358 = x86 & n7356 ;
  assign n21142 = ~n6999 ;
  assign n7359 = n21142 & n7000 ;
  assign n7360 = n153 & n7359 ;
  assign n7361 = n7005 & n7360 ;
  assign n7362 = n7005 | n7360 ;
  assign n21143 = ~n7361 ;
  assign n7363 = n21143 & n7362 ;
  assign n21144 = ~n7358 ;
  assign n7364 = n21144 & n7363 ;
  assign n21145 = ~n7364 ;
  assign n7365 = n7357 & n21145 ;
  assign n7366 = x87 | n7365 ;
  assign n7367 = x87 & n7365 ;
  assign n21146 = ~n7008 ;
  assign n7368 = n21146 & n7009 ;
  assign n7369 = n153 & n7368 ;
  assign n7370 = n21007 & n7369 ;
  assign n21147 = ~n7369 ;
  assign n7371 = n7014 & n21147 ;
  assign n7372 = n7370 | n7371 ;
  assign n21148 = ~n7367 ;
  assign n7373 = n21148 & n7372 ;
  assign n21149 = ~n7373 ;
  assign n7374 = n7366 & n21149 ;
  assign n7375 = x88 | n7374 ;
  assign n7376 = x88 & n7374 ;
  assign n21150 = ~n7017 ;
  assign n7377 = n21150 & n7018 ;
  assign n7378 = n153 & n7377 ;
  assign n7379 = n21010 & n7378 ;
  assign n21151 = ~n7378 ;
  assign n7380 = n7023 & n21151 ;
  assign n7381 = n7379 | n7380 ;
  assign n21152 = ~n7376 ;
  assign n7382 = n21152 & n7381 ;
  assign n21153 = ~n7382 ;
  assign n7383 = n7375 & n21153 ;
  assign n7384 = x89 | n7383 ;
  assign n7385 = x89 & n7383 ;
  assign n21154 = ~n7026 ;
  assign n7386 = n21154 & n7027 ;
  assign n7387 = n153 & n7386 ;
  assign n7388 = n7032 & n7387 ;
  assign n7389 = n7032 | n7387 ;
  assign n21155 = ~n7388 ;
  assign n7390 = n21155 & n7389 ;
  assign n21156 = ~n7385 ;
  assign n7391 = n21156 & n7390 ;
  assign n21157 = ~n7391 ;
  assign n7392 = n7384 & n21157 ;
  assign n7393 = x90 | n7392 ;
  assign n7394 = x90 & n7392 ;
  assign n21158 = ~n7035 ;
  assign n7395 = n21158 & n7036 ;
  assign n7396 = n153 & n7395 ;
  assign n7397 = n21016 & n7396 ;
  assign n21159 = ~n7396 ;
  assign n7398 = n7041 & n21159 ;
  assign n7399 = n7397 | n7398 ;
  assign n21160 = ~n7394 ;
  assign n7400 = n21160 & n7399 ;
  assign n21161 = ~n7400 ;
  assign n7401 = n7393 & n21161 ;
  assign n7402 = x91 | n7401 ;
  assign n7403 = x91 & n7401 ;
  assign n21162 = ~n7044 ;
  assign n7404 = n21162 & n7045 ;
  assign n7405 = n153 & n7404 ;
  assign n7406 = n21019 & n7405 ;
  assign n21163 = ~n7405 ;
  assign n7407 = n7050 & n21163 ;
  assign n7408 = n7406 | n7407 ;
  assign n21164 = ~n7403 ;
  assign n7409 = n21164 & n7408 ;
  assign n21165 = ~n7409 ;
  assign n7410 = n7402 & n21165 ;
  assign n7411 = x92 | n7410 ;
  assign n7412 = x92 & n7410 ;
  assign n21166 = ~n7053 ;
  assign n7413 = n21166 & n7054 ;
  assign n7414 = n153 & n7413 ;
  assign n7415 = n7059 & n7414 ;
  assign n7416 = n7059 | n7414 ;
  assign n21167 = ~n7415 ;
  assign n7417 = n21167 & n7416 ;
  assign n21168 = ~n7412 ;
  assign n7418 = n21168 & n7417 ;
  assign n21169 = ~n7418 ;
  assign n7419 = n7411 & n21169 ;
  assign n7420 = x93 | n7419 ;
  assign n7421 = x93 & n7419 ;
  assign n21170 = ~n7062 ;
  assign n7422 = n21170 & n7063 ;
  assign n7423 = n153 & n7422 ;
  assign n7424 = n7068 & n7423 ;
  assign n7425 = n7068 | n7423 ;
  assign n21171 = ~n7424 ;
  assign n7426 = n21171 & n7425 ;
  assign n21172 = ~n7421 ;
  assign n7427 = n21172 & n7426 ;
  assign n21173 = ~n7427 ;
  assign n7428 = n7420 & n21173 ;
  assign n7429 = x94 | n7428 ;
  assign n7430 = x94 & n7428 ;
  assign n21174 = ~n7071 ;
  assign n7431 = n21174 & n7072 ;
  assign n7432 = n153 & n7431 ;
  assign n7433 = n21028 & n7432 ;
  assign n21175 = ~n7432 ;
  assign n7434 = n7077 & n21175 ;
  assign n7435 = n7433 | n7434 ;
  assign n21176 = ~n7430 ;
  assign n7436 = n21176 & n7435 ;
  assign n21177 = ~n7436 ;
  assign n7437 = n7429 & n21177 ;
  assign n7438 = x95 | n7437 ;
  assign n7439 = x95 & n7437 ;
  assign n21178 = ~n7080 ;
  assign n7440 = n21178 & n7081 ;
  assign n7441 = n153 & n7440 ;
  assign n7442 = n7086 & n7441 ;
  assign n7443 = n7086 | n7441 ;
  assign n21179 = ~n7442 ;
  assign n7444 = n21179 & n7443 ;
  assign n21180 = ~n7439 ;
  assign n7445 = n21180 & n7444 ;
  assign n21181 = ~n7445 ;
  assign n7446 = n7438 & n21181 ;
  assign n7447 = x96 | n7446 ;
  assign n7448 = x96 & n7446 ;
  assign n21182 = ~n7089 ;
  assign n7449 = n21182 & n7090 ;
  assign n7450 = n153 & n7449 ;
  assign n7451 = n21034 & n7450 ;
  assign n21183 = ~n7450 ;
  assign n7452 = n7095 & n21183 ;
  assign n7453 = n7451 | n7452 ;
  assign n21184 = ~n7448 ;
  assign n7454 = n21184 & n7453 ;
  assign n21185 = ~n7454 ;
  assign n7455 = n7447 & n21185 ;
  assign n7456 = x97 | n7455 ;
  assign n7457 = x97 & n7455 ;
  assign n21186 = ~n7098 ;
  assign n7458 = n21186 & n7099 ;
  assign n7459 = n153 & n7458 ;
  assign n7460 = n21037 & n7459 ;
  assign n21187 = ~n7459 ;
  assign n7461 = n7104 & n21187 ;
  assign n7462 = n7460 | n7461 ;
  assign n21188 = ~n7457 ;
  assign n7463 = n21188 & n7462 ;
  assign n21189 = ~n7463 ;
  assign n7464 = n7456 & n21189 ;
  assign n7465 = x98 | n7464 ;
  assign n7466 = x98 & n7464 ;
  assign n21190 = ~n7107 ;
  assign n7467 = n21190 & n7108 ;
  assign n7468 = n153 & n7467 ;
  assign n7469 = n7113 & n7468 ;
  assign n7470 = n7113 | n7468 ;
  assign n21191 = ~n7469 ;
  assign n7471 = n21191 & n7470 ;
  assign n21192 = ~n7466 ;
  assign n7472 = n21192 & n7471 ;
  assign n21193 = ~n7472 ;
  assign n7473 = n7465 & n21193 ;
  assign n7474 = x99 | n7473 ;
  assign n7475 = x99 & n7473 ;
  assign n21194 = ~n7116 ;
  assign n7476 = n21194 & n7117 ;
  assign n7477 = n153 & n7476 ;
  assign n7478 = n7122 & n7477 ;
  assign n7479 = n7122 | n7477 ;
  assign n21195 = ~n7478 ;
  assign n7480 = n21195 & n7479 ;
  assign n21196 = ~n7475 ;
  assign n7481 = n21196 & n7480 ;
  assign n21197 = ~n7481 ;
  assign n7482 = n7474 & n21197 ;
  assign n7483 = x100 | n7482 ;
  assign n7484 = x100 & n7482 ;
  assign n21198 = ~n7125 ;
  assign n7485 = n21198 & n7126 ;
  assign n7486 = n153 & n7485 ;
  assign n7487 = n7131 & n7486 ;
  assign n7488 = n7131 | n7486 ;
  assign n21199 = ~n7487 ;
  assign n7489 = n21199 & n7488 ;
  assign n21200 = ~n7484 ;
  assign n7490 = n21200 & n7489 ;
  assign n21201 = ~n7490 ;
  assign n7491 = n7483 & n21201 ;
  assign n7492 = x101 | n7491 ;
  assign n7493 = x101 & n7491 ;
  assign n21202 = ~n7134 ;
  assign n7494 = n21202 & n7135 ;
  assign n7495 = n153 & n7494 ;
  assign n7496 = n7140 & n7495 ;
  assign n7497 = n7140 | n7495 ;
  assign n21203 = ~n7496 ;
  assign n7498 = n21203 & n7497 ;
  assign n21204 = ~n7493 ;
  assign n7499 = n21204 & n7498 ;
  assign n21205 = ~n7499 ;
  assign n7500 = n7492 & n21205 ;
  assign n7501 = x102 | n7500 ;
  assign n7502 = x102 & n7500 ;
  assign n21206 = ~n7143 ;
  assign n7503 = n21206 & n7144 ;
  assign n7504 = n153 & n7503 ;
  assign n7505 = n7149 & n7504 ;
  assign n7506 = n7149 | n7504 ;
  assign n21207 = ~n7505 ;
  assign n7507 = n21207 & n7506 ;
  assign n21208 = ~n7502 ;
  assign n7508 = n21208 & n7507 ;
  assign n21209 = ~n7508 ;
  assign n7509 = n7501 & n21209 ;
  assign n7511 = x103 | n7509 ;
  assign n7512 = x103 & n7509 ;
  assign n21210 = ~n7512 ;
  assign n7513 = n7166 & n21210 ;
  assign n21211 = ~n7513 ;
  assign n7514 = n7511 & n21211 ;
  assign n21212 = ~n7514 ;
  assign n7515 = n7167 & n21212 ;
  assign n21213 = ~n7515 ;
  assign n7516 = x104 & n21213 ;
  assign n7517 = n18373 | n7516 ;
  assign n21214 = ~n7167 ;
  assign n7519 = n21214 & n7514 ;
  assign n7520 = n7517 | n7519 ;
  assign n21215 = ~n7509 ;
  assign n7510 = x103 & n21215 ;
  assign n21216 = ~x103 ;
  assign n7521 = n21216 & n7509 ;
  assign n7522 = n7510 | n7521 ;
  assign n152 = ~n7520 ;
  assign n7523 = n152 & n7522 ;
  assign n21218 = ~n7166 ;
  assign n7524 = n21218 & n7523 ;
  assign n21219 = ~n7523 ;
  assign n7525 = n7166 & n21219 ;
  assign n7526 = n7524 | n7525 ;
  assign n21220 = ~x22 ;
  assign n7527 = n21220 & x64 ;
  assign n7529 = x65 | n7527 ;
  assign n7528 = x65 & n7527 ;
  assign n7530 = x64 & n152 ;
  assign n7531 = x23 & n7530 ;
  assign n7532 = x23 | n7530 ;
  assign n21221 = ~n7531 ;
  assign n7533 = n21221 & n7532 ;
  assign n21222 = ~n7528 ;
  assign n7534 = n21222 & n7533 ;
  assign n21223 = ~n7534 ;
  assign n7535 = n7529 & n21223 ;
  assign n7536 = x66 & n7535 ;
  assign n7537 = x66 | n7535 ;
  assign n7538 = n21061 & n7170 ;
  assign n7539 = n152 & n7538 ;
  assign n7540 = n7174 & n7539 ;
  assign n7541 = n7174 | n7539 ;
  assign n21224 = ~n7540 ;
  assign n7542 = n21224 & n7541 ;
  assign n21225 = ~n7542 ;
  assign n7543 = n7537 & n21225 ;
  assign n7544 = n7536 | n7543 ;
  assign n7545 = x67 & n7544 ;
  assign n7546 = x67 | n7544 ;
  assign n7547 = n7177 & n21064 ;
  assign n7548 = n152 & n7547 ;
  assign n7549 = n7183 | n7548 ;
  assign n7550 = n7183 & n7548 ;
  assign n21226 = ~n7550 ;
  assign n7551 = n7549 & n21226 ;
  assign n21227 = ~n7551 ;
  assign n7552 = n7546 & n21227 ;
  assign n7553 = n7545 | n7552 ;
  assign n7554 = x68 & n7553 ;
  assign n7555 = x68 | n7553 ;
  assign n7556 = n7186 & n21068 ;
  assign n7557 = n152 & n7556 ;
  assign n21228 = ~n7192 ;
  assign n7558 = n21228 & n7557 ;
  assign n21229 = ~n7557 ;
  assign n7559 = n7192 & n21229 ;
  assign n7560 = n7558 | n7559 ;
  assign n21230 = ~n7560 ;
  assign n7561 = n7555 & n21230 ;
  assign n7562 = n7554 | n7561 ;
  assign n7563 = x69 & n7562 ;
  assign n7564 = x69 | n7562 ;
  assign n7565 = n7195 & n21072 ;
  assign n7566 = n152 & n7565 ;
  assign n21231 = ~n7201 ;
  assign n7567 = n21231 & n7566 ;
  assign n21232 = ~n7566 ;
  assign n7568 = n7201 & n21232 ;
  assign n7569 = n7567 | n7568 ;
  assign n21233 = ~n7569 ;
  assign n7570 = n7564 & n21233 ;
  assign n7571 = n7563 | n7570 ;
  assign n7572 = x70 & n7571 ;
  assign n7573 = x70 | n7571 ;
  assign n7574 = n7204 & n21076 ;
  assign n7575 = n152 & n7574 ;
  assign n7576 = n7210 & n7575 ;
  assign n7577 = n7210 | n7575 ;
  assign n21234 = ~n7576 ;
  assign n7578 = n21234 & n7577 ;
  assign n21235 = ~n7578 ;
  assign n7579 = n7573 & n21235 ;
  assign n7580 = n7572 | n7579 ;
  assign n7581 = x71 & n7580 ;
  assign n7582 = x71 | n7580 ;
  assign n7583 = n7213 & n21080 ;
  assign n7584 = n152 & n7583 ;
  assign n7585 = n7219 & n7584 ;
  assign n7586 = n7219 | n7584 ;
  assign n21236 = ~n7585 ;
  assign n7587 = n21236 & n7586 ;
  assign n21237 = ~n7587 ;
  assign n7588 = n7582 & n21237 ;
  assign n7589 = n7581 | n7588 ;
  assign n7590 = x72 & n7589 ;
  assign n7591 = x72 | n7589 ;
  assign n7592 = n7222 & n21084 ;
  assign n7593 = n152 & n7592 ;
  assign n21238 = ~n7228 ;
  assign n7594 = n21238 & n7593 ;
  assign n21239 = ~n7593 ;
  assign n7595 = n7228 & n21239 ;
  assign n7596 = n7594 | n7595 ;
  assign n21240 = ~n7596 ;
  assign n7597 = n7591 & n21240 ;
  assign n7598 = n7590 | n7597 ;
  assign n7599 = x73 & n7598 ;
  assign n7600 = x73 | n7598 ;
  assign n7601 = n7231 & n21088 ;
  assign n7602 = n152 & n7601 ;
  assign n21241 = ~n7237 ;
  assign n7603 = n21241 & n7602 ;
  assign n21242 = ~n7602 ;
  assign n7604 = n7237 & n21242 ;
  assign n7605 = n7603 | n7604 ;
  assign n21243 = ~n7605 ;
  assign n7606 = n7600 & n21243 ;
  assign n7607 = n7599 | n7606 ;
  assign n7608 = x74 & n7607 ;
  assign n7609 = x74 | n7607 ;
  assign n7610 = n7240 & n21092 ;
  assign n7611 = n152 & n7610 ;
  assign n21244 = ~n7246 ;
  assign n7612 = n21244 & n7611 ;
  assign n21245 = ~n7611 ;
  assign n7613 = n7246 & n21245 ;
  assign n7614 = n7612 | n7613 ;
  assign n21246 = ~n7614 ;
  assign n7615 = n7609 & n21246 ;
  assign n7616 = n7608 | n7615 ;
  assign n7617 = x75 & n7616 ;
  assign n7618 = x75 | n7616 ;
  assign n7619 = n7249 & n21096 ;
  assign n7620 = n152 & n7619 ;
  assign n21247 = ~n7255 ;
  assign n7621 = n21247 & n7620 ;
  assign n21248 = ~n7620 ;
  assign n7622 = n7255 & n21248 ;
  assign n7623 = n7621 | n7622 ;
  assign n21249 = ~n7623 ;
  assign n7624 = n7618 & n21249 ;
  assign n7625 = n7617 | n7624 ;
  assign n7626 = x76 & n7625 ;
  assign n7627 = x76 | n7625 ;
  assign n7628 = n7258 & n21100 ;
  assign n7629 = n152 & n7628 ;
  assign n7630 = n7264 & n7629 ;
  assign n7631 = n7264 | n7629 ;
  assign n21250 = ~n7630 ;
  assign n7632 = n21250 & n7631 ;
  assign n21251 = ~n7632 ;
  assign n7633 = n7627 & n21251 ;
  assign n7634 = n7626 | n7633 ;
  assign n7635 = x77 & n7634 ;
  assign n7636 = x77 | n7634 ;
  assign n7637 = n7267 & n21104 ;
  assign n7638 = n152 & n7637 ;
  assign n7639 = n7273 & n7638 ;
  assign n7640 = n7273 | n7638 ;
  assign n21252 = ~n7639 ;
  assign n7641 = n21252 & n7640 ;
  assign n21253 = ~n7641 ;
  assign n7642 = n7636 & n21253 ;
  assign n7643 = n7635 | n7642 ;
  assign n7644 = x78 & n7643 ;
  assign n7645 = x78 | n7643 ;
  assign n7646 = n7276 & n21108 ;
  assign n7647 = n152 & n7646 ;
  assign n21254 = ~n7282 ;
  assign n7648 = n21254 & n7647 ;
  assign n21255 = ~n7647 ;
  assign n7649 = n7282 & n21255 ;
  assign n7650 = n7648 | n7649 ;
  assign n21256 = ~n7650 ;
  assign n7651 = n7645 & n21256 ;
  assign n7652 = n7644 | n7651 ;
  assign n7653 = x79 & n7652 ;
  assign n7654 = x79 | n7652 ;
  assign n7655 = n7285 & n21112 ;
  assign n7656 = n152 & n7655 ;
  assign n21257 = ~n7291 ;
  assign n7657 = n21257 & n7656 ;
  assign n21258 = ~n7656 ;
  assign n7658 = n7291 & n21258 ;
  assign n7659 = n7657 | n7658 ;
  assign n21259 = ~n7659 ;
  assign n7660 = n7654 & n21259 ;
  assign n7661 = n7653 | n7660 ;
  assign n7662 = x80 & n7661 ;
  assign n7663 = x80 | n7661 ;
  assign n7664 = n7294 & n21116 ;
  assign n7665 = n152 & n7664 ;
  assign n21260 = ~n7300 ;
  assign n7666 = n21260 & n7665 ;
  assign n21261 = ~n7665 ;
  assign n7667 = n7300 & n21261 ;
  assign n7668 = n7666 | n7667 ;
  assign n21262 = ~n7668 ;
  assign n7669 = n7663 & n21262 ;
  assign n7670 = n7662 | n7669 ;
  assign n7671 = x81 & n7670 ;
  assign n7672 = x81 | n7670 ;
  assign n7673 = n7303 & n21120 ;
  assign n7674 = n152 & n7673 ;
  assign n21263 = ~n7309 ;
  assign n7675 = n21263 & n7674 ;
  assign n21264 = ~n7674 ;
  assign n7676 = n7309 & n21264 ;
  assign n7677 = n7675 | n7676 ;
  assign n21265 = ~n7677 ;
  assign n7678 = n7672 & n21265 ;
  assign n7679 = n7671 | n7678 ;
  assign n7680 = x82 & n7679 ;
  assign n7681 = x82 | n7679 ;
  assign n7682 = n7312 & n21124 ;
  assign n7683 = n152 & n7682 ;
  assign n7684 = n7318 & n7683 ;
  assign n7685 = n7318 | n7683 ;
  assign n21266 = ~n7684 ;
  assign n7686 = n21266 & n7685 ;
  assign n21267 = ~n7686 ;
  assign n7687 = n7681 & n21267 ;
  assign n7688 = n7680 | n7687 ;
  assign n7689 = x83 & n7688 ;
  assign n7690 = x83 | n7688 ;
  assign n7691 = n7321 & n21128 ;
  assign n7692 = n152 & n7691 ;
  assign n21268 = ~n7327 ;
  assign n7693 = n21268 & n7692 ;
  assign n21269 = ~n7692 ;
  assign n7694 = n7327 & n21269 ;
  assign n7695 = n7693 | n7694 ;
  assign n21270 = ~n7695 ;
  assign n7696 = n7690 & n21270 ;
  assign n7697 = n7689 | n7696 ;
  assign n7698 = x84 & n7697 ;
  assign n7699 = x84 | n7697 ;
  assign n7700 = n7330 & n21132 ;
  assign n7701 = n152 & n7700 ;
  assign n7702 = n7336 & n7701 ;
  assign n7703 = n7336 | n7701 ;
  assign n21271 = ~n7702 ;
  assign n7704 = n21271 & n7703 ;
  assign n21272 = ~n7704 ;
  assign n7705 = n7699 & n21272 ;
  assign n7706 = n7698 | n7705 ;
  assign n7707 = x85 & n7706 ;
  assign n7708 = x85 | n7706 ;
  assign n7709 = n7339 & n21136 ;
  assign n7710 = n152 & n7709 ;
  assign n21273 = ~n7345 ;
  assign n7711 = n21273 & n7710 ;
  assign n21274 = ~n7710 ;
  assign n7712 = n7345 & n21274 ;
  assign n7713 = n7711 | n7712 ;
  assign n21275 = ~n7713 ;
  assign n7714 = n7708 & n21275 ;
  assign n7715 = n7707 | n7714 ;
  assign n7716 = x86 & n7715 ;
  assign n7717 = x86 | n7715 ;
  assign n7718 = n7348 & n21140 ;
  assign n7719 = n152 & n7718 ;
  assign n21276 = ~n7354 ;
  assign n7720 = n21276 & n7719 ;
  assign n21277 = ~n7719 ;
  assign n7721 = n7354 & n21277 ;
  assign n7722 = n7720 | n7721 ;
  assign n21278 = ~n7722 ;
  assign n7723 = n7717 & n21278 ;
  assign n7724 = n7716 | n7723 ;
  assign n7725 = x87 & n7724 ;
  assign n7726 = x87 | n7724 ;
  assign n7727 = n7357 & n21144 ;
  assign n7728 = n152 & n7727 ;
  assign n21279 = ~n7363 ;
  assign n7729 = n21279 & n7728 ;
  assign n21280 = ~n7728 ;
  assign n7730 = n7363 & n21280 ;
  assign n7731 = n7729 | n7730 ;
  assign n21281 = ~n7731 ;
  assign n7732 = n7726 & n21281 ;
  assign n7733 = n7725 | n7732 ;
  assign n7734 = x88 & n7733 ;
  assign n7735 = x88 | n7733 ;
  assign n7736 = n7366 & n21148 ;
  assign n7737 = n152 & n7736 ;
  assign n21282 = ~n7372 ;
  assign n7738 = n21282 & n7737 ;
  assign n21283 = ~n7737 ;
  assign n7739 = n7372 & n21283 ;
  assign n7740 = n7738 | n7739 ;
  assign n21284 = ~n7740 ;
  assign n7741 = n7735 & n21284 ;
  assign n7742 = n7734 | n7741 ;
  assign n7743 = x89 & n7742 ;
  assign n7744 = x89 | n7742 ;
  assign n7745 = n7375 & n21152 ;
  assign n7746 = n152 & n7745 ;
  assign n21285 = ~n7381 ;
  assign n7747 = n21285 & n7746 ;
  assign n21286 = ~n7746 ;
  assign n7748 = n7381 & n21286 ;
  assign n7749 = n7747 | n7748 ;
  assign n21287 = ~n7749 ;
  assign n7750 = n7744 & n21287 ;
  assign n7751 = n7743 | n7750 ;
  assign n7752 = x90 & n7751 ;
  assign n7753 = x90 | n7751 ;
  assign n7754 = n7384 & n21156 ;
  assign n7755 = n152 & n7754 ;
  assign n7756 = n7390 & n7755 ;
  assign n7757 = n7390 | n7755 ;
  assign n21288 = ~n7756 ;
  assign n7758 = n21288 & n7757 ;
  assign n21289 = ~n7758 ;
  assign n7759 = n7753 & n21289 ;
  assign n7760 = n7752 | n7759 ;
  assign n7761 = x91 & n7760 ;
  assign n7762 = x91 | n7760 ;
  assign n7763 = n7393 & n21160 ;
  assign n7764 = n152 & n7763 ;
  assign n21290 = ~n7399 ;
  assign n7765 = n21290 & n7764 ;
  assign n21291 = ~n7764 ;
  assign n7766 = n7399 & n21291 ;
  assign n7767 = n7765 | n7766 ;
  assign n21292 = ~n7767 ;
  assign n7768 = n7762 & n21292 ;
  assign n7769 = n7761 | n7768 ;
  assign n7770 = x92 & n7769 ;
  assign n7771 = x92 | n7769 ;
  assign n7772 = n7402 & n21164 ;
  assign n7773 = n152 & n7772 ;
  assign n21293 = ~n7408 ;
  assign n7774 = n21293 & n7773 ;
  assign n21294 = ~n7773 ;
  assign n7775 = n7408 & n21294 ;
  assign n7776 = n7774 | n7775 ;
  assign n21295 = ~n7776 ;
  assign n7777 = n7771 & n21295 ;
  assign n7778 = n7770 | n7777 ;
  assign n7779 = x93 & n7778 ;
  assign n7780 = x93 | n7778 ;
  assign n7781 = n7411 & n21168 ;
  assign n7782 = n152 & n7781 ;
  assign n7783 = n7417 & n7782 ;
  assign n7784 = n7417 | n7782 ;
  assign n21296 = ~n7783 ;
  assign n7785 = n21296 & n7784 ;
  assign n21297 = ~n7785 ;
  assign n7786 = n7780 & n21297 ;
  assign n7787 = n7779 | n7786 ;
  assign n7788 = x94 & n7787 ;
  assign n7789 = x94 | n7787 ;
  assign n7790 = n7420 & n21172 ;
  assign n7791 = n152 & n7790 ;
  assign n7792 = n7426 & n7791 ;
  assign n7793 = n7426 | n7791 ;
  assign n21298 = ~n7792 ;
  assign n7794 = n21298 & n7793 ;
  assign n21299 = ~n7794 ;
  assign n7795 = n7789 & n21299 ;
  assign n7796 = n7788 | n7795 ;
  assign n7797 = x95 & n7796 ;
  assign n7798 = x95 | n7796 ;
  assign n7799 = n7429 & n21176 ;
  assign n7800 = n152 & n7799 ;
  assign n21300 = ~n7435 ;
  assign n7801 = n21300 & n7800 ;
  assign n21301 = ~n7800 ;
  assign n7802 = n7435 & n21301 ;
  assign n7803 = n7801 | n7802 ;
  assign n21302 = ~n7803 ;
  assign n7804 = n7798 & n21302 ;
  assign n7805 = n7797 | n7804 ;
  assign n7806 = x96 & n7805 ;
  assign n7807 = x96 | n7805 ;
  assign n7808 = n7438 & n21180 ;
  assign n7809 = n152 & n7808 ;
  assign n7810 = n7444 & n7809 ;
  assign n7811 = n7444 | n7809 ;
  assign n21303 = ~n7810 ;
  assign n7812 = n21303 & n7811 ;
  assign n21304 = ~n7812 ;
  assign n7813 = n7807 & n21304 ;
  assign n7814 = n7806 | n7813 ;
  assign n7815 = x97 & n7814 ;
  assign n7816 = x97 | n7814 ;
  assign n7817 = n7447 & n21184 ;
  assign n7818 = n152 & n7817 ;
  assign n21305 = ~n7453 ;
  assign n7819 = n21305 & n7818 ;
  assign n21306 = ~n7818 ;
  assign n7820 = n7453 & n21306 ;
  assign n7821 = n7819 | n7820 ;
  assign n21307 = ~n7821 ;
  assign n7822 = n7816 & n21307 ;
  assign n7823 = n7815 | n7822 ;
  assign n7824 = x98 & n7823 ;
  assign n7825 = x98 | n7823 ;
  assign n7826 = n7456 & n21188 ;
  assign n7827 = n152 & n7826 ;
  assign n21308 = ~n7462 ;
  assign n7828 = n21308 & n7827 ;
  assign n21309 = ~n7827 ;
  assign n7829 = n7462 & n21309 ;
  assign n7830 = n7828 | n7829 ;
  assign n21310 = ~n7830 ;
  assign n7831 = n7825 & n21310 ;
  assign n7832 = n7824 | n7831 ;
  assign n7833 = x99 & n7832 ;
  assign n7834 = x99 | n7832 ;
  assign n7835 = n7465 & n21192 ;
  assign n7836 = n152 & n7835 ;
  assign n7837 = n7471 & n7836 ;
  assign n7838 = n7471 | n7836 ;
  assign n21311 = ~n7837 ;
  assign n7839 = n21311 & n7838 ;
  assign n21312 = ~n7839 ;
  assign n7840 = n7834 & n21312 ;
  assign n7841 = n7833 | n7840 ;
  assign n7842 = x100 & n7841 ;
  assign n7843 = x100 | n7841 ;
  assign n7844 = n7474 & n21196 ;
  assign n7845 = n152 & n7844 ;
  assign n7846 = n7480 & n7845 ;
  assign n7847 = n7480 | n7845 ;
  assign n21313 = ~n7846 ;
  assign n7848 = n21313 & n7847 ;
  assign n21314 = ~n7848 ;
  assign n7849 = n7843 & n21314 ;
  assign n7850 = n7842 | n7849 ;
  assign n7851 = x101 & n7850 ;
  assign n7852 = x101 | n7850 ;
  assign n7853 = n7483 & n21200 ;
  assign n7854 = n152 & n7853 ;
  assign n7855 = n7489 & n7854 ;
  assign n7856 = n7489 | n7854 ;
  assign n21315 = ~n7855 ;
  assign n7857 = n21315 & n7856 ;
  assign n21316 = ~n7857 ;
  assign n7858 = n7852 & n21316 ;
  assign n7859 = n7851 | n7858 ;
  assign n7860 = x102 & n7859 ;
  assign n7861 = x102 | n7859 ;
  assign n7862 = n7492 & n21204 ;
  assign n7863 = n152 & n7862 ;
  assign n7864 = n7498 & n7863 ;
  assign n7865 = n7498 | n7863 ;
  assign n21317 = ~n7864 ;
  assign n7866 = n21317 & n7865 ;
  assign n21318 = ~n7866 ;
  assign n7867 = n7861 & n21318 ;
  assign n7868 = n7860 | n7867 ;
  assign n7869 = x103 & n7868 ;
  assign n7870 = x103 | n7868 ;
  assign n7871 = n7501 & n21208 ;
  assign n7872 = n152 & n7871 ;
  assign n7873 = n7507 & n7872 ;
  assign n7874 = n7507 | n7872 ;
  assign n21319 = ~n7873 ;
  assign n7875 = n21319 & n7874 ;
  assign n21320 = ~n7875 ;
  assign n7876 = n7870 & n21320 ;
  assign n7877 = n7869 | n7876 ;
  assign n7879 = x104 & n7877 ;
  assign n7878 = x104 | n7877 ;
  assign n21321 = ~n7879 ;
  assign n7880 = n7526 & n21321 ;
  assign n7518 = n21884 | n7517 ;
  assign n7881 = n7167 & n7518 ;
  assign n21322 = ~x105 ;
  assign n7882 = n21322 & n7881 ;
  assign n21323 = ~n7882 ;
  assign n7883 = n7878 & n21323 ;
  assign n21324 = ~n7880 ;
  assign n7884 = n21324 & n7883 ;
  assign n7885 = n18368 | n7884 ;
  assign n21325 = ~n7881 ;
  assign n7887 = x105 & n21325 ;
  assign n7888 = n7885 | n7887 ;
  assign n151 = ~n7888 ;
  assign n7889 = n7878 & n151 ;
  assign n7890 = n21321 & n7889 ;
  assign n7891 = n7526 | n7890 ;
  assign n7892 = n7880 & n7889 ;
  assign n21327 = ~n7892 ;
  assign n7893 = n7891 & n21327 ;
  assign n21328 = ~x21 ;
  assign n7894 = n21328 & x64 ;
  assign n7896 = x65 | n7894 ;
  assign n7895 = x65 & n7894 ;
  assign n7897 = x64 & n151 ;
  assign n7898 = x22 & n7897 ;
  assign n7899 = x22 | n7897 ;
  assign n21329 = ~n7898 ;
  assign n7900 = n21329 & n7899 ;
  assign n21330 = ~n7895 ;
  assign n7901 = n21330 & n7900 ;
  assign n21331 = ~n7901 ;
  assign n7902 = n7896 & n21331 ;
  assign n7903 = x66 & n7902 ;
  assign n7904 = x66 | n7902 ;
  assign n7905 = n21222 & n7529 ;
  assign n7906 = n151 & n7905 ;
  assign n7907 = n7533 & n7906 ;
  assign n7908 = n7533 | n7906 ;
  assign n21332 = ~n7907 ;
  assign n7909 = n21332 & n7908 ;
  assign n21333 = ~n7909 ;
  assign n7910 = n7904 & n21333 ;
  assign n7911 = n7903 | n7910 ;
  assign n7912 = x67 & n7911 ;
  assign n7913 = x67 | n7911 ;
  assign n21334 = ~n7536 ;
  assign n7914 = n21334 & n7537 ;
  assign n7915 = n151 & n7914 ;
  assign n7916 = n7542 & n7915 ;
  assign n7917 = n7542 | n7915 ;
  assign n21335 = ~n7916 ;
  assign n7918 = n21335 & n7917 ;
  assign n21336 = ~n7918 ;
  assign n7919 = n7913 & n21336 ;
  assign n7920 = n7912 | n7919 ;
  assign n7921 = x68 & n7920 ;
  assign n7922 = x68 | n7920 ;
  assign n21337 = ~n7545 ;
  assign n7923 = n21337 & n7546 ;
  assign n7924 = n151 & n7923 ;
  assign n7925 = n7551 & n7924 ;
  assign n7926 = n7551 | n7924 ;
  assign n21338 = ~n7925 ;
  assign n7927 = n21338 & n7926 ;
  assign n21339 = ~n7927 ;
  assign n7928 = n7922 & n21339 ;
  assign n7929 = n7921 | n7928 ;
  assign n7930 = x69 & n7929 ;
  assign n7931 = x69 | n7929 ;
  assign n21340 = ~n7554 ;
  assign n7932 = n21340 & n7555 ;
  assign n7933 = n151 & n7932 ;
  assign n7934 = n7560 & n7933 ;
  assign n7935 = n7560 | n7933 ;
  assign n21341 = ~n7934 ;
  assign n7936 = n21341 & n7935 ;
  assign n21342 = ~n7936 ;
  assign n7937 = n7931 & n21342 ;
  assign n7938 = n7930 | n7937 ;
  assign n7939 = x70 & n7938 ;
  assign n7940 = x70 | n7938 ;
  assign n21343 = ~n7563 ;
  assign n7941 = n21343 & n7564 ;
  assign n7942 = n151 & n7941 ;
  assign n7943 = n21233 & n7942 ;
  assign n21344 = ~n7942 ;
  assign n7944 = n7569 & n21344 ;
  assign n7945 = n7943 | n7944 ;
  assign n21345 = ~n7945 ;
  assign n7946 = n7940 & n21345 ;
  assign n7947 = n7939 | n7946 ;
  assign n7948 = x71 & n7947 ;
  assign n7949 = x71 | n7947 ;
  assign n21346 = ~n7572 ;
  assign n7950 = n21346 & n7573 ;
  assign n7951 = n151 & n7950 ;
  assign n7952 = n7578 & n7951 ;
  assign n7953 = n7578 | n7951 ;
  assign n21347 = ~n7952 ;
  assign n7954 = n21347 & n7953 ;
  assign n21348 = ~n7954 ;
  assign n7955 = n7949 & n21348 ;
  assign n7956 = n7948 | n7955 ;
  assign n7957 = x72 & n7956 ;
  assign n7958 = x72 | n7956 ;
  assign n21349 = ~n7581 ;
  assign n7959 = n21349 & n7582 ;
  assign n7960 = n151 & n7959 ;
  assign n7961 = n7587 & n7960 ;
  assign n7962 = n7587 | n7960 ;
  assign n21350 = ~n7961 ;
  assign n7963 = n21350 & n7962 ;
  assign n21351 = ~n7963 ;
  assign n7964 = n7958 & n21351 ;
  assign n7965 = n7957 | n7964 ;
  assign n7966 = x73 & n7965 ;
  assign n7967 = x73 | n7965 ;
  assign n21352 = ~n7590 ;
  assign n7968 = n21352 & n7591 ;
  assign n7969 = n151 & n7968 ;
  assign n7970 = n21240 & n7969 ;
  assign n21353 = ~n7969 ;
  assign n7971 = n7596 & n21353 ;
  assign n7972 = n7970 | n7971 ;
  assign n21354 = ~n7972 ;
  assign n7973 = n7967 & n21354 ;
  assign n7974 = n7966 | n7973 ;
  assign n7975 = x74 & n7974 ;
  assign n7976 = x74 | n7974 ;
  assign n21355 = ~n7599 ;
  assign n7977 = n21355 & n7600 ;
  assign n7978 = n151 & n7977 ;
  assign n7979 = n21243 & n7978 ;
  assign n21356 = ~n7978 ;
  assign n7980 = n7605 & n21356 ;
  assign n7981 = n7979 | n7980 ;
  assign n21357 = ~n7981 ;
  assign n7982 = n7976 & n21357 ;
  assign n7983 = n7975 | n7982 ;
  assign n7984 = x75 & n7983 ;
  assign n7985 = x75 | n7983 ;
  assign n21358 = ~n7608 ;
  assign n7986 = n21358 & n7609 ;
  assign n7987 = n151 & n7986 ;
  assign n7988 = n7614 & n7987 ;
  assign n7989 = n7614 | n7987 ;
  assign n21359 = ~n7988 ;
  assign n7990 = n21359 & n7989 ;
  assign n21360 = ~n7990 ;
  assign n7991 = n7985 & n21360 ;
  assign n7992 = n7984 | n7991 ;
  assign n7993 = x76 & n7992 ;
  assign n7994 = x76 | n7992 ;
  assign n21361 = ~n7617 ;
  assign n7995 = n21361 & n7618 ;
  assign n7996 = n151 & n7995 ;
  assign n7997 = n21249 & n7996 ;
  assign n21362 = ~n7996 ;
  assign n7998 = n7623 & n21362 ;
  assign n7999 = n7997 | n7998 ;
  assign n21363 = ~n7999 ;
  assign n8000 = n7994 & n21363 ;
  assign n8001 = n7993 | n8000 ;
  assign n8002 = x77 & n8001 ;
  assign n8003 = x77 | n8001 ;
  assign n21364 = ~n7626 ;
  assign n8004 = n21364 & n7627 ;
  assign n8005 = n151 & n8004 ;
  assign n8006 = n7632 & n8005 ;
  assign n8007 = n7632 | n8005 ;
  assign n21365 = ~n8006 ;
  assign n8008 = n21365 & n8007 ;
  assign n21366 = ~n8008 ;
  assign n8009 = n8003 & n21366 ;
  assign n8010 = n8002 | n8009 ;
  assign n8011 = x78 & n8010 ;
  assign n8012 = x78 | n8010 ;
  assign n21367 = ~n7635 ;
  assign n8013 = n21367 & n7636 ;
  assign n8014 = n151 & n8013 ;
  assign n8015 = n7641 & n8014 ;
  assign n8016 = n7641 | n8014 ;
  assign n21368 = ~n8015 ;
  assign n8017 = n21368 & n8016 ;
  assign n21369 = ~n8017 ;
  assign n8018 = n8012 & n21369 ;
  assign n8019 = n8011 | n8018 ;
  assign n8020 = x79 & n8019 ;
  assign n8021 = x79 | n8019 ;
  assign n21370 = ~n7644 ;
  assign n8022 = n21370 & n7645 ;
  assign n8023 = n151 & n8022 ;
  assign n8024 = n21256 & n8023 ;
  assign n21371 = ~n8023 ;
  assign n8025 = n7650 & n21371 ;
  assign n8026 = n8024 | n8025 ;
  assign n21372 = ~n8026 ;
  assign n8027 = n8021 & n21372 ;
  assign n8028 = n8020 | n8027 ;
  assign n8029 = x80 & n8028 ;
  assign n8030 = x80 | n8028 ;
  assign n21373 = ~n7653 ;
  assign n8031 = n21373 & n7654 ;
  assign n8032 = n151 & n8031 ;
  assign n8033 = n21259 & n8032 ;
  assign n21374 = ~n8032 ;
  assign n8034 = n7659 & n21374 ;
  assign n8035 = n8033 | n8034 ;
  assign n21375 = ~n8035 ;
  assign n8036 = n8030 & n21375 ;
  assign n8037 = n8029 | n8036 ;
  assign n8038 = x81 & n8037 ;
  assign n8039 = x81 | n8037 ;
  assign n21376 = ~n7662 ;
  assign n8040 = n21376 & n7663 ;
  assign n8041 = n151 & n8040 ;
  assign n8042 = n21262 & n8041 ;
  assign n21377 = ~n8041 ;
  assign n8043 = n7668 & n21377 ;
  assign n8044 = n8042 | n8043 ;
  assign n21378 = ~n8044 ;
  assign n8045 = n8039 & n21378 ;
  assign n8046 = n8038 | n8045 ;
  assign n8047 = x82 & n8046 ;
  assign n8048 = x82 | n8046 ;
  assign n21379 = ~n7671 ;
  assign n8049 = n21379 & n7672 ;
  assign n8050 = n151 & n8049 ;
  assign n8051 = n21265 & n8050 ;
  assign n21380 = ~n8050 ;
  assign n8052 = n7677 & n21380 ;
  assign n8053 = n8051 | n8052 ;
  assign n21381 = ~n8053 ;
  assign n8054 = n8048 & n21381 ;
  assign n8055 = n8047 | n8054 ;
  assign n8056 = x83 & n8055 ;
  assign n8057 = x83 | n8055 ;
  assign n21382 = ~n7680 ;
  assign n8058 = n21382 & n7681 ;
  assign n8059 = n151 & n8058 ;
  assign n8060 = n7686 & n8059 ;
  assign n8061 = n7686 | n8059 ;
  assign n21383 = ~n8060 ;
  assign n8062 = n21383 & n8061 ;
  assign n21384 = ~n8062 ;
  assign n8063 = n8057 & n21384 ;
  assign n8064 = n8056 | n8063 ;
  assign n8065 = x84 & n8064 ;
  assign n8066 = x84 | n8064 ;
  assign n21385 = ~n7689 ;
  assign n8067 = n21385 & n7690 ;
  assign n8068 = n151 & n8067 ;
  assign n8069 = n7695 & n8068 ;
  assign n8070 = n7695 | n8068 ;
  assign n21386 = ~n8069 ;
  assign n8071 = n21386 & n8070 ;
  assign n21387 = ~n8071 ;
  assign n8072 = n8066 & n21387 ;
  assign n8073 = n8065 | n8072 ;
  assign n8074 = x85 & n8073 ;
  assign n8075 = x85 | n8073 ;
  assign n21388 = ~n7698 ;
  assign n8076 = n21388 & n7699 ;
  assign n8077 = n151 & n8076 ;
  assign n8078 = n7704 & n8077 ;
  assign n8079 = n7704 | n8077 ;
  assign n21389 = ~n8078 ;
  assign n8080 = n21389 & n8079 ;
  assign n21390 = ~n8080 ;
  assign n8081 = n8075 & n21390 ;
  assign n8082 = n8074 | n8081 ;
  assign n8083 = x86 & n8082 ;
  assign n8084 = x86 | n8082 ;
  assign n21391 = ~n7707 ;
  assign n8085 = n21391 & n7708 ;
  assign n8086 = n151 & n8085 ;
  assign n8087 = n21275 & n8086 ;
  assign n21392 = ~n8086 ;
  assign n8088 = n7713 & n21392 ;
  assign n8089 = n8087 | n8088 ;
  assign n21393 = ~n8089 ;
  assign n8090 = n8084 & n21393 ;
  assign n8091 = n8083 | n8090 ;
  assign n8092 = x87 & n8091 ;
  assign n8093 = x87 | n8091 ;
  assign n21394 = ~n7716 ;
  assign n8094 = n21394 & n7717 ;
  assign n8095 = n151 & n8094 ;
  assign n8096 = n21278 & n8095 ;
  assign n21395 = ~n8095 ;
  assign n8097 = n7722 & n21395 ;
  assign n8098 = n8096 | n8097 ;
  assign n21396 = ~n8098 ;
  assign n8099 = n8093 & n21396 ;
  assign n8100 = n8092 | n8099 ;
  assign n8101 = x88 & n8100 ;
  assign n8102 = x88 | n8100 ;
  assign n21397 = ~n7725 ;
  assign n8103 = n21397 & n7726 ;
  assign n8104 = n151 & n8103 ;
  assign n8105 = n21281 & n8104 ;
  assign n21398 = ~n8104 ;
  assign n8106 = n7731 & n21398 ;
  assign n8107 = n8105 | n8106 ;
  assign n21399 = ~n8107 ;
  assign n8108 = n8102 & n21399 ;
  assign n8109 = n8101 | n8108 ;
  assign n8110 = x89 & n8109 ;
  assign n8111 = x89 | n8109 ;
  assign n21400 = ~n7734 ;
  assign n8112 = n21400 & n7735 ;
  assign n8113 = n151 & n8112 ;
  assign n8114 = n7740 & n8113 ;
  assign n8115 = n7740 | n8113 ;
  assign n21401 = ~n8114 ;
  assign n8116 = n21401 & n8115 ;
  assign n21402 = ~n8116 ;
  assign n8117 = n8111 & n21402 ;
  assign n8118 = n8110 | n8117 ;
  assign n8119 = x90 & n8118 ;
  assign n8120 = x90 | n8118 ;
  assign n21403 = ~n7743 ;
  assign n8121 = n21403 & n7744 ;
  assign n8122 = n151 & n8121 ;
  assign n8123 = n7749 & n8122 ;
  assign n8124 = n7749 | n8122 ;
  assign n21404 = ~n8123 ;
  assign n8125 = n21404 & n8124 ;
  assign n21405 = ~n8125 ;
  assign n8126 = n8120 & n21405 ;
  assign n8127 = n8119 | n8126 ;
  assign n8128 = x91 & n8127 ;
  assign n8129 = x91 | n8127 ;
  assign n21406 = ~n7752 ;
  assign n8130 = n21406 & n7753 ;
  assign n8131 = n151 & n8130 ;
  assign n8132 = n7758 & n8131 ;
  assign n8133 = n7758 | n8131 ;
  assign n21407 = ~n8132 ;
  assign n8134 = n21407 & n8133 ;
  assign n21408 = ~n8134 ;
  assign n8135 = n8129 & n21408 ;
  assign n8136 = n8128 | n8135 ;
  assign n8137 = x92 & n8136 ;
  assign n8138 = x92 | n8136 ;
  assign n21409 = ~n7761 ;
  assign n8139 = n21409 & n7762 ;
  assign n8140 = n151 & n8139 ;
  assign n8141 = n21292 & n8140 ;
  assign n21410 = ~n8140 ;
  assign n8142 = n7767 & n21410 ;
  assign n8143 = n8141 | n8142 ;
  assign n21411 = ~n8143 ;
  assign n8144 = n8138 & n21411 ;
  assign n8145 = n8137 | n8144 ;
  assign n8146 = x93 & n8145 ;
  assign n8147 = x93 | n8145 ;
  assign n21412 = ~n7770 ;
  assign n8148 = n21412 & n7771 ;
  assign n8149 = n151 & n8148 ;
  assign n8150 = n21295 & n8149 ;
  assign n21413 = ~n8149 ;
  assign n8151 = n7776 & n21413 ;
  assign n8152 = n8150 | n8151 ;
  assign n21414 = ~n8152 ;
  assign n8153 = n8147 & n21414 ;
  assign n8154 = n8146 | n8153 ;
  assign n8155 = x94 & n8154 ;
  assign n8156 = x94 | n8154 ;
  assign n21415 = ~n7779 ;
  assign n8157 = n21415 & n7780 ;
  assign n8158 = n151 & n8157 ;
  assign n8159 = n7785 & n8158 ;
  assign n8160 = n7785 | n8158 ;
  assign n21416 = ~n8159 ;
  assign n8161 = n21416 & n8160 ;
  assign n21417 = ~n8161 ;
  assign n8162 = n8156 & n21417 ;
  assign n8163 = n8155 | n8162 ;
  assign n8164 = x95 & n8163 ;
  assign n8165 = x95 | n8163 ;
  assign n21418 = ~n7788 ;
  assign n8166 = n21418 & n7789 ;
  assign n8167 = n151 & n8166 ;
  assign n8168 = n7794 & n8167 ;
  assign n8169 = n7794 | n8167 ;
  assign n21419 = ~n8168 ;
  assign n8170 = n21419 & n8169 ;
  assign n21420 = ~n8170 ;
  assign n8171 = n8165 & n21420 ;
  assign n8172 = n8164 | n8171 ;
  assign n8173 = x96 & n8172 ;
  assign n8174 = x96 | n8172 ;
  assign n21421 = ~n7797 ;
  assign n8175 = n21421 & n7798 ;
  assign n8176 = n151 & n8175 ;
  assign n8177 = n21302 & n8176 ;
  assign n21422 = ~n8176 ;
  assign n8178 = n7803 & n21422 ;
  assign n8179 = n8177 | n8178 ;
  assign n21423 = ~n8179 ;
  assign n8180 = n8174 & n21423 ;
  assign n8181 = n8173 | n8180 ;
  assign n8182 = x97 & n8181 ;
  assign n8183 = x97 | n8181 ;
  assign n21424 = ~n7806 ;
  assign n8184 = n21424 & n7807 ;
  assign n8185 = n151 & n8184 ;
  assign n8186 = n7812 & n8185 ;
  assign n8187 = n7812 | n8185 ;
  assign n21425 = ~n8186 ;
  assign n8188 = n21425 & n8187 ;
  assign n21426 = ~n8188 ;
  assign n8189 = n8183 & n21426 ;
  assign n8190 = n8182 | n8189 ;
  assign n8191 = x98 & n8190 ;
  assign n8192 = x98 | n8190 ;
  assign n21427 = ~n7815 ;
  assign n8193 = n21427 & n7816 ;
  assign n8194 = n151 & n8193 ;
  assign n8195 = n21307 & n8194 ;
  assign n21428 = ~n8194 ;
  assign n8196 = n7821 & n21428 ;
  assign n8197 = n8195 | n8196 ;
  assign n21429 = ~n8197 ;
  assign n8198 = n8192 & n21429 ;
  assign n8199 = n8191 | n8198 ;
  assign n8200 = x99 & n8199 ;
  assign n8201 = x99 | n8199 ;
  assign n21430 = ~n7824 ;
  assign n8202 = n21430 & n7825 ;
  assign n8203 = n151 & n8202 ;
  assign n8204 = n21310 & n8203 ;
  assign n21431 = ~n8203 ;
  assign n8205 = n7830 & n21431 ;
  assign n8206 = n8204 | n8205 ;
  assign n21432 = ~n8206 ;
  assign n8207 = n8201 & n21432 ;
  assign n8208 = n8200 | n8207 ;
  assign n8209 = x100 & n8208 ;
  assign n8210 = x100 | n8208 ;
  assign n21433 = ~n7833 ;
  assign n8211 = n21433 & n7834 ;
  assign n8212 = n151 & n8211 ;
  assign n8213 = n7839 & n8212 ;
  assign n8214 = n7839 | n8212 ;
  assign n21434 = ~n8213 ;
  assign n8215 = n21434 & n8214 ;
  assign n21435 = ~n8215 ;
  assign n8216 = n8210 & n21435 ;
  assign n8217 = n8209 | n8216 ;
  assign n8218 = x101 & n8217 ;
  assign n8219 = x101 | n8217 ;
  assign n21436 = ~n7842 ;
  assign n8220 = n21436 & n7843 ;
  assign n8221 = n151 & n8220 ;
  assign n8222 = n7848 & n8221 ;
  assign n8223 = n7848 | n8221 ;
  assign n21437 = ~n8222 ;
  assign n8224 = n21437 & n8223 ;
  assign n21438 = ~n8224 ;
  assign n8225 = n8219 & n21438 ;
  assign n8226 = n8218 | n8225 ;
  assign n8227 = x102 & n8226 ;
  assign n8228 = x102 | n8226 ;
  assign n21439 = ~n7851 ;
  assign n8229 = n21439 & n7852 ;
  assign n8230 = n151 & n8229 ;
  assign n8231 = n7857 & n8230 ;
  assign n8232 = n7857 | n8230 ;
  assign n21440 = ~n8231 ;
  assign n8233 = n21440 & n8232 ;
  assign n21441 = ~n8233 ;
  assign n8234 = n8228 & n21441 ;
  assign n8235 = n8227 | n8234 ;
  assign n8236 = x103 & n8235 ;
  assign n8237 = x103 | n8235 ;
  assign n21442 = ~n7860 ;
  assign n8238 = n21442 & n7861 ;
  assign n8239 = n151 & n8238 ;
  assign n8240 = n7866 & n8239 ;
  assign n8241 = n7866 | n8239 ;
  assign n21443 = ~n8240 ;
  assign n8242 = n21443 & n8241 ;
  assign n21444 = ~n8242 ;
  assign n8243 = n8237 & n21444 ;
  assign n8244 = n8236 | n8243 ;
  assign n8245 = x104 & n8244 ;
  assign n8246 = x104 | n8244 ;
  assign n21445 = ~n7869 ;
  assign n8247 = n21445 & n7870 ;
  assign n8248 = n151 & n8247 ;
  assign n8249 = n21320 & n8248 ;
  assign n21446 = ~n8248 ;
  assign n8250 = n7875 & n21446 ;
  assign n8251 = n8249 | n8250 ;
  assign n21447 = ~n8251 ;
  assign n8252 = n8246 & n21447 ;
  assign n8253 = n8245 | n8252 ;
  assign n8254 = x105 & n8253 ;
  assign n8255 = x105 | n8253 ;
  assign n21448 = ~n7893 ;
  assign n8256 = n21448 & n8255 ;
  assign n8257 = n8254 | n8256 ;
  assign n7886 = n21884 | n7885 ;
  assign n8259 = n7881 & n7886 ;
  assign n21449 = ~x106 ;
  assign n8261 = n21449 & n8259 ;
  assign n21450 = ~n8261 ;
  assign n8262 = n8257 & n21450 ;
  assign n21451 = ~n18363 ;
  assign n8263 = n21451 & n8259 ;
  assign n21452 = ~n8263 ;
  assign n8264 = n18368 & n21452 ;
  assign n8265 = n8262 | n8264 ;
  assign n21453 = ~n8254 ;
  assign n8266 = n21453 & n8255 ;
  assign n150 = ~n8265 ;
  assign n8267 = n150 & n8266 ;
  assign n8268 = n7893 & n8267 ;
  assign n8269 = n7893 | n8267 ;
  assign n21455 = ~n8268 ;
  assign n8270 = n21455 & n8269 ;
  assign n8258 = n18368 & n8257 ;
  assign n8271 = n21884 | n8258 ;
  assign n8272 = n8263 & n8271 ;
  assign n21456 = ~x20 ;
  assign n8273 = n21456 & x64 ;
  assign n8275 = x65 | n8273 ;
  assign n8274 = x65 & n8273 ;
  assign n8276 = x64 & n150 ;
  assign n8277 = x21 & n8276 ;
  assign n8278 = x21 | n8276 ;
  assign n21457 = ~n8277 ;
  assign n8279 = n21457 & n8278 ;
  assign n21458 = ~n8274 ;
  assign n8280 = n21458 & n8279 ;
  assign n21459 = ~n8280 ;
  assign n8281 = n8275 & n21459 ;
  assign n8282 = x66 & n8281 ;
  assign n8283 = x66 | n8281 ;
  assign n8284 = n21330 & n7896 ;
  assign n8285 = n150 & n8284 ;
  assign n8286 = n7900 & n8285 ;
  assign n8287 = n7900 | n8285 ;
  assign n21460 = ~n8286 ;
  assign n8288 = n21460 & n8287 ;
  assign n21461 = ~n8288 ;
  assign n8289 = n8283 & n21461 ;
  assign n8290 = n8282 | n8289 ;
  assign n8291 = x67 & n8290 ;
  assign n8292 = x67 | n8290 ;
  assign n21462 = ~n7903 ;
  assign n8293 = n21462 & n7904 ;
  assign n8294 = n150 & n8293 ;
  assign n8295 = n7909 & n8294 ;
  assign n8296 = n7909 | n8294 ;
  assign n21463 = ~n8295 ;
  assign n8297 = n21463 & n8296 ;
  assign n21464 = ~n8297 ;
  assign n8298 = n8292 & n21464 ;
  assign n8299 = n8291 | n8298 ;
  assign n8300 = x68 & n8299 ;
  assign n8301 = x68 | n8299 ;
  assign n21465 = ~n7912 ;
  assign n8302 = n21465 & n7913 ;
  assign n8303 = n150 & n8302 ;
  assign n8304 = n7918 & n8303 ;
  assign n8305 = n7918 | n8303 ;
  assign n21466 = ~n8304 ;
  assign n8306 = n21466 & n8305 ;
  assign n21467 = ~n8306 ;
  assign n8307 = n8301 & n21467 ;
  assign n8308 = n8300 | n8307 ;
  assign n8309 = x69 & n8308 ;
  assign n8310 = x69 | n8308 ;
  assign n21468 = ~n7921 ;
  assign n8311 = n21468 & n7922 ;
  assign n8312 = n150 & n8311 ;
  assign n8313 = n21339 & n8312 ;
  assign n21469 = ~n8312 ;
  assign n8314 = n7927 & n21469 ;
  assign n8315 = n8313 | n8314 ;
  assign n21470 = ~n8315 ;
  assign n8316 = n8310 & n21470 ;
  assign n8317 = n8309 | n8316 ;
  assign n8318 = x70 & n8317 ;
  assign n8319 = x70 | n8317 ;
  assign n21471 = ~n7930 ;
  assign n8320 = n21471 & n7931 ;
  assign n8321 = n150 & n8320 ;
  assign n8322 = n7936 & n8321 ;
  assign n8323 = n7936 | n8321 ;
  assign n21472 = ~n8322 ;
  assign n8324 = n21472 & n8323 ;
  assign n21473 = ~n8324 ;
  assign n8325 = n8319 & n21473 ;
  assign n8326 = n8318 | n8325 ;
  assign n8327 = x71 & n8326 ;
  assign n8328 = x71 | n8326 ;
  assign n21474 = ~n7939 ;
  assign n8329 = n21474 & n7940 ;
  assign n8330 = n150 & n8329 ;
  assign n8331 = n21345 & n8330 ;
  assign n21475 = ~n8330 ;
  assign n8332 = n7945 & n21475 ;
  assign n8333 = n8331 | n8332 ;
  assign n21476 = ~n8333 ;
  assign n8334 = n8328 & n21476 ;
  assign n8335 = n8327 | n8334 ;
  assign n8336 = x72 & n8335 ;
  assign n8337 = x72 | n8335 ;
  assign n21477 = ~n7948 ;
  assign n8338 = n21477 & n7949 ;
  assign n8339 = n150 & n8338 ;
  assign n8340 = n7954 & n8339 ;
  assign n8341 = n7954 | n8339 ;
  assign n21478 = ~n8340 ;
  assign n8342 = n21478 & n8341 ;
  assign n21479 = ~n8342 ;
  assign n8343 = n8337 & n21479 ;
  assign n8344 = n8336 | n8343 ;
  assign n8345 = x73 & n8344 ;
  assign n8346 = x73 | n8344 ;
  assign n21480 = ~n7957 ;
  assign n8347 = n21480 & n7958 ;
  assign n8348 = n150 & n8347 ;
  assign n8349 = n21351 & n8348 ;
  assign n21481 = ~n8348 ;
  assign n8350 = n7963 & n21481 ;
  assign n8351 = n8349 | n8350 ;
  assign n21482 = ~n8351 ;
  assign n8352 = n8346 & n21482 ;
  assign n8353 = n8345 | n8352 ;
  assign n8354 = x74 & n8353 ;
  assign n8355 = x74 | n8353 ;
  assign n21483 = ~n7966 ;
  assign n8356 = n21483 & n7967 ;
  assign n8357 = n150 & n8356 ;
  assign n8358 = n21354 & n8357 ;
  assign n21484 = ~n8357 ;
  assign n8359 = n7972 & n21484 ;
  assign n8360 = n8358 | n8359 ;
  assign n21485 = ~n8360 ;
  assign n8361 = n8355 & n21485 ;
  assign n8362 = n8354 | n8361 ;
  assign n8363 = x75 & n8362 ;
  assign n8364 = x75 | n8362 ;
  assign n21486 = ~n7975 ;
  assign n8365 = n21486 & n7976 ;
  assign n8366 = n150 & n8365 ;
  assign n8367 = n21357 & n8366 ;
  assign n21487 = ~n8366 ;
  assign n8368 = n7981 & n21487 ;
  assign n8369 = n8367 | n8368 ;
  assign n21488 = ~n8369 ;
  assign n8370 = n8364 & n21488 ;
  assign n8371 = n8363 | n8370 ;
  assign n8372 = x76 & n8371 ;
  assign n8373 = x76 | n8371 ;
  assign n21489 = ~n7984 ;
  assign n8374 = n21489 & n7985 ;
  assign n8375 = n150 & n8374 ;
  assign n8376 = n7990 & n8375 ;
  assign n8377 = n7990 | n8375 ;
  assign n21490 = ~n8376 ;
  assign n8378 = n21490 & n8377 ;
  assign n21491 = ~n8378 ;
  assign n8379 = n8373 & n21491 ;
  assign n8380 = n8372 | n8379 ;
  assign n8381 = x77 & n8380 ;
  assign n8382 = x77 | n8380 ;
  assign n21492 = ~n7993 ;
  assign n8383 = n21492 & n7994 ;
  assign n8384 = n150 & n8383 ;
  assign n8385 = n21363 & n8384 ;
  assign n21493 = ~n8384 ;
  assign n8386 = n7999 & n21493 ;
  assign n8387 = n8385 | n8386 ;
  assign n21494 = ~n8387 ;
  assign n8388 = n8382 & n21494 ;
  assign n8389 = n8381 | n8388 ;
  assign n8390 = x78 & n8389 ;
  assign n8391 = x78 | n8389 ;
  assign n21495 = ~n8002 ;
  assign n8392 = n21495 & n8003 ;
  assign n8393 = n150 & n8392 ;
  assign n8394 = n21366 & n8393 ;
  assign n21496 = ~n8393 ;
  assign n8395 = n8008 & n21496 ;
  assign n8396 = n8394 | n8395 ;
  assign n21497 = ~n8396 ;
  assign n8397 = n8391 & n21497 ;
  assign n8398 = n8390 | n8397 ;
  assign n8399 = x79 & n8398 ;
  assign n8400 = x79 | n8398 ;
  assign n21498 = ~n8011 ;
  assign n8401 = n21498 & n8012 ;
  assign n8402 = n150 & n8401 ;
  assign n8403 = n21369 & n8402 ;
  assign n21499 = ~n8402 ;
  assign n8404 = n8017 & n21499 ;
  assign n8405 = n8403 | n8404 ;
  assign n21500 = ~n8405 ;
  assign n8406 = n8400 & n21500 ;
  assign n8407 = n8399 | n8406 ;
  assign n8408 = x80 & n8407 ;
  assign n8409 = x80 | n8407 ;
  assign n21501 = ~n8020 ;
  assign n8410 = n21501 & n8021 ;
  assign n8411 = n150 & n8410 ;
  assign n8412 = n21372 & n8411 ;
  assign n21502 = ~n8411 ;
  assign n8413 = n8026 & n21502 ;
  assign n8414 = n8412 | n8413 ;
  assign n21503 = ~n8414 ;
  assign n8415 = n8409 & n21503 ;
  assign n8416 = n8408 | n8415 ;
  assign n8417 = x81 & n8416 ;
  assign n8418 = x81 | n8416 ;
  assign n21504 = ~n8029 ;
  assign n8419 = n21504 & n8030 ;
  assign n8420 = n150 & n8419 ;
  assign n8421 = n21375 & n8420 ;
  assign n21505 = ~n8420 ;
  assign n8422 = n8035 & n21505 ;
  assign n8423 = n8421 | n8422 ;
  assign n21506 = ~n8423 ;
  assign n8424 = n8418 & n21506 ;
  assign n8425 = n8417 | n8424 ;
  assign n8426 = x82 & n8425 ;
  assign n8427 = x82 | n8425 ;
  assign n21507 = ~n8038 ;
  assign n8428 = n21507 & n8039 ;
  assign n8429 = n150 & n8428 ;
  assign n8430 = n21378 & n8429 ;
  assign n21508 = ~n8429 ;
  assign n8431 = n8044 & n21508 ;
  assign n8432 = n8430 | n8431 ;
  assign n21509 = ~n8432 ;
  assign n8433 = n8427 & n21509 ;
  assign n8434 = n8426 | n8433 ;
  assign n8435 = x83 & n8434 ;
  assign n8436 = x83 | n8434 ;
  assign n21510 = ~n8047 ;
  assign n8437 = n21510 & n8048 ;
  assign n8438 = n150 & n8437 ;
  assign n8439 = n21381 & n8438 ;
  assign n21511 = ~n8438 ;
  assign n8440 = n8053 & n21511 ;
  assign n8441 = n8439 | n8440 ;
  assign n21512 = ~n8441 ;
  assign n8442 = n8436 & n21512 ;
  assign n8443 = n8435 | n8442 ;
  assign n8444 = x84 & n8443 ;
  assign n8445 = x84 | n8443 ;
  assign n21513 = ~n8056 ;
  assign n8446 = n21513 & n8057 ;
  assign n8447 = n150 & n8446 ;
  assign n8448 = n8062 & n8447 ;
  assign n8449 = n8062 | n8447 ;
  assign n21514 = ~n8448 ;
  assign n8450 = n21514 & n8449 ;
  assign n21515 = ~n8450 ;
  assign n8451 = n8445 & n21515 ;
  assign n8452 = n8444 | n8451 ;
  assign n8453 = x85 & n8452 ;
  assign n8454 = x85 | n8452 ;
  assign n21516 = ~n8065 ;
  assign n8455 = n21516 & n8066 ;
  assign n8456 = n150 & n8455 ;
  assign n8457 = n8071 & n8456 ;
  assign n8458 = n8071 | n8456 ;
  assign n21517 = ~n8457 ;
  assign n8459 = n21517 & n8458 ;
  assign n21518 = ~n8459 ;
  assign n8460 = n8454 & n21518 ;
  assign n8461 = n8453 | n8460 ;
  assign n8462 = x86 & n8461 ;
  assign n8463 = x86 | n8461 ;
  assign n21519 = ~n8074 ;
  assign n8464 = n21519 & n8075 ;
  assign n8465 = n150 & n8464 ;
  assign n8466 = n21390 & n8465 ;
  assign n21520 = ~n8465 ;
  assign n8467 = n8080 & n21520 ;
  assign n8468 = n8466 | n8467 ;
  assign n21521 = ~n8468 ;
  assign n8469 = n8463 & n21521 ;
  assign n8470 = n8462 | n8469 ;
  assign n8471 = x87 & n8470 ;
  assign n8472 = x87 | n8470 ;
  assign n21522 = ~n8083 ;
  assign n8473 = n21522 & n8084 ;
  assign n8474 = n150 & n8473 ;
  assign n8475 = n21393 & n8474 ;
  assign n21523 = ~n8474 ;
  assign n8476 = n8089 & n21523 ;
  assign n8477 = n8475 | n8476 ;
  assign n21524 = ~n8477 ;
  assign n8478 = n8472 & n21524 ;
  assign n8479 = n8471 | n8478 ;
  assign n8480 = x88 & n8479 ;
  assign n8481 = x88 | n8479 ;
  assign n21525 = ~n8092 ;
  assign n8482 = n21525 & n8093 ;
  assign n8483 = n150 & n8482 ;
  assign n8484 = n21396 & n8483 ;
  assign n21526 = ~n8483 ;
  assign n8485 = n8098 & n21526 ;
  assign n8486 = n8484 | n8485 ;
  assign n21527 = ~n8486 ;
  assign n8487 = n8481 & n21527 ;
  assign n8488 = n8480 | n8487 ;
  assign n8489 = x89 & n8488 ;
  assign n8490 = x89 | n8488 ;
  assign n21528 = ~n8101 ;
  assign n8491 = n21528 & n8102 ;
  assign n8492 = n150 & n8491 ;
  assign n8493 = n8107 & n8492 ;
  assign n8494 = n8107 | n8492 ;
  assign n21529 = ~n8493 ;
  assign n8495 = n21529 & n8494 ;
  assign n21530 = ~n8495 ;
  assign n8496 = n8490 & n21530 ;
  assign n8497 = n8489 | n8496 ;
  assign n8498 = x90 & n8497 ;
  assign n8499 = x90 | n8497 ;
  assign n21531 = ~n8110 ;
  assign n8500 = n21531 & n8111 ;
  assign n8501 = n150 & n8500 ;
  assign n8502 = n8116 & n8501 ;
  assign n8503 = n8116 | n8501 ;
  assign n21532 = ~n8502 ;
  assign n8504 = n21532 & n8503 ;
  assign n21533 = ~n8504 ;
  assign n8505 = n8499 & n21533 ;
  assign n8506 = n8498 | n8505 ;
  assign n8507 = x91 & n8506 ;
  assign n8508 = x91 | n8506 ;
  assign n21534 = ~n8119 ;
  assign n8509 = n21534 & n8120 ;
  assign n8510 = n150 & n8509 ;
  assign n8511 = n8125 & n8510 ;
  assign n8512 = n8125 | n8510 ;
  assign n21535 = ~n8511 ;
  assign n8513 = n21535 & n8512 ;
  assign n21536 = ~n8513 ;
  assign n8514 = n8508 & n21536 ;
  assign n8515 = n8507 | n8514 ;
  assign n8516 = x92 & n8515 ;
  assign n8517 = x92 | n8515 ;
  assign n21537 = ~n8128 ;
  assign n8518 = n21537 & n8129 ;
  assign n8519 = n150 & n8518 ;
  assign n8520 = n21408 & n8519 ;
  assign n21538 = ~n8519 ;
  assign n8521 = n8134 & n21538 ;
  assign n8522 = n8520 | n8521 ;
  assign n21539 = ~n8522 ;
  assign n8523 = n8517 & n21539 ;
  assign n8524 = n8516 | n8523 ;
  assign n8525 = x93 & n8524 ;
  assign n8526 = x93 | n8524 ;
  assign n21540 = ~n8137 ;
  assign n8527 = n21540 & n8138 ;
  assign n8528 = n150 & n8527 ;
  assign n8529 = n21411 & n8528 ;
  assign n21541 = ~n8528 ;
  assign n8530 = n8143 & n21541 ;
  assign n8531 = n8529 | n8530 ;
  assign n21542 = ~n8531 ;
  assign n8532 = n8526 & n21542 ;
  assign n8533 = n8525 | n8532 ;
  assign n8534 = x94 & n8533 ;
  assign n8535 = x94 | n8533 ;
  assign n21543 = ~n8146 ;
  assign n8536 = n21543 & n8147 ;
  assign n8537 = n150 & n8536 ;
  assign n8538 = n21414 & n8537 ;
  assign n21544 = ~n8537 ;
  assign n8539 = n8152 & n21544 ;
  assign n8540 = n8538 | n8539 ;
  assign n21545 = ~n8540 ;
  assign n8541 = n8535 & n21545 ;
  assign n8542 = n8534 | n8541 ;
  assign n8543 = x95 & n8542 ;
  assign n8544 = x95 | n8542 ;
  assign n21546 = ~n8155 ;
  assign n8545 = n21546 & n8156 ;
  assign n8546 = n150 & n8545 ;
  assign n8547 = n21417 & n8546 ;
  assign n21547 = ~n8546 ;
  assign n8548 = n8161 & n21547 ;
  assign n8549 = n8547 | n8548 ;
  assign n21548 = ~n8549 ;
  assign n8550 = n8544 & n21548 ;
  assign n8551 = n8543 | n8550 ;
  assign n8552 = x96 & n8551 ;
  assign n8553 = x96 | n8551 ;
  assign n21549 = ~n8164 ;
  assign n8554 = n21549 & n8165 ;
  assign n8555 = n150 & n8554 ;
  assign n8556 = n21420 & n8555 ;
  assign n21550 = ~n8555 ;
  assign n8557 = n8170 & n21550 ;
  assign n8558 = n8556 | n8557 ;
  assign n21551 = ~n8558 ;
  assign n8559 = n8553 & n21551 ;
  assign n8560 = n8552 | n8559 ;
  assign n8561 = x97 & n8560 ;
  assign n8562 = x97 | n8560 ;
  assign n21552 = ~n8173 ;
  assign n8563 = n21552 & n8174 ;
  assign n8564 = n150 & n8563 ;
  assign n8565 = n21423 & n8564 ;
  assign n21553 = ~n8564 ;
  assign n8566 = n8179 & n21553 ;
  assign n8567 = n8565 | n8566 ;
  assign n21554 = ~n8567 ;
  assign n8568 = n8562 & n21554 ;
  assign n8569 = n8561 | n8568 ;
  assign n8570 = x98 & n8569 ;
  assign n8571 = x98 | n8569 ;
  assign n21555 = ~n8182 ;
  assign n8572 = n21555 & n8183 ;
  assign n8573 = n150 & n8572 ;
  assign n8574 = n21426 & n8573 ;
  assign n21556 = ~n8573 ;
  assign n8575 = n8188 & n21556 ;
  assign n8576 = n8574 | n8575 ;
  assign n21557 = ~n8576 ;
  assign n8577 = n8571 & n21557 ;
  assign n8578 = n8570 | n8577 ;
  assign n8579 = x99 & n8578 ;
  assign n8580 = x99 | n8578 ;
  assign n21558 = ~n8191 ;
  assign n8581 = n21558 & n8192 ;
  assign n8582 = n150 & n8581 ;
  assign n8583 = n21429 & n8582 ;
  assign n21559 = ~n8582 ;
  assign n8584 = n8197 & n21559 ;
  assign n8585 = n8583 | n8584 ;
  assign n21560 = ~n8585 ;
  assign n8586 = n8580 & n21560 ;
  assign n8587 = n8579 | n8586 ;
  assign n8588 = x100 & n8587 ;
  assign n8589 = x100 | n8587 ;
  assign n21561 = ~n8200 ;
  assign n8590 = n21561 & n8201 ;
  assign n8591 = n150 & n8590 ;
  assign n8592 = n21432 & n8591 ;
  assign n21562 = ~n8591 ;
  assign n8593 = n8206 & n21562 ;
  assign n8594 = n8592 | n8593 ;
  assign n21563 = ~n8594 ;
  assign n8595 = n8589 & n21563 ;
  assign n8596 = n8588 | n8595 ;
  assign n8597 = x101 & n8596 ;
  assign n8598 = x101 | n8596 ;
  assign n21564 = ~n8209 ;
  assign n8599 = n21564 & n8210 ;
  assign n8600 = n150 & n8599 ;
  assign n8601 = n21435 & n8600 ;
  assign n21565 = ~n8600 ;
  assign n8602 = n8215 & n21565 ;
  assign n8603 = n8601 | n8602 ;
  assign n21566 = ~n8603 ;
  assign n8604 = n8598 & n21566 ;
  assign n8605 = n8597 | n8604 ;
  assign n8606 = x102 & n8605 ;
  assign n8607 = x102 | n8605 ;
  assign n21567 = ~n8218 ;
  assign n8608 = n21567 & n8219 ;
  assign n8609 = n150 & n8608 ;
  assign n8610 = n21438 & n8609 ;
  assign n21568 = ~n8609 ;
  assign n8611 = n8224 & n21568 ;
  assign n8612 = n8610 | n8611 ;
  assign n21569 = ~n8612 ;
  assign n8613 = n8607 & n21569 ;
  assign n8614 = n8606 | n8613 ;
  assign n8615 = x103 & n8614 ;
  assign n8616 = x103 | n8614 ;
  assign n21570 = ~n8227 ;
  assign n8617 = n21570 & n8228 ;
  assign n8618 = n150 & n8617 ;
  assign n8619 = n21441 & n8618 ;
  assign n21571 = ~n8618 ;
  assign n8620 = n8233 & n21571 ;
  assign n8621 = n8619 | n8620 ;
  assign n21572 = ~n8621 ;
  assign n8622 = n8616 & n21572 ;
  assign n8623 = n8615 | n8622 ;
  assign n8624 = x104 & n8623 ;
  assign n8625 = x104 | n8623 ;
  assign n21573 = ~n8236 ;
  assign n8626 = n21573 & n8237 ;
  assign n8627 = n150 & n8626 ;
  assign n8628 = n21444 & n8627 ;
  assign n21574 = ~n8627 ;
  assign n8629 = n8242 & n21574 ;
  assign n8630 = n8628 | n8629 ;
  assign n21575 = ~n8630 ;
  assign n8631 = n8625 & n21575 ;
  assign n8632 = n8624 | n8631 ;
  assign n8633 = x105 & n8632 ;
  assign n8634 = x105 | n8632 ;
  assign n21576 = ~n8245 ;
  assign n8635 = n21576 & n8246 ;
  assign n8636 = n150 & n8635 ;
  assign n8637 = n21447 & n8636 ;
  assign n21577 = ~n8636 ;
  assign n8638 = n8251 & n21577 ;
  assign n8639 = n8637 | n8638 ;
  assign n21578 = ~n8639 ;
  assign n8640 = n8634 & n21578 ;
  assign n8641 = n8633 | n8640 ;
  assign n8643 = x106 | n8641 ;
  assign n21579 = ~n8270 ;
  assign n8644 = n21579 & n8643 ;
  assign n8642 = x106 & n8641 ;
  assign n21580 = ~n8259 ;
  assign n8260 = x107 & n21580 ;
  assign n8645 = n18357 | n8260 ;
  assign n8646 = n8272 | n8645 ;
  assign n8647 = n8642 | n8646 ;
  assign n8648 = n8644 | n8647 ;
  assign n21581 = ~n8272 ;
  assign n8649 = n21581 & n8648 ;
  assign n21582 = ~n8642 ;
  assign n8650 = n21582 & n8643 ;
  assign n149 = ~n8649 ;
  assign n8651 = n149 & n8650 ;
  assign n8652 = n21579 & n8651 ;
  assign n21584 = ~n8651 ;
  assign n8653 = n8270 & n21584 ;
  assign n8654 = n8652 | n8653 ;
  assign n21585 = ~x19 ;
  assign n8655 = n21585 & x64 ;
  assign n8656 = x65 | n8655 ;
  assign n8657 = x64 & n149 ;
  assign n21586 = ~n8657 ;
  assign n8658 = x20 & n21586 ;
  assign n8659 = n8273 & n149 ;
  assign n8660 = n8658 | n8659 ;
  assign n8661 = x65 & n8655 ;
  assign n21587 = ~n8661 ;
  assign n8662 = n8660 & n21587 ;
  assign n21588 = ~n8662 ;
  assign n8663 = n8656 & n21588 ;
  assign n8664 = x66 | n8663 ;
  assign n8665 = x66 & n8663 ;
  assign n8666 = n21458 & n8275 ;
  assign n8667 = n149 & n8666 ;
  assign n8668 = n8279 & n8667 ;
  assign n8669 = n8279 | n8667 ;
  assign n21589 = ~n8668 ;
  assign n8670 = n21589 & n8669 ;
  assign n21590 = ~n8665 ;
  assign n8671 = n21590 & n8670 ;
  assign n21591 = ~n8671 ;
  assign n8672 = n8664 & n21591 ;
  assign n8674 = x67 | n8672 ;
  assign n8673 = x67 & n8672 ;
  assign n21592 = ~n8282 ;
  assign n8675 = n21592 & n8283 ;
  assign n8676 = n149 & n8675 ;
  assign n8677 = n8288 & n8676 ;
  assign n8678 = n8288 | n8676 ;
  assign n21593 = ~n8677 ;
  assign n8679 = n21593 & n8678 ;
  assign n21594 = ~n8673 ;
  assign n8680 = n21594 & n8679 ;
  assign n21595 = ~n8680 ;
  assign n8681 = n8674 & n21595 ;
  assign n8682 = x68 | n8681 ;
  assign n8683 = x68 & n8681 ;
  assign n21596 = ~n8291 ;
  assign n8684 = n21596 & n8292 ;
  assign n8685 = n149 & n8684 ;
  assign n8686 = n8297 & n8685 ;
  assign n8687 = n8297 | n8685 ;
  assign n21597 = ~n8686 ;
  assign n8688 = n21597 & n8687 ;
  assign n21598 = ~n8683 ;
  assign n8689 = n21598 & n8688 ;
  assign n21599 = ~n8689 ;
  assign n8690 = n8682 & n21599 ;
  assign n8691 = x69 | n8690 ;
  assign n8692 = x69 & n8690 ;
  assign n21600 = ~n8300 ;
  assign n8693 = n21600 & n8301 ;
  assign n8694 = n149 & n8693 ;
  assign n8695 = n8306 & n8694 ;
  assign n8696 = n8306 | n8694 ;
  assign n21601 = ~n8695 ;
  assign n8697 = n21601 & n8696 ;
  assign n21602 = ~n8692 ;
  assign n8698 = n21602 & n8697 ;
  assign n21603 = ~n8698 ;
  assign n8699 = n8691 & n21603 ;
  assign n8700 = x70 | n8699 ;
  assign n8701 = x70 & n8699 ;
  assign n21604 = ~n8309 ;
  assign n8702 = n21604 & n8310 ;
  assign n8703 = n149 & n8702 ;
  assign n8704 = n21470 & n8703 ;
  assign n21605 = ~n8703 ;
  assign n8705 = n8315 & n21605 ;
  assign n8706 = n8704 | n8705 ;
  assign n21606 = ~n8701 ;
  assign n8707 = n21606 & n8706 ;
  assign n21607 = ~n8707 ;
  assign n8708 = n8700 & n21607 ;
  assign n8709 = x71 | n8708 ;
  assign n8710 = x71 & n8708 ;
  assign n21608 = ~n8318 ;
  assign n8711 = n21608 & n8319 ;
  assign n8712 = n149 & n8711 ;
  assign n8713 = n8324 & n8712 ;
  assign n8714 = n8324 | n8712 ;
  assign n21609 = ~n8713 ;
  assign n8715 = n21609 & n8714 ;
  assign n21610 = ~n8710 ;
  assign n8716 = n21610 & n8715 ;
  assign n21611 = ~n8716 ;
  assign n8717 = n8709 & n21611 ;
  assign n8718 = x72 | n8717 ;
  assign n8719 = x72 & n8717 ;
  assign n21612 = ~n8327 ;
  assign n8720 = n21612 & n8328 ;
  assign n8721 = n149 & n8720 ;
  assign n8722 = n8333 & n8721 ;
  assign n8723 = n8333 | n8721 ;
  assign n21613 = ~n8722 ;
  assign n8724 = n21613 & n8723 ;
  assign n21614 = ~n8719 ;
  assign n8725 = n21614 & n8724 ;
  assign n21615 = ~n8725 ;
  assign n8726 = n8718 & n21615 ;
  assign n8727 = x73 | n8726 ;
  assign n8728 = x73 & n8726 ;
  assign n21616 = ~n8336 ;
  assign n8729 = n21616 & n8337 ;
  assign n8730 = n149 & n8729 ;
  assign n8731 = n21479 & n8730 ;
  assign n21617 = ~n8730 ;
  assign n8732 = n8342 & n21617 ;
  assign n8733 = n8731 | n8732 ;
  assign n21618 = ~n8728 ;
  assign n8734 = n21618 & n8733 ;
  assign n21619 = ~n8734 ;
  assign n8735 = n8727 & n21619 ;
  assign n8736 = x74 | n8735 ;
  assign n8737 = x74 & n8735 ;
  assign n21620 = ~n8345 ;
  assign n8738 = n21620 & n8346 ;
  assign n8739 = n149 & n8738 ;
  assign n8740 = n21482 & n8739 ;
  assign n21621 = ~n8739 ;
  assign n8741 = n8351 & n21621 ;
  assign n8742 = n8740 | n8741 ;
  assign n21622 = ~n8737 ;
  assign n8743 = n21622 & n8742 ;
  assign n21623 = ~n8743 ;
  assign n8744 = n8736 & n21623 ;
  assign n8745 = x75 | n8744 ;
  assign n8746 = x75 & n8744 ;
  assign n21624 = ~n8354 ;
  assign n8747 = n21624 & n8355 ;
  assign n8748 = n149 & n8747 ;
  assign n8749 = n8360 & n8748 ;
  assign n8750 = n8360 | n8748 ;
  assign n21625 = ~n8749 ;
  assign n8751 = n21625 & n8750 ;
  assign n21626 = ~n8746 ;
  assign n8752 = n21626 & n8751 ;
  assign n21627 = ~n8752 ;
  assign n8753 = n8745 & n21627 ;
  assign n8754 = x76 | n8753 ;
  assign n8755 = x76 & n8753 ;
  assign n21628 = ~n8363 ;
  assign n8756 = n21628 & n8364 ;
  assign n8757 = n149 & n8756 ;
  assign n8758 = n8369 & n8757 ;
  assign n8759 = n8369 | n8757 ;
  assign n21629 = ~n8758 ;
  assign n8760 = n21629 & n8759 ;
  assign n21630 = ~n8755 ;
  assign n8761 = n21630 & n8760 ;
  assign n21631 = ~n8761 ;
  assign n8762 = n8754 & n21631 ;
  assign n8763 = x77 | n8762 ;
  assign n8764 = x77 & n8762 ;
  assign n21632 = ~n8372 ;
  assign n8765 = n21632 & n8373 ;
  assign n8766 = n149 & n8765 ;
  assign n8767 = n8378 & n8766 ;
  assign n8768 = n8378 | n8766 ;
  assign n21633 = ~n8767 ;
  assign n8769 = n21633 & n8768 ;
  assign n21634 = ~n8764 ;
  assign n8770 = n21634 & n8769 ;
  assign n21635 = ~n8770 ;
  assign n8771 = n8763 & n21635 ;
  assign n8772 = x78 | n8771 ;
  assign n8773 = x78 & n8771 ;
  assign n21636 = ~n8381 ;
  assign n8774 = n21636 & n8382 ;
  assign n8775 = n149 & n8774 ;
  assign n8776 = n21494 & n8775 ;
  assign n21637 = ~n8775 ;
  assign n8777 = n8387 & n21637 ;
  assign n8778 = n8776 | n8777 ;
  assign n21638 = ~n8773 ;
  assign n8779 = n21638 & n8778 ;
  assign n21639 = ~n8779 ;
  assign n8780 = n8772 & n21639 ;
  assign n8781 = x79 | n8780 ;
  assign n8782 = x79 & n8780 ;
  assign n21640 = ~n8390 ;
  assign n8783 = n21640 & n8391 ;
  assign n8784 = n149 & n8783 ;
  assign n8785 = n21497 & n8784 ;
  assign n21641 = ~n8784 ;
  assign n8786 = n8396 & n21641 ;
  assign n8787 = n8785 | n8786 ;
  assign n21642 = ~n8782 ;
  assign n8788 = n21642 & n8787 ;
  assign n21643 = ~n8788 ;
  assign n8789 = n8781 & n21643 ;
  assign n8790 = x80 | n8789 ;
  assign n8791 = x80 & n8789 ;
  assign n21644 = ~n8399 ;
  assign n8792 = n21644 & n8400 ;
  assign n8793 = n149 & n8792 ;
  assign n8794 = n21500 & n8793 ;
  assign n21645 = ~n8793 ;
  assign n8795 = n8405 & n21645 ;
  assign n8796 = n8794 | n8795 ;
  assign n21646 = ~n8791 ;
  assign n8797 = n21646 & n8796 ;
  assign n21647 = ~n8797 ;
  assign n8798 = n8790 & n21647 ;
  assign n8799 = x81 | n8798 ;
  assign n8800 = x81 & n8798 ;
  assign n21648 = ~n8408 ;
  assign n8801 = n21648 & n8409 ;
  assign n8802 = n149 & n8801 ;
  assign n8803 = n21503 & n8802 ;
  assign n21649 = ~n8802 ;
  assign n8804 = n8414 & n21649 ;
  assign n8805 = n8803 | n8804 ;
  assign n21650 = ~n8800 ;
  assign n8806 = n21650 & n8805 ;
  assign n21651 = ~n8806 ;
  assign n8807 = n8799 & n21651 ;
  assign n8808 = x82 | n8807 ;
  assign n8809 = x82 & n8807 ;
  assign n21652 = ~n8417 ;
  assign n8810 = n21652 & n8418 ;
  assign n8811 = n149 & n8810 ;
  assign n8812 = n21506 & n8811 ;
  assign n21653 = ~n8811 ;
  assign n8813 = n8423 & n21653 ;
  assign n8814 = n8812 | n8813 ;
  assign n21654 = ~n8809 ;
  assign n8815 = n21654 & n8814 ;
  assign n21655 = ~n8815 ;
  assign n8816 = n8808 & n21655 ;
  assign n8817 = x83 | n8816 ;
  assign n8818 = x83 & n8816 ;
  assign n21656 = ~n8426 ;
  assign n8819 = n21656 & n8427 ;
  assign n8820 = n149 & n8819 ;
  assign n8821 = n21509 & n8820 ;
  assign n21657 = ~n8820 ;
  assign n8822 = n8432 & n21657 ;
  assign n8823 = n8821 | n8822 ;
  assign n21658 = ~n8818 ;
  assign n8824 = n21658 & n8823 ;
  assign n21659 = ~n8824 ;
  assign n8825 = n8817 & n21659 ;
  assign n8826 = x84 | n8825 ;
  assign n8827 = x84 & n8825 ;
  assign n21660 = ~n8435 ;
  assign n8828 = n21660 & n8436 ;
  assign n8829 = n149 & n8828 ;
  assign n8830 = n21512 & n8829 ;
  assign n21661 = ~n8829 ;
  assign n8831 = n8441 & n21661 ;
  assign n8832 = n8830 | n8831 ;
  assign n21662 = ~n8827 ;
  assign n8833 = n21662 & n8832 ;
  assign n21663 = ~n8833 ;
  assign n8834 = n8826 & n21663 ;
  assign n8835 = x85 | n8834 ;
  assign n8836 = x85 & n8834 ;
  assign n21664 = ~n8444 ;
  assign n8837 = n21664 & n8445 ;
  assign n8838 = n149 & n8837 ;
  assign n8839 = n21515 & n8838 ;
  assign n21665 = ~n8838 ;
  assign n8840 = n8450 & n21665 ;
  assign n8841 = n8839 | n8840 ;
  assign n21666 = ~n8836 ;
  assign n8842 = n21666 & n8841 ;
  assign n21667 = ~n8842 ;
  assign n8843 = n8835 & n21667 ;
  assign n8844 = x86 | n8843 ;
  assign n8845 = x86 & n8843 ;
  assign n21668 = ~n8453 ;
  assign n8846 = n21668 & n8454 ;
  assign n8847 = n149 & n8846 ;
  assign n8848 = n8459 & n8847 ;
  assign n8849 = n8459 | n8847 ;
  assign n21669 = ~n8848 ;
  assign n8850 = n21669 & n8849 ;
  assign n21670 = ~n8845 ;
  assign n8851 = n21670 & n8850 ;
  assign n21671 = ~n8851 ;
  assign n8852 = n8844 & n21671 ;
  assign n8853 = x87 | n8852 ;
  assign n8854 = x87 & n8852 ;
  assign n21672 = ~n8462 ;
  assign n8855 = n21672 & n8463 ;
  assign n8856 = n149 & n8855 ;
  assign n8857 = n21521 & n8856 ;
  assign n21673 = ~n8856 ;
  assign n8858 = n8468 & n21673 ;
  assign n8859 = n8857 | n8858 ;
  assign n21674 = ~n8854 ;
  assign n8860 = n21674 & n8859 ;
  assign n21675 = ~n8860 ;
  assign n8861 = n8853 & n21675 ;
  assign n8862 = x88 | n8861 ;
  assign n8863 = x88 & n8861 ;
  assign n21676 = ~n8471 ;
  assign n8864 = n21676 & n8472 ;
  assign n8865 = n149 & n8864 ;
  assign n8866 = n8477 & n8865 ;
  assign n8867 = n8477 | n8865 ;
  assign n21677 = ~n8866 ;
  assign n8868 = n21677 & n8867 ;
  assign n21678 = ~n8863 ;
  assign n8869 = n21678 & n8868 ;
  assign n21679 = ~n8869 ;
  assign n8870 = n8862 & n21679 ;
  assign n8871 = x89 | n8870 ;
  assign n8872 = x89 & n8870 ;
  assign n21680 = ~n8480 ;
  assign n8873 = n21680 & n8481 ;
  assign n8874 = n149 & n8873 ;
  assign n8875 = n8486 & n8874 ;
  assign n8876 = n8486 | n8874 ;
  assign n21681 = ~n8875 ;
  assign n8877 = n21681 & n8876 ;
  assign n21682 = ~n8872 ;
  assign n8878 = n21682 & n8877 ;
  assign n21683 = ~n8878 ;
  assign n8879 = n8871 & n21683 ;
  assign n8880 = x90 | n8879 ;
  assign n8881 = x90 & n8879 ;
  assign n21684 = ~n8489 ;
  assign n8882 = n21684 & n8490 ;
  assign n8883 = n149 & n8882 ;
  assign n8884 = n8495 & n8883 ;
  assign n8885 = n8495 | n8883 ;
  assign n21685 = ~n8884 ;
  assign n8886 = n21685 & n8885 ;
  assign n21686 = ~n8881 ;
  assign n8887 = n21686 & n8886 ;
  assign n21687 = ~n8887 ;
  assign n8888 = n8880 & n21687 ;
  assign n8889 = x91 | n8888 ;
  assign n8890 = x91 & n8888 ;
  assign n21688 = ~n8498 ;
  assign n8891 = n21688 & n8499 ;
  assign n8892 = n149 & n8891 ;
  assign n8893 = n8504 & n8892 ;
  assign n8894 = n8504 | n8892 ;
  assign n21689 = ~n8893 ;
  assign n8895 = n21689 & n8894 ;
  assign n21690 = ~n8890 ;
  assign n8896 = n21690 & n8895 ;
  assign n21691 = ~n8896 ;
  assign n8897 = n8889 & n21691 ;
  assign n8898 = x92 | n8897 ;
  assign n8899 = x92 & n8897 ;
  assign n21692 = ~n8507 ;
  assign n8900 = n21692 & n8508 ;
  assign n8901 = n149 & n8900 ;
  assign n8902 = n8513 & n8901 ;
  assign n8903 = n8513 | n8901 ;
  assign n21693 = ~n8902 ;
  assign n8904 = n21693 & n8903 ;
  assign n21694 = ~n8899 ;
  assign n8905 = n21694 & n8904 ;
  assign n21695 = ~n8905 ;
  assign n8906 = n8898 & n21695 ;
  assign n8907 = x93 | n8906 ;
  assign n8908 = x93 & n8906 ;
  assign n21696 = ~n8516 ;
  assign n8909 = n21696 & n8517 ;
  assign n8910 = n149 & n8909 ;
  assign n8911 = n21539 & n8910 ;
  assign n21697 = ~n8910 ;
  assign n8912 = n8522 & n21697 ;
  assign n8913 = n8911 | n8912 ;
  assign n21698 = ~n8908 ;
  assign n8914 = n21698 & n8913 ;
  assign n21699 = ~n8914 ;
  assign n8915 = n8907 & n21699 ;
  assign n8916 = x94 | n8915 ;
  assign n8917 = x94 & n8915 ;
  assign n21700 = ~n8525 ;
  assign n8918 = n21700 & n8526 ;
  assign n8919 = n149 & n8918 ;
  assign n8920 = n21542 & n8919 ;
  assign n21701 = ~n8919 ;
  assign n8921 = n8531 & n21701 ;
  assign n8922 = n8920 | n8921 ;
  assign n21702 = ~n8917 ;
  assign n8923 = n21702 & n8922 ;
  assign n21703 = ~n8923 ;
  assign n8924 = n8916 & n21703 ;
  assign n8925 = x95 | n8924 ;
  assign n8926 = x95 & n8924 ;
  assign n21704 = ~n8534 ;
  assign n8927 = n21704 & n8535 ;
  assign n8928 = n149 & n8927 ;
  assign n8929 = n21545 & n8928 ;
  assign n21705 = ~n8928 ;
  assign n8930 = n8540 & n21705 ;
  assign n8931 = n8929 | n8930 ;
  assign n21706 = ~n8926 ;
  assign n8932 = n21706 & n8931 ;
  assign n21707 = ~n8932 ;
  assign n8933 = n8925 & n21707 ;
  assign n8934 = x96 | n8933 ;
  assign n8935 = x96 & n8933 ;
  assign n21708 = ~n8543 ;
  assign n8936 = n21708 & n8544 ;
  assign n8937 = n149 & n8936 ;
  assign n8938 = n21548 & n8937 ;
  assign n21709 = ~n8937 ;
  assign n8939 = n8549 & n21709 ;
  assign n8940 = n8938 | n8939 ;
  assign n21710 = ~n8935 ;
  assign n8941 = n21710 & n8940 ;
  assign n21711 = ~n8941 ;
  assign n8942 = n8934 & n21711 ;
  assign n8943 = x97 | n8942 ;
  assign n8944 = x97 & n8942 ;
  assign n21712 = ~n8552 ;
  assign n8945 = n21712 & n8553 ;
  assign n8946 = n149 & n8945 ;
  assign n8947 = n21551 & n8946 ;
  assign n21713 = ~n8946 ;
  assign n8948 = n8558 & n21713 ;
  assign n8949 = n8947 | n8948 ;
  assign n21714 = ~n8944 ;
  assign n8950 = n21714 & n8949 ;
  assign n21715 = ~n8950 ;
  assign n8951 = n8943 & n21715 ;
  assign n8952 = x98 | n8951 ;
  assign n8953 = x98 & n8951 ;
  assign n21716 = ~n8561 ;
  assign n8954 = n21716 & n8562 ;
  assign n8955 = n149 & n8954 ;
  assign n8956 = n21554 & n8955 ;
  assign n21717 = ~n8955 ;
  assign n8957 = n8567 & n21717 ;
  assign n8958 = n8956 | n8957 ;
  assign n21718 = ~n8953 ;
  assign n8959 = n21718 & n8958 ;
  assign n21719 = ~n8959 ;
  assign n8960 = n8952 & n21719 ;
  assign n8961 = x99 | n8960 ;
  assign n8962 = x99 & n8960 ;
  assign n21720 = ~n8570 ;
  assign n8963 = n21720 & n8571 ;
  assign n8964 = n149 & n8963 ;
  assign n8965 = n21557 & n8964 ;
  assign n21721 = ~n8964 ;
  assign n8966 = n8576 & n21721 ;
  assign n8967 = n8965 | n8966 ;
  assign n21722 = ~n8962 ;
  assign n8968 = n21722 & n8967 ;
  assign n21723 = ~n8968 ;
  assign n8969 = n8961 & n21723 ;
  assign n8970 = x100 | n8969 ;
  assign n8971 = x100 & n8969 ;
  assign n21724 = ~n8579 ;
  assign n8972 = n21724 & n8580 ;
  assign n8973 = n149 & n8972 ;
  assign n8974 = n21560 & n8973 ;
  assign n21725 = ~n8973 ;
  assign n8975 = n8585 & n21725 ;
  assign n8976 = n8974 | n8975 ;
  assign n21726 = ~n8971 ;
  assign n8977 = n21726 & n8976 ;
  assign n21727 = ~n8977 ;
  assign n8978 = n8970 & n21727 ;
  assign n8979 = x101 | n8978 ;
  assign n8980 = x101 & n8978 ;
  assign n21728 = ~n8588 ;
  assign n8981 = n21728 & n8589 ;
  assign n8982 = n149 & n8981 ;
  assign n8983 = n21563 & n8982 ;
  assign n21729 = ~n8982 ;
  assign n8984 = n8594 & n21729 ;
  assign n8985 = n8983 | n8984 ;
  assign n21730 = ~n8980 ;
  assign n8986 = n21730 & n8985 ;
  assign n21731 = ~n8986 ;
  assign n8987 = n8979 & n21731 ;
  assign n8988 = x102 | n8987 ;
  assign n8989 = x102 & n8987 ;
  assign n21732 = ~n8597 ;
  assign n8990 = n21732 & n8598 ;
  assign n8991 = n149 & n8990 ;
  assign n8992 = n21566 & n8991 ;
  assign n21733 = ~n8991 ;
  assign n8993 = n8603 & n21733 ;
  assign n8994 = n8992 | n8993 ;
  assign n21734 = ~n8989 ;
  assign n8995 = n21734 & n8994 ;
  assign n21735 = ~n8995 ;
  assign n8996 = n8988 & n21735 ;
  assign n8997 = x103 | n8996 ;
  assign n8998 = x103 & n8996 ;
  assign n21736 = ~n8606 ;
  assign n8999 = n21736 & n8607 ;
  assign n9000 = n149 & n8999 ;
  assign n9001 = n21569 & n9000 ;
  assign n21737 = ~n9000 ;
  assign n9002 = n8612 & n21737 ;
  assign n9003 = n9001 | n9002 ;
  assign n21738 = ~n8998 ;
  assign n9004 = n21738 & n9003 ;
  assign n21739 = ~n9004 ;
  assign n9005 = n8997 & n21739 ;
  assign n9006 = x104 | n9005 ;
  assign n9007 = x104 & n9005 ;
  assign n21740 = ~n8615 ;
  assign n9008 = n21740 & n8616 ;
  assign n9009 = n149 & n9008 ;
  assign n9010 = n21572 & n9009 ;
  assign n21741 = ~n9009 ;
  assign n9011 = n8621 & n21741 ;
  assign n9012 = n9010 | n9011 ;
  assign n21742 = ~n9007 ;
  assign n9013 = n21742 & n9012 ;
  assign n21743 = ~n9013 ;
  assign n9014 = n9006 & n21743 ;
  assign n9015 = x105 | n9014 ;
  assign n9016 = x105 & n9014 ;
  assign n21744 = ~n8624 ;
  assign n9017 = n21744 & n8625 ;
  assign n9018 = n149 & n9017 ;
  assign n9019 = n21575 & n9018 ;
  assign n21745 = ~n9018 ;
  assign n9020 = n8630 & n21745 ;
  assign n9021 = n9019 | n9020 ;
  assign n21746 = ~n9016 ;
  assign n9022 = n21746 & n9021 ;
  assign n21747 = ~n9022 ;
  assign n9023 = n9015 & n21747 ;
  assign n9024 = x106 | n9023 ;
  assign n9025 = x106 & n9023 ;
  assign n21748 = ~n8633 ;
  assign n9026 = n21748 & n8634 ;
  assign n9027 = n149 & n9026 ;
  assign n9028 = n21578 & n9027 ;
  assign n21749 = ~n9027 ;
  assign n9029 = n8639 & n21749 ;
  assign n9030 = n9028 | n9029 ;
  assign n21750 = ~n9025 ;
  assign n9031 = n21750 & n9030 ;
  assign n21751 = ~n9031 ;
  assign n9032 = n9024 & n21751 ;
  assign n9033 = x107 | n9032 ;
  assign n9034 = x107 & n9032 ;
  assign n21752 = ~n9034 ;
  assign n9035 = n8654 & n21752 ;
  assign n21753 = ~n9035 ;
  assign n9036 = n9033 & n21753 ;
  assign n9038 = x108 & n9036 ;
  assign n9039 = n18353 | n9038 ;
  assign n9037 = x108 | n9036 ;
  assign n9040 = n8259 & n8648 ;
  assign n9041 = n18363 & n9040 ;
  assign n9043 = n21884 | n9041 ;
  assign n21754 = ~n9043 ;
  assign n9044 = n9037 & n21754 ;
  assign n9045 = n9039 | n9044 ;
  assign n9049 = n9033 & n21752 ;
  assign n148 = ~n9045 ;
  assign n9050 = n148 & n9049 ;
  assign n21756 = ~n8654 ;
  assign n9051 = n21756 & n9050 ;
  assign n21757 = ~n9050 ;
  assign n9052 = n8654 & n21757 ;
  assign n9053 = n9051 | n9052 ;
  assign n9042 = n9039 & n9040 ;
  assign n9054 = n21884 | n9042 ;
  assign n21758 = ~n9054 ;
  assign n9055 = x109 & n21758 ;
  assign n21759 = ~x109 ;
  assign n9057 = n21759 & n9054 ;
  assign n21760 = ~x18 ;
  assign n9058 = n21760 & x64 ;
  assign n9060 = x65 | n9058 ;
  assign n9059 = x65 & n9058 ;
  assign n9061 = x64 & n148 ;
  assign n9062 = x19 & n9061 ;
  assign n9063 = x19 | n9061 ;
  assign n21761 = ~n9062 ;
  assign n9064 = n21761 & n9063 ;
  assign n21762 = ~n9059 ;
  assign n9065 = n21762 & n9064 ;
  assign n21763 = ~n9065 ;
  assign n9066 = n9060 & n21763 ;
  assign n9067 = x66 | n9066 ;
  assign n9068 = x66 & n9066 ;
  assign n9046 = n8656 & n148 ;
  assign n9069 = n21587 & n9046 ;
  assign n9070 = n8660 | n9069 ;
  assign n9071 = n8662 & n9046 ;
  assign n21764 = ~n9071 ;
  assign n9072 = n9070 & n21764 ;
  assign n21765 = ~n9068 ;
  assign n9073 = n21765 & n9072 ;
  assign n21766 = ~n9073 ;
  assign n9074 = n9067 & n21766 ;
  assign n9076 = x67 & n9074 ;
  assign n9075 = x67 | n9074 ;
  assign n9047 = n8664 & n148 ;
  assign n9048 = n8671 & n9047 ;
  assign n9077 = n21590 & n9047 ;
  assign n9078 = n8670 | n9077 ;
  assign n21767 = ~n9048 ;
  assign n9079 = n21767 & n9078 ;
  assign n21768 = ~n9079 ;
  assign n9080 = n9075 & n21768 ;
  assign n9081 = n9076 | n9080 ;
  assign n9082 = x68 & n9081 ;
  assign n9083 = x68 | n9081 ;
  assign n9084 = n8674 & n148 ;
  assign n9085 = n8680 & n9084 ;
  assign n9086 = n21594 & n9084 ;
  assign n9087 = n8679 | n9086 ;
  assign n21769 = ~n9085 ;
  assign n9088 = n21769 & n9087 ;
  assign n21770 = ~n9088 ;
  assign n9089 = n9083 & n21770 ;
  assign n9090 = n9082 | n9089 ;
  assign n9091 = x69 & n9090 ;
  assign n9092 = x69 | n9090 ;
  assign n9093 = n8682 & n21598 ;
  assign n9094 = n148 & n9093 ;
  assign n21771 = ~n8688 ;
  assign n9095 = n21771 & n9094 ;
  assign n21772 = ~n9094 ;
  assign n9096 = n8688 & n21772 ;
  assign n9097 = n9095 | n9096 ;
  assign n21773 = ~n9097 ;
  assign n9098 = n9092 & n21773 ;
  assign n9099 = n9091 | n9098 ;
  assign n9100 = x70 & n9099 ;
  assign n9101 = x70 | n9099 ;
  assign n9102 = n8691 & n21602 ;
  assign n9103 = n148 & n9102 ;
  assign n9104 = n8697 & n9103 ;
  assign n9105 = n8697 | n9103 ;
  assign n21774 = ~n9104 ;
  assign n9106 = n21774 & n9105 ;
  assign n21775 = ~n9106 ;
  assign n9107 = n9101 & n21775 ;
  assign n9108 = n9100 | n9107 ;
  assign n9109 = x71 & n9108 ;
  assign n9110 = x71 | n9108 ;
  assign n9111 = n8700 & n21606 ;
  assign n9112 = n148 & n9111 ;
  assign n21776 = ~n8706 ;
  assign n9113 = n21776 & n9112 ;
  assign n21777 = ~n9112 ;
  assign n9114 = n8706 & n21777 ;
  assign n9115 = n9113 | n9114 ;
  assign n21778 = ~n9115 ;
  assign n9116 = n9110 & n21778 ;
  assign n9117 = n9109 | n9116 ;
  assign n9118 = x72 & n9117 ;
  assign n9119 = x72 | n9117 ;
  assign n9120 = n8709 & n21610 ;
  assign n9121 = n148 & n9120 ;
  assign n21779 = ~n8715 ;
  assign n9122 = n21779 & n9121 ;
  assign n21780 = ~n9121 ;
  assign n9123 = n8715 & n21780 ;
  assign n9124 = n9122 | n9123 ;
  assign n21781 = ~n9124 ;
  assign n9125 = n9119 & n21781 ;
  assign n9126 = n9118 | n9125 ;
  assign n9127 = x73 & n9126 ;
  assign n9128 = x73 | n9126 ;
  assign n9129 = n8718 & n21614 ;
  assign n9130 = n148 & n9129 ;
  assign n9131 = n8724 & n9130 ;
  assign n9132 = n8724 | n9130 ;
  assign n21782 = ~n9131 ;
  assign n9133 = n21782 & n9132 ;
  assign n21783 = ~n9133 ;
  assign n9134 = n9128 & n21783 ;
  assign n9135 = n9127 | n9134 ;
  assign n9136 = x74 & n9135 ;
  assign n9137 = x74 | n9135 ;
  assign n9138 = n8727 & n21618 ;
  assign n9139 = n148 & n9138 ;
  assign n21784 = ~n8733 ;
  assign n9140 = n21784 & n9139 ;
  assign n21785 = ~n9139 ;
  assign n9141 = n8733 & n21785 ;
  assign n9142 = n9140 | n9141 ;
  assign n21786 = ~n9142 ;
  assign n9143 = n9137 & n21786 ;
  assign n9144 = n9136 | n9143 ;
  assign n9145 = x75 & n9144 ;
  assign n9146 = x75 | n9144 ;
  assign n9147 = n8736 & n21622 ;
  assign n9148 = n148 & n9147 ;
  assign n21787 = ~n8742 ;
  assign n9149 = n21787 & n9148 ;
  assign n21788 = ~n9148 ;
  assign n9150 = n8742 & n21788 ;
  assign n9151 = n9149 | n9150 ;
  assign n21789 = ~n9151 ;
  assign n9152 = n9146 & n21789 ;
  assign n9153 = n9145 | n9152 ;
  assign n9154 = x76 & n9153 ;
  assign n9155 = x76 | n9153 ;
  assign n9156 = n8745 & n21626 ;
  assign n9157 = n148 & n9156 ;
  assign n9158 = n8751 & n9157 ;
  assign n9159 = n8751 | n9157 ;
  assign n21790 = ~n9158 ;
  assign n9160 = n21790 & n9159 ;
  assign n21791 = ~n9160 ;
  assign n9161 = n9155 & n21791 ;
  assign n9162 = n9154 | n9161 ;
  assign n9163 = x77 & n9162 ;
  assign n9164 = x77 | n9162 ;
  assign n9165 = n8754 & n21630 ;
  assign n9166 = n148 & n9165 ;
  assign n9167 = n8760 & n9166 ;
  assign n9168 = n8760 | n9166 ;
  assign n21792 = ~n9167 ;
  assign n9169 = n21792 & n9168 ;
  assign n21793 = ~n9169 ;
  assign n9170 = n9164 & n21793 ;
  assign n9171 = n9163 | n9170 ;
  assign n9172 = x78 & n9171 ;
  assign n9173 = x78 | n9171 ;
  assign n9174 = n8763 & n21634 ;
  assign n9175 = n148 & n9174 ;
  assign n21794 = ~n8769 ;
  assign n9176 = n21794 & n9175 ;
  assign n21795 = ~n9175 ;
  assign n9177 = n8769 & n21795 ;
  assign n9178 = n9176 | n9177 ;
  assign n21796 = ~n9178 ;
  assign n9179 = n9173 & n21796 ;
  assign n9180 = n9172 | n9179 ;
  assign n9181 = x79 & n9180 ;
  assign n9182 = x79 | n9180 ;
  assign n9183 = n8772 & n21638 ;
  assign n9184 = n148 & n9183 ;
  assign n21797 = ~n8778 ;
  assign n9185 = n21797 & n9184 ;
  assign n21798 = ~n9184 ;
  assign n9186 = n8778 & n21798 ;
  assign n9187 = n9185 | n9186 ;
  assign n21799 = ~n9187 ;
  assign n9188 = n9182 & n21799 ;
  assign n9189 = n9181 | n9188 ;
  assign n9190 = x80 & n9189 ;
  assign n9191 = x80 | n9189 ;
  assign n9192 = n8781 & n21642 ;
  assign n9193 = n148 & n9192 ;
  assign n21800 = ~n8787 ;
  assign n9194 = n21800 & n9193 ;
  assign n21801 = ~n9193 ;
  assign n9195 = n8787 & n21801 ;
  assign n9196 = n9194 | n9195 ;
  assign n21802 = ~n9196 ;
  assign n9197 = n9191 & n21802 ;
  assign n9198 = n9190 | n9197 ;
  assign n9199 = x81 & n9198 ;
  assign n9200 = x81 | n9198 ;
  assign n9201 = n8790 & n21646 ;
  assign n9202 = n148 & n9201 ;
  assign n21803 = ~n8796 ;
  assign n9203 = n21803 & n9202 ;
  assign n21804 = ~n9202 ;
  assign n9204 = n8796 & n21804 ;
  assign n9205 = n9203 | n9204 ;
  assign n21805 = ~n9205 ;
  assign n9206 = n9200 & n21805 ;
  assign n9207 = n9199 | n9206 ;
  assign n9208 = x82 & n9207 ;
  assign n9209 = x82 | n9207 ;
  assign n9210 = n8799 & n21650 ;
  assign n9211 = n148 & n9210 ;
  assign n21806 = ~n8805 ;
  assign n9212 = n21806 & n9211 ;
  assign n21807 = ~n9211 ;
  assign n9213 = n8805 & n21807 ;
  assign n9214 = n9212 | n9213 ;
  assign n21808 = ~n9214 ;
  assign n9215 = n9209 & n21808 ;
  assign n9216 = n9208 | n9215 ;
  assign n9217 = x83 & n9216 ;
  assign n9218 = x83 | n9216 ;
  assign n9219 = n8808 & n21654 ;
  assign n9220 = n148 & n9219 ;
  assign n21809 = ~n8814 ;
  assign n9221 = n21809 & n9220 ;
  assign n21810 = ~n9220 ;
  assign n9222 = n8814 & n21810 ;
  assign n9223 = n9221 | n9222 ;
  assign n21811 = ~n9223 ;
  assign n9224 = n9218 & n21811 ;
  assign n9225 = n9217 | n9224 ;
  assign n9226 = x84 & n9225 ;
  assign n9227 = x84 | n9225 ;
  assign n9228 = n8817 & n21658 ;
  assign n9229 = n148 & n9228 ;
  assign n21812 = ~n8823 ;
  assign n9230 = n21812 & n9229 ;
  assign n21813 = ~n9229 ;
  assign n9231 = n8823 & n21813 ;
  assign n9232 = n9230 | n9231 ;
  assign n21814 = ~n9232 ;
  assign n9233 = n9227 & n21814 ;
  assign n9234 = n9226 | n9233 ;
  assign n9235 = x85 & n9234 ;
  assign n9236 = x85 | n9234 ;
  assign n9237 = n8826 & n21662 ;
  assign n9238 = n148 & n9237 ;
  assign n21815 = ~n8832 ;
  assign n9239 = n21815 & n9238 ;
  assign n21816 = ~n9238 ;
  assign n9240 = n8832 & n21816 ;
  assign n9241 = n9239 | n9240 ;
  assign n21817 = ~n9241 ;
  assign n9242 = n9236 & n21817 ;
  assign n9243 = n9235 | n9242 ;
  assign n9244 = x86 & n9243 ;
  assign n9245 = x86 | n9243 ;
  assign n9246 = n8835 & n21666 ;
  assign n9247 = n148 & n9246 ;
  assign n21818 = ~n8841 ;
  assign n9248 = n21818 & n9247 ;
  assign n21819 = ~n9247 ;
  assign n9249 = n8841 & n21819 ;
  assign n9250 = n9248 | n9249 ;
  assign n21820 = ~n9250 ;
  assign n9251 = n9245 & n21820 ;
  assign n9252 = n9244 | n9251 ;
  assign n9253 = x87 & n9252 ;
  assign n9254 = x87 | n9252 ;
  assign n9255 = n8844 & n21670 ;
  assign n9256 = n148 & n9255 ;
  assign n21821 = ~n8850 ;
  assign n9257 = n21821 & n9256 ;
  assign n21822 = ~n9256 ;
  assign n9258 = n8850 & n21822 ;
  assign n9259 = n9257 | n9258 ;
  assign n21823 = ~n9259 ;
  assign n9260 = n9254 & n21823 ;
  assign n9261 = n9253 | n9260 ;
  assign n9262 = x88 & n9261 ;
  assign n9263 = x88 | n9261 ;
  assign n9264 = n8853 & n21674 ;
  assign n9265 = n148 & n9264 ;
  assign n21824 = ~n8859 ;
  assign n9266 = n21824 & n9265 ;
  assign n21825 = ~n9265 ;
  assign n9267 = n8859 & n21825 ;
  assign n9268 = n9266 | n9267 ;
  assign n21826 = ~n9268 ;
  assign n9269 = n9263 & n21826 ;
  assign n9270 = n9262 | n9269 ;
  assign n9271 = x89 & n9270 ;
  assign n9272 = x89 | n9270 ;
  assign n9273 = n8862 & n21678 ;
  assign n9274 = n148 & n9273 ;
  assign n9275 = n8868 & n9274 ;
  assign n9276 = n8868 | n9274 ;
  assign n21827 = ~n9275 ;
  assign n9277 = n21827 & n9276 ;
  assign n21828 = ~n9277 ;
  assign n9278 = n9272 & n21828 ;
  assign n9279 = n9271 | n9278 ;
  assign n9280 = x90 & n9279 ;
  assign n9281 = x90 | n9279 ;
  assign n9282 = n8871 & n21682 ;
  assign n9283 = n148 & n9282 ;
  assign n9284 = n8877 & n9283 ;
  assign n9285 = n8877 | n9283 ;
  assign n21829 = ~n9284 ;
  assign n9286 = n21829 & n9285 ;
  assign n21830 = ~n9286 ;
  assign n9287 = n9281 & n21830 ;
  assign n9288 = n9280 | n9287 ;
  assign n9289 = x91 & n9288 ;
  assign n9290 = x91 | n9288 ;
  assign n9291 = n8880 & n21686 ;
  assign n9292 = n148 & n9291 ;
  assign n9293 = n8886 & n9292 ;
  assign n9294 = n8886 | n9292 ;
  assign n21831 = ~n9293 ;
  assign n9295 = n21831 & n9294 ;
  assign n21832 = ~n9295 ;
  assign n9296 = n9290 & n21832 ;
  assign n9297 = n9289 | n9296 ;
  assign n9298 = x92 & n9297 ;
  assign n9299 = x92 | n9297 ;
  assign n9300 = n8889 & n21690 ;
  assign n9301 = n148 & n9300 ;
  assign n21833 = ~n8895 ;
  assign n9302 = n21833 & n9301 ;
  assign n21834 = ~n9301 ;
  assign n9303 = n8895 & n21834 ;
  assign n9304 = n9302 | n9303 ;
  assign n21835 = ~n9304 ;
  assign n9305 = n9299 & n21835 ;
  assign n9306 = n9298 | n9305 ;
  assign n9307 = x93 & n9306 ;
  assign n9308 = x93 | n9306 ;
  assign n9309 = n8898 & n21694 ;
  assign n9310 = n148 & n9309 ;
  assign n21836 = ~n8904 ;
  assign n9311 = n21836 & n9310 ;
  assign n21837 = ~n9310 ;
  assign n9312 = n8904 & n21837 ;
  assign n9313 = n9311 | n9312 ;
  assign n21838 = ~n9313 ;
  assign n9314 = n9308 & n21838 ;
  assign n9315 = n9307 | n9314 ;
  assign n9316 = x94 & n9315 ;
  assign n9317 = x94 | n9315 ;
  assign n9318 = n8907 & n21698 ;
  assign n9319 = n148 & n9318 ;
  assign n21839 = ~n8913 ;
  assign n9320 = n21839 & n9319 ;
  assign n21840 = ~n9319 ;
  assign n9321 = n8913 & n21840 ;
  assign n9322 = n9320 | n9321 ;
  assign n21841 = ~n9322 ;
  assign n9323 = n9317 & n21841 ;
  assign n9324 = n9316 | n9323 ;
  assign n9325 = x95 & n9324 ;
  assign n9326 = x95 | n9324 ;
  assign n9327 = n8916 & n21702 ;
  assign n9328 = n148 & n9327 ;
  assign n21842 = ~n8922 ;
  assign n9329 = n21842 & n9328 ;
  assign n21843 = ~n9328 ;
  assign n9330 = n8922 & n21843 ;
  assign n9331 = n9329 | n9330 ;
  assign n21844 = ~n9331 ;
  assign n9332 = n9326 & n21844 ;
  assign n9333 = n9325 | n9332 ;
  assign n9334 = x96 & n9333 ;
  assign n9335 = x96 | n9333 ;
  assign n9336 = n8925 & n21706 ;
  assign n9337 = n148 & n9336 ;
  assign n21845 = ~n8931 ;
  assign n9338 = n21845 & n9337 ;
  assign n21846 = ~n9337 ;
  assign n9339 = n8931 & n21846 ;
  assign n9340 = n9338 | n9339 ;
  assign n21847 = ~n9340 ;
  assign n9341 = n9335 & n21847 ;
  assign n9342 = n9334 | n9341 ;
  assign n9343 = x97 & n9342 ;
  assign n9344 = x97 | n9342 ;
  assign n9345 = n8934 & n21710 ;
  assign n9346 = n148 & n9345 ;
  assign n21848 = ~n8940 ;
  assign n9347 = n21848 & n9346 ;
  assign n21849 = ~n9346 ;
  assign n9348 = n8940 & n21849 ;
  assign n9349 = n9347 | n9348 ;
  assign n21850 = ~n9349 ;
  assign n9350 = n9344 & n21850 ;
  assign n9351 = n9343 | n9350 ;
  assign n9352 = x98 & n9351 ;
  assign n9353 = x98 | n9351 ;
  assign n9354 = n8943 & n21714 ;
  assign n9355 = n148 & n9354 ;
  assign n21851 = ~n8949 ;
  assign n9356 = n21851 & n9355 ;
  assign n21852 = ~n9355 ;
  assign n9357 = n8949 & n21852 ;
  assign n9358 = n9356 | n9357 ;
  assign n21853 = ~n9358 ;
  assign n9359 = n9353 & n21853 ;
  assign n9360 = n9352 | n9359 ;
  assign n9361 = x99 & n9360 ;
  assign n9362 = x99 | n9360 ;
  assign n9363 = n8952 & n21718 ;
  assign n9364 = n148 & n9363 ;
  assign n21854 = ~n8958 ;
  assign n9365 = n21854 & n9364 ;
  assign n21855 = ~n9364 ;
  assign n9366 = n8958 & n21855 ;
  assign n9367 = n9365 | n9366 ;
  assign n21856 = ~n9367 ;
  assign n9368 = n9362 & n21856 ;
  assign n9369 = n9361 | n9368 ;
  assign n9370 = x100 & n9369 ;
  assign n9371 = x100 | n9369 ;
  assign n9372 = n8961 & n21722 ;
  assign n9373 = n148 & n9372 ;
  assign n21857 = ~n8967 ;
  assign n9374 = n21857 & n9373 ;
  assign n21858 = ~n9373 ;
  assign n9375 = n8967 & n21858 ;
  assign n9376 = n9374 | n9375 ;
  assign n21859 = ~n9376 ;
  assign n9377 = n9371 & n21859 ;
  assign n9378 = n9370 | n9377 ;
  assign n9379 = x101 & n9378 ;
  assign n9380 = x101 | n9378 ;
  assign n9381 = n8970 & n21726 ;
  assign n9382 = n148 & n9381 ;
  assign n21860 = ~n8976 ;
  assign n9383 = n21860 & n9382 ;
  assign n21861 = ~n9382 ;
  assign n9384 = n8976 & n21861 ;
  assign n9385 = n9383 | n9384 ;
  assign n21862 = ~n9385 ;
  assign n9386 = n9380 & n21862 ;
  assign n9387 = n9379 | n9386 ;
  assign n9388 = x102 & n9387 ;
  assign n9389 = x102 | n9387 ;
  assign n9390 = n8979 & n21730 ;
  assign n9391 = n148 & n9390 ;
  assign n21863 = ~n8985 ;
  assign n9392 = n21863 & n9391 ;
  assign n21864 = ~n9391 ;
  assign n9393 = n8985 & n21864 ;
  assign n9394 = n9392 | n9393 ;
  assign n21865 = ~n9394 ;
  assign n9395 = n9389 & n21865 ;
  assign n9396 = n9388 | n9395 ;
  assign n9397 = x103 & n9396 ;
  assign n9398 = x103 | n9396 ;
  assign n9399 = n8988 & n21734 ;
  assign n9400 = n148 & n9399 ;
  assign n21866 = ~n8994 ;
  assign n9401 = n21866 & n9400 ;
  assign n21867 = ~n9400 ;
  assign n9402 = n8994 & n21867 ;
  assign n9403 = n9401 | n9402 ;
  assign n21868 = ~n9403 ;
  assign n9404 = n9398 & n21868 ;
  assign n9405 = n9397 | n9404 ;
  assign n9406 = x104 & n9405 ;
  assign n9407 = x104 | n9405 ;
  assign n9408 = n8997 & n21738 ;
  assign n9409 = n148 & n9408 ;
  assign n21869 = ~n9003 ;
  assign n9410 = n21869 & n9409 ;
  assign n21870 = ~n9409 ;
  assign n9411 = n9003 & n21870 ;
  assign n9412 = n9410 | n9411 ;
  assign n21871 = ~n9412 ;
  assign n9413 = n9407 & n21871 ;
  assign n9414 = n9406 | n9413 ;
  assign n9415 = x105 & n9414 ;
  assign n9416 = x105 | n9414 ;
  assign n9417 = n9006 & n21742 ;
  assign n9418 = n148 & n9417 ;
  assign n21872 = ~n9012 ;
  assign n9419 = n21872 & n9418 ;
  assign n21873 = ~n9418 ;
  assign n9420 = n9012 & n21873 ;
  assign n9421 = n9419 | n9420 ;
  assign n21874 = ~n9421 ;
  assign n9422 = n9416 & n21874 ;
  assign n9423 = n9415 | n9422 ;
  assign n9424 = x106 & n9423 ;
  assign n9425 = x106 | n9423 ;
  assign n9426 = n9015 & n21746 ;
  assign n9427 = n148 & n9426 ;
  assign n21875 = ~n9021 ;
  assign n9428 = n21875 & n9427 ;
  assign n21876 = ~n9427 ;
  assign n9429 = n9021 & n21876 ;
  assign n9430 = n9428 | n9429 ;
  assign n21877 = ~n9430 ;
  assign n9431 = n9425 & n21877 ;
  assign n9432 = n9424 | n9431 ;
  assign n9433 = x107 & n9432 ;
  assign n9434 = x107 | n9432 ;
  assign n9435 = n9024 & n21750 ;
  assign n9436 = n148 & n9435 ;
  assign n21878 = ~n9030 ;
  assign n9437 = n21878 & n9436 ;
  assign n21879 = ~n9436 ;
  assign n9438 = n9030 & n21879 ;
  assign n9439 = n9437 | n9438 ;
  assign n21880 = ~n9439 ;
  assign n9440 = n9434 & n21880 ;
  assign n9441 = n9433 | n9440 ;
  assign n9442 = x108 & n9441 ;
  assign n9443 = x108 | n9441 ;
  assign n21881 = ~n9053 ;
  assign n9444 = n21881 & n9443 ;
  assign n9445 = n9442 | n9444 ;
  assign n21882 = ~n9057 ;
  assign n9446 = n21882 & n9445 ;
  assign n9447 = n18348 | n9446 ;
  assign n9448 = n9055 | n9447 ;
  assign n21883 = ~n9442 ;
  assign n9449 = n21883 & n9443 ;
  assign n147 = ~n9448 ;
  assign n9450 = n147 & n9449 ;
  assign n9451 = n21881 & n9450 ;
  assign n21885 = ~n9450 ;
  assign n9452 = n9053 & n21885 ;
  assign n9453 = n9451 | n9452 ;
  assign n21886 = ~x110 ;
  assign n9455 = n21886 & n9054 ;
  assign n9454 = x109 | n9445 ;
  assign n21887 = ~n9447 ;
  assign n9456 = n21887 & n9454 ;
  assign n21888 = ~n9456 ;
  assign n9457 = n9455 & n21888 ;
  assign n9056 = x110 & n21758 ;
  assign n21889 = ~x17 ;
  assign n9458 = n21889 & x64 ;
  assign n9460 = x65 | n9458 ;
  assign n9459 = x65 & n9458 ;
  assign n9461 = x64 & n147 ;
  assign n9462 = x18 & n9461 ;
  assign n9463 = x18 | n9461 ;
  assign n21890 = ~n9462 ;
  assign n9464 = n21890 & n9463 ;
  assign n21891 = ~n9459 ;
  assign n9465 = n21891 & n9464 ;
  assign n21892 = ~n9465 ;
  assign n9466 = n9460 & n21892 ;
  assign n9467 = x66 & n9466 ;
  assign n9468 = x66 | n9466 ;
  assign n9469 = n21762 & n9060 ;
  assign n9470 = n147 & n9469 ;
  assign n9471 = n9064 & n9470 ;
  assign n9472 = n9064 | n9470 ;
  assign n21893 = ~n9471 ;
  assign n9473 = n21893 & n9472 ;
  assign n21894 = ~n9473 ;
  assign n9474 = n9468 & n21894 ;
  assign n9475 = n9467 | n9474 ;
  assign n9476 = x67 & n9475 ;
  assign n9477 = x67 | n9475 ;
  assign n9478 = n9067 & n21765 ;
  assign n9479 = n147 & n9478 ;
  assign n21895 = ~n9072 ;
  assign n9480 = n21895 & n9479 ;
  assign n21896 = ~n9479 ;
  assign n9481 = n9072 & n21896 ;
  assign n9482 = n9480 | n9481 ;
  assign n21897 = ~n9482 ;
  assign n9483 = n9477 & n21897 ;
  assign n9484 = n9476 | n9483 ;
  assign n9485 = x68 & n9484 ;
  assign n9486 = x68 | n9484 ;
  assign n9487 = n9076 | n9448 ;
  assign n21898 = ~n9487 ;
  assign n9488 = n9080 & n21898 ;
  assign n9489 = n9075 & n21898 ;
  assign n21899 = ~n9489 ;
  assign n9490 = n9079 & n21899 ;
  assign n9491 = n9488 | n9490 ;
  assign n21900 = ~n9491 ;
  assign n9492 = n9486 & n21900 ;
  assign n9493 = n9485 | n9492 ;
  assign n9494 = x69 & n9493 ;
  assign n9495 = x69 | n9493 ;
  assign n21901 = ~n9082 ;
  assign n9496 = n21901 & n9083 ;
  assign n9497 = n147 & n9496 ;
  assign n9498 = n9088 & n9497 ;
  assign n9499 = n9088 | n9497 ;
  assign n21902 = ~n9498 ;
  assign n9500 = n21902 & n9499 ;
  assign n21903 = ~n9500 ;
  assign n9501 = n9495 & n21903 ;
  assign n9502 = n9494 | n9501 ;
  assign n9503 = x70 & n9502 ;
  assign n9504 = x70 | n9502 ;
  assign n21904 = ~n9091 ;
  assign n9505 = n21904 & n9092 ;
  assign n9506 = n147 & n9505 ;
  assign n9507 = n9097 & n9506 ;
  assign n9508 = n9097 | n9506 ;
  assign n21905 = ~n9507 ;
  assign n9509 = n21905 & n9508 ;
  assign n21906 = ~n9509 ;
  assign n9510 = n9504 & n21906 ;
  assign n9511 = n9503 | n9510 ;
  assign n9512 = x71 & n9511 ;
  assign n9513 = x71 | n9511 ;
  assign n21907 = ~n9100 ;
  assign n9514 = n21907 & n9101 ;
  assign n9515 = n147 & n9514 ;
  assign n9516 = n9106 & n9515 ;
  assign n9517 = n9106 | n9515 ;
  assign n21908 = ~n9516 ;
  assign n9518 = n21908 & n9517 ;
  assign n21909 = ~n9518 ;
  assign n9519 = n9513 & n21909 ;
  assign n9520 = n9512 | n9519 ;
  assign n9521 = x72 & n9520 ;
  assign n9522 = x72 | n9520 ;
  assign n21910 = ~n9109 ;
  assign n9523 = n21910 & n9110 ;
  assign n9524 = n147 & n9523 ;
  assign n9525 = n21778 & n9524 ;
  assign n21911 = ~n9524 ;
  assign n9526 = n9115 & n21911 ;
  assign n9527 = n9525 | n9526 ;
  assign n21912 = ~n9527 ;
  assign n9528 = n9522 & n21912 ;
  assign n9529 = n9521 | n9528 ;
  assign n9530 = x73 & n9529 ;
  assign n9531 = x73 | n9529 ;
  assign n21913 = ~n9118 ;
  assign n9532 = n21913 & n9119 ;
  assign n9533 = n147 & n9532 ;
  assign n9534 = n21781 & n9533 ;
  assign n21914 = ~n9533 ;
  assign n9535 = n9124 & n21914 ;
  assign n9536 = n9534 | n9535 ;
  assign n21915 = ~n9536 ;
  assign n9537 = n9531 & n21915 ;
  assign n9538 = n9530 | n9537 ;
  assign n9539 = x74 & n9538 ;
  assign n9540 = x74 | n9538 ;
  assign n21916 = ~n9127 ;
  assign n9541 = n21916 & n9128 ;
  assign n9542 = n147 & n9541 ;
  assign n9543 = n9133 & n9542 ;
  assign n9544 = n9133 | n9542 ;
  assign n21917 = ~n9543 ;
  assign n9545 = n21917 & n9544 ;
  assign n21918 = ~n9545 ;
  assign n9546 = n9540 & n21918 ;
  assign n9547 = n9539 | n9546 ;
  assign n9548 = x75 & n9547 ;
  assign n9549 = x75 | n9547 ;
  assign n21919 = ~n9136 ;
  assign n9550 = n21919 & n9137 ;
  assign n9551 = n147 & n9550 ;
  assign n9552 = n21786 & n9551 ;
  assign n21920 = ~n9551 ;
  assign n9553 = n9142 & n21920 ;
  assign n9554 = n9552 | n9553 ;
  assign n21921 = ~n9554 ;
  assign n9555 = n9549 & n21921 ;
  assign n9556 = n9548 | n9555 ;
  assign n9557 = x76 & n9556 ;
  assign n9558 = x76 | n9556 ;
  assign n21922 = ~n9145 ;
  assign n9559 = n21922 & n9146 ;
  assign n9560 = n147 & n9559 ;
  assign n9561 = n9151 & n9560 ;
  assign n9562 = n9151 | n9560 ;
  assign n21923 = ~n9561 ;
  assign n9563 = n21923 & n9562 ;
  assign n21924 = ~n9563 ;
  assign n9564 = n9558 & n21924 ;
  assign n9565 = n9557 | n9564 ;
  assign n9566 = x77 & n9565 ;
  assign n9567 = x77 | n9565 ;
  assign n21925 = ~n9154 ;
  assign n9568 = n21925 & n9155 ;
  assign n9569 = n147 & n9568 ;
  assign n9570 = n9160 & n9569 ;
  assign n9571 = n9160 | n9569 ;
  assign n21926 = ~n9570 ;
  assign n9572 = n21926 & n9571 ;
  assign n21927 = ~n9572 ;
  assign n9573 = n9567 & n21927 ;
  assign n9574 = n9566 | n9573 ;
  assign n9575 = x78 & n9574 ;
  assign n9576 = x78 | n9574 ;
  assign n21928 = ~n9163 ;
  assign n9577 = n21928 & n9164 ;
  assign n9578 = n147 & n9577 ;
  assign n9579 = n9169 & n9578 ;
  assign n9580 = n9169 | n9578 ;
  assign n21929 = ~n9579 ;
  assign n9581 = n21929 & n9580 ;
  assign n21930 = ~n9581 ;
  assign n9582 = n9576 & n21930 ;
  assign n9583 = n9575 | n9582 ;
  assign n9584 = x79 & n9583 ;
  assign n9585 = x79 | n9583 ;
  assign n21931 = ~n9172 ;
  assign n9586 = n21931 & n9173 ;
  assign n9587 = n147 & n9586 ;
  assign n9588 = n21796 & n9587 ;
  assign n21932 = ~n9587 ;
  assign n9589 = n9178 & n21932 ;
  assign n9590 = n9588 | n9589 ;
  assign n21933 = ~n9590 ;
  assign n9591 = n9585 & n21933 ;
  assign n9592 = n9584 | n9591 ;
  assign n9593 = x80 & n9592 ;
  assign n9594 = x80 | n9592 ;
  assign n21934 = ~n9181 ;
  assign n9595 = n21934 & n9182 ;
  assign n9596 = n147 & n9595 ;
  assign n9597 = n21799 & n9596 ;
  assign n21935 = ~n9596 ;
  assign n9598 = n9187 & n21935 ;
  assign n9599 = n9597 | n9598 ;
  assign n21936 = ~n9599 ;
  assign n9600 = n9594 & n21936 ;
  assign n9601 = n9593 | n9600 ;
  assign n9602 = x81 & n9601 ;
  assign n9603 = x81 | n9601 ;
  assign n21937 = ~n9190 ;
  assign n9604 = n21937 & n9191 ;
  assign n9605 = n147 & n9604 ;
  assign n9606 = n9196 & n9605 ;
  assign n9607 = n9196 | n9605 ;
  assign n21938 = ~n9606 ;
  assign n9608 = n21938 & n9607 ;
  assign n21939 = ~n9608 ;
  assign n9609 = n9603 & n21939 ;
  assign n9610 = n9602 | n9609 ;
  assign n9611 = x82 & n9610 ;
  assign n9612 = x82 | n9610 ;
  assign n21940 = ~n9199 ;
  assign n9613 = n21940 & n9200 ;
  assign n9614 = n147 & n9613 ;
  assign n9615 = n9205 & n9614 ;
  assign n9616 = n9205 | n9614 ;
  assign n21941 = ~n9615 ;
  assign n9617 = n21941 & n9616 ;
  assign n21942 = ~n9617 ;
  assign n9618 = n9612 & n21942 ;
  assign n9619 = n9611 | n9618 ;
  assign n9620 = x83 & n9619 ;
  assign n9621 = x83 | n9619 ;
  assign n21943 = ~n9208 ;
  assign n9622 = n21943 & n9209 ;
  assign n9623 = n147 & n9622 ;
  assign n9624 = n21808 & n9623 ;
  assign n21944 = ~n9623 ;
  assign n9625 = n9214 & n21944 ;
  assign n9626 = n9624 | n9625 ;
  assign n21945 = ~n9626 ;
  assign n9627 = n9621 & n21945 ;
  assign n9628 = n9620 | n9627 ;
  assign n9629 = x84 & n9628 ;
  assign n9630 = x84 | n9628 ;
  assign n21946 = ~n9217 ;
  assign n9631 = n21946 & n9218 ;
  assign n9632 = n147 & n9631 ;
  assign n9633 = n21811 & n9632 ;
  assign n21947 = ~n9632 ;
  assign n9634 = n9223 & n21947 ;
  assign n9635 = n9633 | n9634 ;
  assign n21948 = ~n9635 ;
  assign n9636 = n9630 & n21948 ;
  assign n9637 = n9629 | n9636 ;
  assign n9638 = x85 & n9637 ;
  assign n9639 = x85 | n9637 ;
  assign n21949 = ~n9226 ;
  assign n9640 = n21949 & n9227 ;
  assign n9641 = n147 & n9640 ;
  assign n9642 = n21814 & n9641 ;
  assign n21950 = ~n9641 ;
  assign n9643 = n9232 & n21950 ;
  assign n9644 = n9642 | n9643 ;
  assign n21951 = ~n9644 ;
  assign n9645 = n9639 & n21951 ;
  assign n9646 = n9638 | n9645 ;
  assign n9647 = x86 & n9646 ;
  assign n9648 = x86 | n9646 ;
  assign n21952 = ~n9235 ;
  assign n9649 = n21952 & n9236 ;
  assign n9650 = n147 & n9649 ;
  assign n9651 = n21817 & n9650 ;
  assign n21953 = ~n9650 ;
  assign n9652 = n9241 & n21953 ;
  assign n9653 = n9651 | n9652 ;
  assign n21954 = ~n9653 ;
  assign n9654 = n9648 & n21954 ;
  assign n9655 = n9647 | n9654 ;
  assign n9656 = x87 & n9655 ;
  assign n9657 = x87 | n9655 ;
  assign n21955 = ~n9244 ;
  assign n9658 = n21955 & n9245 ;
  assign n9659 = n147 & n9658 ;
  assign n9660 = n9250 & n9659 ;
  assign n9661 = n9250 | n9659 ;
  assign n21956 = ~n9660 ;
  assign n9662 = n21956 & n9661 ;
  assign n21957 = ~n9662 ;
  assign n9663 = n9657 & n21957 ;
  assign n9664 = n9656 | n9663 ;
  assign n9665 = x88 & n9664 ;
  assign n9666 = x88 | n9664 ;
  assign n21958 = ~n9253 ;
  assign n9667 = n21958 & n9254 ;
  assign n9668 = n147 & n9667 ;
  assign n9669 = n21823 & n9668 ;
  assign n21959 = ~n9668 ;
  assign n9670 = n9259 & n21959 ;
  assign n9671 = n9669 | n9670 ;
  assign n21960 = ~n9671 ;
  assign n9672 = n9666 & n21960 ;
  assign n9673 = n9665 | n9672 ;
  assign n9674 = x89 & n9673 ;
  assign n9675 = x89 | n9673 ;
  assign n21961 = ~n9262 ;
  assign n9676 = n21961 & n9263 ;
  assign n9677 = n147 & n9676 ;
  assign n9678 = n21826 & n9677 ;
  assign n21962 = ~n9677 ;
  assign n9679 = n9268 & n21962 ;
  assign n9680 = n9678 | n9679 ;
  assign n21963 = ~n9680 ;
  assign n9681 = n9675 & n21963 ;
  assign n9682 = n9674 | n9681 ;
  assign n9683 = x90 & n9682 ;
  assign n9684 = x90 | n9682 ;
  assign n21964 = ~n9271 ;
  assign n9685 = n21964 & n9272 ;
  assign n9686 = n147 & n9685 ;
  assign n9687 = n9277 & n9686 ;
  assign n9688 = n9277 | n9686 ;
  assign n21965 = ~n9687 ;
  assign n9689 = n21965 & n9688 ;
  assign n21966 = ~n9689 ;
  assign n9690 = n9684 & n21966 ;
  assign n9691 = n9683 | n9690 ;
  assign n9692 = x91 & n9691 ;
  assign n9693 = x91 | n9691 ;
  assign n21967 = ~n9280 ;
  assign n9694 = n21967 & n9281 ;
  assign n9695 = n147 & n9694 ;
  assign n9696 = n9286 & n9695 ;
  assign n9697 = n9286 | n9695 ;
  assign n21968 = ~n9696 ;
  assign n9698 = n21968 & n9697 ;
  assign n21969 = ~n9698 ;
  assign n9699 = n9693 & n21969 ;
  assign n9700 = n9692 | n9699 ;
  assign n9701 = x92 & n9700 ;
  assign n9702 = x92 | n9700 ;
  assign n21970 = ~n9289 ;
  assign n9703 = n21970 & n9290 ;
  assign n9704 = n147 & n9703 ;
  assign n9705 = n9295 & n9704 ;
  assign n9706 = n9295 | n9704 ;
  assign n21971 = ~n9705 ;
  assign n9707 = n21971 & n9706 ;
  assign n21972 = ~n9707 ;
  assign n9708 = n9702 & n21972 ;
  assign n9709 = n9701 | n9708 ;
  assign n9710 = x93 & n9709 ;
  assign n9711 = x93 | n9709 ;
  assign n21973 = ~n9298 ;
  assign n9712 = n21973 & n9299 ;
  assign n9713 = n147 & n9712 ;
  assign n9714 = n21835 & n9713 ;
  assign n21974 = ~n9713 ;
  assign n9715 = n9304 & n21974 ;
  assign n9716 = n9714 | n9715 ;
  assign n21975 = ~n9716 ;
  assign n9717 = n9711 & n21975 ;
  assign n9718 = n9710 | n9717 ;
  assign n9719 = x94 & n9718 ;
  assign n9720 = x94 | n9718 ;
  assign n21976 = ~n9307 ;
  assign n9721 = n21976 & n9308 ;
  assign n9722 = n147 & n9721 ;
  assign n9723 = n21838 & n9722 ;
  assign n21977 = ~n9722 ;
  assign n9724 = n9313 & n21977 ;
  assign n9725 = n9723 | n9724 ;
  assign n21978 = ~n9725 ;
  assign n9726 = n9720 & n21978 ;
  assign n9727 = n9719 | n9726 ;
  assign n9728 = x95 & n9727 ;
  assign n9729 = x95 | n9727 ;
  assign n21979 = ~n9316 ;
  assign n9730 = n21979 & n9317 ;
  assign n9731 = n147 & n9730 ;
  assign n9732 = n9322 & n9731 ;
  assign n9733 = n9322 | n9731 ;
  assign n21980 = ~n9732 ;
  assign n9734 = n21980 & n9733 ;
  assign n21981 = ~n9734 ;
  assign n9735 = n9729 & n21981 ;
  assign n9736 = n9728 | n9735 ;
  assign n9737 = x96 & n9736 ;
  assign n9738 = x96 | n9736 ;
  assign n21982 = ~n9325 ;
  assign n9739 = n21982 & n9326 ;
  assign n9740 = n147 & n9739 ;
  assign n9741 = n21844 & n9740 ;
  assign n21983 = ~n9740 ;
  assign n9742 = n9331 & n21983 ;
  assign n9743 = n9741 | n9742 ;
  assign n21984 = ~n9743 ;
  assign n9744 = n9738 & n21984 ;
  assign n9745 = n9737 | n9744 ;
  assign n9746 = x97 & n9745 ;
  assign n9747 = x97 | n9745 ;
  assign n21985 = ~n9334 ;
  assign n9748 = n21985 & n9335 ;
  assign n9749 = n147 & n9748 ;
  assign n9750 = n21847 & n9749 ;
  assign n21986 = ~n9749 ;
  assign n9751 = n9340 & n21986 ;
  assign n9752 = n9750 | n9751 ;
  assign n21987 = ~n9752 ;
  assign n9753 = n9747 & n21987 ;
  assign n9754 = n9746 | n9753 ;
  assign n9755 = x98 & n9754 ;
  assign n9756 = x98 | n9754 ;
  assign n21988 = ~n9343 ;
  assign n9757 = n21988 & n9344 ;
  assign n9758 = n147 & n9757 ;
  assign n9759 = n9349 & n9758 ;
  assign n9760 = n9349 | n9758 ;
  assign n21989 = ~n9759 ;
  assign n9761 = n21989 & n9760 ;
  assign n21990 = ~n9761 ;
  assign n9762 = n9756 & n21990 ;
  assign n9763 = n9755 | n9762 ;
  assign n9764 = x99 & n9763 ;
  assign n9765 = x99 | n9763 ;
  assign n21991 = ~n9352 ;
  assign n9766 = n21991 & n9353 ;
  assign n9767 = n147 & n9766 ;
  assign n9768 = n9358 & n9767 ;
  assign n9769 = n9358 | n9767 ;
  assign n21992 = ~n9768 ;
  assign n9770 = n21992 & n9769 ;
  assign n21993 = ~n9770 ;
  assign n9771 = n9765 & n21993 ;
  assign n9772 = n9764 | n9771 ;
  assign n9773 = x100 & n9772 ;
  assign n9774 = x100 | n9772 ;
  assign n21994 = ~n9361 ;
  assign n9775 = n21994 & n9362 ;
  assign n9776 = n147 & n9775 ;
  assign n9777 = n9367 & n9776 ;
  assign n9778 = n9367 | n9776 ;
  assign n21995 = ~n9777 ;
  assign n9779 = n21995 & n9778 ;
  assign n21996 = ~n9779 ;
  assign n9780 = n9774 & n21996 ;
  assign n9781 = n9773 | n9780 ;
  assign n9782 = x101 & n9781 ;
  assign n9783 = x101 | n9781 ;
  assign n21997 = ~n9370 ;
  assign n9784 = n21997 & n9371 ;
  assign n9785 = n147 & n9784 ;
  assign n9786 = n21859 & n9785 ;
  assign n21998 = ~n9785 ;
  assign n9787 = n9376 & n21998 ;
  assign n9788 = n9786 | n9787 ;
  assign n21999 = ~n9788 ;
  assign n9789 = n9783 & n21999 ;
  assign n9790 = n9782 | n9789 ;
  assign n9791 = x102 & n9790 ;
  assign n9792 = x102 | n9790 ;
  assign n22000 = ~n9379 ;
  assign n9793 = n22000 & n9380 ;
  assign n9794 = n147 & n9793 ;
  assign n9795 = n21862 & n9794 ;
  assign n22001 = ~n9794 ;
  assign n9796 = n9385 & n22001 ;
  assign n9797 = n9795 | n9796 ;
  assign n22002 = ~n9797 ;
  assign n9798 = n9792 & n22002 ;
  assign n9799 = n9791 | n9798 ;
  assign n9800 = x103 & n9799 ;
  assign n9801 = x103 | n9799 ;
  assign n22003 = ~n9388 ;
  assign n9802 = n22003 & n9389 ;
  assign n9803 = n147 & n9802 ;
  assign n9804 = n21865 & n9803 ;
  assign n22004 = ~n9803 ;
  assign n9805 = n9394 & n22004 ;
  assign n9806 = n9804 | n9805 ;
  assign n22005 = ~n9806 ;
  assign n9807 = n9801 & n22005 ;
  assign n9808 = n9800 | n9807 ;
  assign n9809 = x104 & n9808 ;
  assign n9810 = x104 | n9808 ;
  assign n22006 = ~n9397 ;
  assign n9811 = n22006 & n9398 ;
  assign n9812 = n147 & n9811 ;
  assign n9813 = n9403 & n9812 ;
  assign n9814 = n9403 | n9812 ;
  assign n22007 = ~n9813 ;
  assign n9815 = n22007 & n9814 ;
  assign n22008 = ~n9815 ;
  assign n9816 = n9810 & n22008 ;
  assign n9817 = n9809 | n9816 ;
  assign n9818 = x105 & n9817 ;
  assign n9819 = x105 | n9817 ;
  assign n22009 = ~n9406 ;
  assign n9820 = n22009 & n9407 ;
  assign n9821 = n147 & n9820 ;
  assign n9822 = n9412 & n9821 ;
  assign n9823 = n9412 | n9821 ;
  assign n22010 = ~n9822 ;
  assign n9824 = n22010 & n9823 ;
  assign n22011 = ~n9824 ;
  assign n9825 = n9819 & n22011 ;
  assign n9826 = n9818 | n9825 ;
  assign n9827 = x106 & n9826 ;
  assign n9828 = x106 | n9826 ;
  assign n22012 = ~n9415 ;
  assign n9829 = n22012 & n9416 ;
  assign n9830 = n147 & n9829 ;
  assign n9831 = n9421 & n9830 ;
  assign n9832 = n9421 | n9830 ;
  assign n22013 = ~n9831 ;
  assign n9833 = n22013 & n9832 ;
  assign n22014 = ~n9833 ;
  assign n9834 = n9828 & n22014 ;
  assign n9835 = n9827 | n9834 ;
  assign n9836 = x107 & n9835 ;
  assign n9837 = x107 | n9835 ;
  assign n22015 = ~n9424 ;
  assign n9838 = n22015 & n9425 ;
  assign n9839 = n147 & n9838 ;
  assign n9840 = n21877 & n9839 ;
  assign n22016 = ~n9839 ;
  assign n9841 = n9430 & n22016 ;
  assign n9842 = n9840 | n9841 ;
  assign n22017 = ~n9842 ;
  assign n9843 = n9837 & n22017 ;
  assign n9844 = n9836 | n9843 ;
  assign n9845 = x108 & n9844 ;
  assign n9846 = x108 | n9844 ;
  assign n22018 = ~n9433 ;
  assign n9847 = n22018 & n9434 ;
  assign n9848 = n147 & n9847 ;
  assign n9849 = n9439 & n9848 ;
  assign n9850 = n9439 | n9848 ;
  assign n22019 = ~n9849 ;
  assign n9851 = n22019 & n9850 ;
  assign n22020 = ~n9851 ;
  assign n9852 = n9846 & n22020 ;
  assign n9853 = n9845 | n9852 ;
  assign n9854 = x109 & n9853 ;
  assign n9857 = n9056 | n9854 ;
  assign n9856 = x109 | n9853 ;
  assign n22021 = ~n9453 ;
  assign n9858 = n22021 & n9856 ;
  assign n9859 = n9857 | n9858 ;
  assign n22022 = ~n9457 ;
  assign n9860 = n22022 & n9859 ;
  assign n9861 = n18343 | n9860 ;
  assign n9855 = n21759 & n9853 ;
  assign n22023 = ~n9853 ;
  assign n9865 = x109 & n22023 ;
  assign n9866 = n9855 | n9865 ;
  assign n146 = ~n9861 ;
  assign n9867 = n146 & n9866 ;
  assign n9868 = n9453 & n9867 ;
  assign n9869 = n9453 | n9867 ;
  assign n22025 = ~n9868 ;
  assign n9870 = n22025 & n9869 ;
  assign n22026 = ~x16 ;
  assign n9871 = n22026 & x64 ;
  assign n9872 = x65 | n9871 ;
  assign n9873 = x65 & n9871 ;
  assign n9863 = n9458 & n146 ;
  assign n9862 = x64 & n146 ;
  assign n22027 = ~n9862 ;
  assign n9874 = x17 & n22027 ;
  assign n9875 = n9863 | n9874 ;
  assign n22028 = ~n9873 ;
  assign n9876 = n22028 & n9875 ;
  assign n22029 = ~n9876 ;
  assign n9877 = n9872 & n22029 ;
  assign n9880 = x66 & n9877 ;
  assign n9878 = x66 | n9877 ;
  assign n9881 = n21891 & n9460 ;
  assign n9882 = n146 & n9881 ;
  assign n9883 = n9464 & n9882 ;
  assign n9884 = n9464 | n9882 ;
  assign n22030 = ~n9883 ;
  assign n9885 = n22030 & n9884 ;
  assign n22031 = ~n9885 ;
  assign n9886 = n9878 & n22031 ;
  assign n9887 = n9880 | n9886 ;
  assign n9888 = x67 & n9887 ;
  assign n9889 = x67 | n9887 ;
  assign n22032 = ~n9467 ;
  assign n9890 = n22032 & n9468 ;
  assign n9891 = n146 & n9890 ;
  assign n9892 = n9473 & n9891 ;
  assign n9893 = n9473 | n9891 ;
  assign n22033 = ~n9892 ;
  assign n9894 = n22033 & n9893 ;
  assign n22034 = ~n9894 ;
  assign n9895 = n9889 & n22034 ;
  assign n9896 = n9888 | n9895 ;
  assign n9897 = x68 & n9896 ;
  assign n9898 = x68 | n9896 ;
  assign n22035 = ~n9476 ;
  assign n9899 = n22035 & n9477 ;
  assign n9900 = n146 & n9899 ;
  assign n9901 = n9482 & n9900 ;
  assign n9902 = n9482 | n9900 ;
  assign n22036 = ~n9901 ;
  assign n9903 = n22036 & n9902 ;
  assign n22037 = ~n9903 ;
  assign n9904 = n9898 & n22037 ;
  assign n9905 = n9897 | n9904 ;
  assign n9906 = x69 & n9905 ;
  assign n9907 = x69 | n9905 ;
  assign n22038 = ~n9485 ;
  assign n9908 = n22038 & n9486 ;
  assign n9909 = n146 & n9908 ;
  assign n9910 = n9491 & n9909 ;
  assign n9911 = n9491 | n9909 ;
  assign n22039 = ~n9910 ;
  assign n9912 = n22039 & n9911 ;
  assign n22040 = ~n9912 ;
  assign n9913 = n9907 & n22040 ;
  assign n9914 = n9906 | n9913 ;
  assign n9915 = x70 & n9914 ;
  assign n9916 = x70 | n9914 ;
  assign n22041 = ~n9494 ;
  assign n9917 = n22041 & n9495 ;
  assign n9918 = n146 & n9917 ;
  assign n9919 = n21903 & n9918 ;
  assign n22042 = ~n9918 ;
  assign n9920 = n9500 & n22042 ;
  assign n9921 = n9919 | n9920 ;
  assign n22043 = ~n9921 ;
  assign n9922 = n9916 & n22043 ;
  assign n9923 = n9915 | n9922 ;
  assign n9924 = x71 & n9923 ;
  assign n9925 = x71 | n9923 ;
  assign n22044 = ~n9503 ;
  assign n9926 = n22044 & n9504 ;
  assign n9927 = n146 & n9926 ;
  assign n9928 = n9509 & n9927 ;
  assign n9929 = n9509 | n9927 ;
  assign n22045 = ~n9928 ;
  assign n9930 = n22045 & n9929 ;
  assign n22046 = ~n9930 ;
  assign n9931 = n9925 & n22046 ;
  assign n9932 = n9924 | n9931 ;
  assign n9933 = x72 & n9932 ;
  assign n9934 = x72 | n9932 ;
  assign n22047 = ~n9512 ;
  assign n9935 = n22047 & n9513 ;
  assign n9936 = n146 & n9935 ;
  assign n9937 = n9518 & n9936 ;
  assign n9938 = n9518 | n9936 ;
  assign n22048 = ~n9937 ;
  assign n9939 = n22048 & n9938 ;
  assign n22049 = ~n9939 ;
  assign n9940 = n9934 & n22049 ;
  assign n9941 = n9933 | n9940 ;
  assign n9942 = x73 & n9941 ;
  assign n9943 = x73 | n9941 ;
  assign n22050 = ~n9521 ;
  assign n9944 = n22050 & n9522 ;
  assign n9945 = n146 & n9944 ;
  assign n9946 = n21912 & n9945 ;
  assign n22051 = ~n9945 ;
  assign n9947 = n9527 & n22051 ;
  assign n9948 = n9946 | n9947 ;
  assign n22052 = ~n9948 ;
  assign n9949 = n9943 & n22052 ;
  assign n9950 = n9942 | n9949 ;
  assign n9951 = x74 & n9950 ;
  assign n9952 = x74 | n9950 ;
  assign n22053 = ~n9530 ;
  assign n9953 = n22053 & n9531 ;
  assign n9954 = n146 & n9953 ;
  assign n9955 = n21915 & n9954 ;
  assign n22054 = ~n9954 ;
  assign n9956 = n9536 & n22054 ;
  assign n9957 = n9955 | n9956 ;
  assign n22055 = ~n9957 ;
  assign n9958 = n9952 & n22055 ;
  assign n9959 = n9951 | n9958 ;
  assign n9960 = x75 & n9959 ;
  assign n9961 = x75 | n9959 ;
  assign n22056 = ~n9539 ;
  assign n9962 = n22056 & n9540 ;
  assign n9963 = n146 & n9962 ;
  assign n9964 = n9545 & n9963 ;
  assign n9965 = n9545 | n9963 ;
  assign n22057 = ~n9964 ;
  assign n9966 = n22057 & n9965 ;
  assign n22058 = ~n9966 ;
  assign n9967 = n9961 & n22058 ;
  assign n9968 = n9960 | n9967 ;
  assign n9969 = x76 & n9968 ;
  assign n9970 = x76 | n9968 ;
  assign n22059 = ~n9548 ;
  assign n9971 = n22059 & n9549 ;
  assign n9972 = n146 & n9971 ;
  assign n9973 = n21921 & n9972 ;
  assign n22060 = ~n9972 ;
  assign n9974 = n9554 & n22060 ;
  assign n9975 = n9973 | n9974 ;
  assign n22061 = ~n9975 ;
  assign n9976 = n9970 & n22061 ;
  assign n9977 = n9969 | n9976 ;
  assign n9978 = x77 & n9977 ;
  assign n9979 = x77 | n9977 ;
  assign n22062 = ~n9557 ;
  assign n9980 = n22062 & n9558 ;
  assign n9981 = n146 & n9980 ;
  assign n9982 = n9563 & n9981 ;
  assign n9983 = n9563 | n9981 ;
  assign n22063 = ~n9982 ;
  assign n9984 = n22063 & n9983 ;
  assign n22064 = ~n9984 ;
  assign n9985 = n9979 & n22064 ;
  assign n9986 = n9978 | n9985 ;
  assign n9987 = x78 & n9986 ;
  assign n9988 = x78 | n9986 ;
  assign n22065 = ~n9566 ;
  assign n9989 = n22065 & n9567 ;
  assign n9990 = n146 & n9989 ;
  assign n9991 = n9572 & n9990 ;
  assign n9992 = n9572 | n9990 ;
  assign n22066 = ~n9991 ;
  assign n9993 = n22066 & n9992 ;
  assign n22067 = ~n9993 ;
  assign n9994 = n9988 & n22067 ;
  assign n9995 = n9987 | n9994 ;
  assign n9996 = x79 & n9995 ;
  assign n9997 = x79 | n9995 ;
  assign n22068 = ~n9575 ;
  assign n9998 = n22068 & n9576 ;
  assign n9999 = n146 & n9998 ;
  assign n10000 = n9581 & n9999 ;
  assign n10001 = n9581 | n9999 ;
  assign n22069 = ~n10000 ;
  assign n10002 = n22069 & n10001 ;
  assign n22070 = ~n10002 ;
  assign n10003 = n9997 & n22070 ;
  assign n10004 = n9996 | n10003 ;
  assign n10005 = x80 & n10004 ;
  assign n10006 = x80 | n10004 ;
  assign n22071 = ~n9584 ;
  assign n10007 = n22071 & n9585 ;
  assign n10008 = n146 & n10007 ;
  assign n10009 = n21933 & n10008 ;
  assign n22072 = ~n10008 ;
  assign n10010 = n9590 & n22072 ;
  assign n10011 = n10009 | n10010 ;
  assign n22073 = ~n10011 ;
  assign n10012 = n10006 & n22073 ;
  assign n10013 = n10005 | n10012 ;
  assign n10014 = x81 & n10013 ;
  assign n10015 = x81 | n10013 ;
  assign n22074 = ~n9593 ;
  assign n10016 = n22074 & n9594 ;
  assign n10017 = n146 & n10016 ;
  assign n10018 = n21936 & n10017 ;
  assign n22075 = ~n10017 ;
  assign n10019 = n9599 & n22075 ;
  assign n10020 = n10018 | n10019 ;
  assign n22076 = ~n10020 ;
  assign n10021 = n10015 & n22076 ;
  assign n10022 = n10014 | n10021 ;
  assign n10023 = x82 & n10022 ;
  assign n10024 = x82 | n10022 ;
  assign n22077 = ~n9602 ;
  assign n10025 = n22077 & n9603 ;
  assign n10026 = n146 & n10025 ;
  assign n10027 = n9608 & n10026 ;
  assign n10028 = n9608 | n10026 ;
  assign n22078 = ~n10027 ;
  assign n10029 = n22078 & n10028 ;
  assign n22079 = ~n10029 ;
  assign n10030 = n10024 & n22079 ;
  assign n10031 = n10023 | n10030 ;
  assign n10032 = x83 & n10031 ;
  assign n10033 = x83 | n10031 ;
  assign n22080 = ~n9611 ;
  assign n10034 = n22080 & n9612 ;
  assign n10035 = n146 & n10034 ;
  assign n10036 = n9617 & n10035 ;
  assign n10037 = n9617 | n10035 ;
  assign n22081 = ~n10036 ;
  assign n10038 = n22081 & n10037 ;
  assign n22082 = ~n10038 ;
  assign n10039 = n10033 & n22082 ;
  assign n10040 = n10032 | n10039 ;
  assign n10041 = x84 & n10040 ;
  assign n10042 = x84 | n10040 ;
  assign n22083 = ~n9620 ;
  assign n10043 = n22083 & n9621 ;
  assign n10044 = n146 & n10043 ;
  assign n10045 = n9626 & n10044 ;
  assign n10046 = n9626 | n10044 ;
  assign n22084 = ~n10045 ;
  assign n10047 = n22084 & n10046 ;
  assign n22085 = ~n10047 ;
  assign n10048 = n10042 & n22085 ;
  assign n10049 = n10041 | n10048 ;
  assign n10050 = x85 & n10049 ;
  assign n10051 = x85 | n10049 ;
  assign n22086 = ~n9629 ;
  assign n10052 = n22086 & n9630 ;
  assign n10053 = n146 & n10052 ;
  assign n10054 = n21948 & n10053 ;
  assign n22087 = ~n10053 ;
  assign n10055 = n9635 & n22087 ;
  assign n10056 = n10054 | n10055 ;
  assign n22088 = ~n10056 ;
  assign n10057 = n10051 & n22088 ;
  assign n10058 = n10050 | n10057 ;
  assign n10059 = x86 & n10058 ;
  assign n10060 = x86 | n10058 ;
  assign n22089 = ~n9638 ;
  assign n10061 = n22089 & n9639 ;
  assign n10062 = n146 & n10061 ;
  assign n10063 = n9644 & n10062 ;
  assign n10064 = n9644 | n10062 ;
  assign n22090 = ~n10063 ;
  assign n10065 = n22090 & n10064 ;
  assign n22091 = ~n10065 ;
  assign n10066 = n10060 & n22091 ;
  assign n10067 = n10059 | n10066 ;
  assign n10068 = x87 & n10067 ;
  assign n10069 = x87 | n10067 ;
  assign n22092 = ~n9647 ;
  assign n10070 = n22092 & n9648 ;
  assign n10071 = n146 & n10070 ;
  assign n10072 = n21954 & n10071 ;
  assign n22093 = ~n10071 ;
  assign n10073 = n9653 & n22093 ;
  assign n10074 = n10072 | n10073 ;
  assign n22094 = ~n10074 ;
  assign n10075 = n10069 & n22094 ;
  assign n10076 = n10068 | n10075 ;
  assign n10077 = x88 & n10076 ;
  assign n10078 = x88 | n10076 ;
  assign n22095 = ~n9656 ;
  assign n10079 = n22095 & n9657 ;
  assign n10080 = n146 & n10079 ;
  assign n10081 = n9662 & n10080 ;
  assign n10082 = n9662 | n10080 ;
  assign n22096 = ~n10081 ;
  assign n10083 = n22096 & n10082 ;
  assign n22097 = ~n10083 ;
  assign n10084 = n10078 & n22097 ;
  assign n10085 = n10077 | n10084 ;
  assign n10086 = x89 & n10085 ;
  assign n10087 = x89 | n10085 ;
  assign n22098 = ~n9665 ;
  assign n10088 = n22098 & n9666 ;
  assign n10089 = n146 & n10088 ;
  assign n10090 = n21960 & n10089 ;
  assign n22099 = ~n10089 ;
  assign n10091 = n9671 & n22099 ;
  assign n10092 = n10090 | n10091 ;
  assign n22100 = ~n10092 ;
  assign n10093 = n10087 & n22100 ;
  assign n10094 = n10086 | n10093 ;
  assign n10095 = x90 & n10094 ;
  assign n10096 = x90 | n10094 ;
  assign n22101 = ~n9674 ;
  assign n10097 = n22101 & n9675 ;
  assign n10098 = n146 & n10097 ;
  assign n10099 = n21963 & n10098 ;
  assign n22102 = ~n10098 ;
  assign n10100 = n9680 & n22102 ;
  assign n10101 = n10099 | n10100 ;
  assign n22103 = ~n10101 ;
  assign n10102 = n10096 & n22103 ;
  assign n10103 = n10095 | n10102 ;
  assign n10104 = x91 & n10103 ;
  assign n10105 = x91 | n10103 ;
  assign n22104 = ~n9683 ;
  assign n10106 = n22104 & n9684 ;
  assign n10107 = n146 & n10106 ;
  assign n10108 = n9689 & n10107 ;
  assign n10109 = n9689 | n10107 ;
  assign n22105 = ~n10108 ;
  assign n10110 = n22105 & n10109 ;
  assign n22106 = ~n10110 ;
  assign n10111 = n10105 & n22106 ;
  assign n10112 = n10104 | n10111 ;
  assign n10113 = x92 & n10112 ;
  assign n10114 = x92 | n10112 ;
  assign n22107 = ~n9692 ;
  assign n10115 = n22107 & n9693 ;
  assign n10116 = n146 & n10115 ;
  assign n10117 = n9698 & n10116 ;
  assign n10118 = n9698 | n10116 ;
  assign n22108 = ~n10117 ;
  assign n10119 = n22108 & n10118 ;
  assign n22109 = ~n10119 ;
  assign n10120 = n10114 & n22109 ;
  assign n10121 = n10113 | n10120 ;
  assign n10122 = x93 & n10121 ;
  assign n10123 = x93 | n10121 ;
  assign n22110 = ~n9701 ;
  assign n10124 = n22110 & n9702 ;
  assign n10125 = n146 & n10124 ;
  assign n10126 = n21972 & n10125 ;
  assign n22111 = ~n10125 ;
  assign n10127 = n9707 & n22111 ;
  assign n10128 = n10126 | n10127 ;
  assign n22112 = ~n10128 ;
  assign n10129 = n10123 & n22112 ;
  assign n10130 = n10122 | n10129 ;
  assign n10131 = x94 & n10130 ;
  assign n10132 = x94 | n10130 ;
  assign n22113 = ~n9710 ;
  assign n10133 = n22113 & n9711 ;
  assign n10134 = n146 & n10133 ;
  assign n10135 = n21975 & n10134 ;
  assign n22114 = ~n10134 ;
  assign n10136 = n9716 & n22114 ;
  assign n10137 = n10135 | n10136 ;
  assign n22115 = ~n10137 ;
  assign n10138 = n10132 & n22115 ;
  assign n10139 = n10131 | n10138 ;
  assign n10140 = x95 & n10139 ;
  assign n10141 = x95 | n10139 ;
  assign n22116 = ~n9719 ;
  assign n10142 = n22116 & n9720 ;
  assign n10143 = n146 & n10142 ;
  assign n10144 = n9725 & n10143 ;
  assign n10145 = n9725 | n10143 ;
  assign n22117 = ~n10144 ;
  assign n10146 = n22117 & n10145 ;
  assign n22118 = ~n10146 ;
  assign n10147 = n10141 & n22118 ;
  assign n10148 = n10140 | n10147 ;
  assign n10149 = x96 & n10148 ;
  assign n10150 = x96 | n10148 ;
  assign n22119 = ~n9728 ;
  assign n10151 = n22119 & n9729 ;
  assign n10152 = n146 & n10151 ;
  assign n10153 = n9734 & n10152 ;
  assign n10154 = n9734 | n10152 ;
  assign n22120 = ~n10153 ;
  assign n10155 = n22120 & n10154 ;
  assign n22121 = ~n10155 ;
  assign n10156 = n10150 & n22121 ;
  assign n10157 = n10149 | n10156 ;
  assign n10158 = x97 & n10157 ;
  assign n10159 = x97 | n10157 ;
  assign n22122 = ~n9737 ;
  assign n10160 = n22122 & n9738 ;
  assign n10161 = n146 & n10160 ;
  assign n10162 = n21984 & n10161 ;
  assign n22123 = ~n10161 ;
  assign n10163 = n9743 & n22123 ;
  assign n10164 = n10162 | n10163 ;
  assign n22124 = ~n10164 ;
  assign n10165 = n10159 & n22124 ;
  assign n10166 = n10158 | n10165 ;
  assign n10167 = x98 & n10166 ;
  assign n10168 = x98 | n10166 ;
  assign n22125 = ~n9746 ;
  assign n10169 = n22125 & n9747 ;
  assign n10170 = n146 & n10169 ;
  assign n10171 = n9752 & n10170 ;
  assign n10172 = n9752 | n10170 ;
  assign n22126 = ~n10171 ;
  assign n10173 = n22126 & n10172 ;
  assign n22127 = ~n10173 ;
  assign n10174 = n10168 & n22127 ;
  assign n10175 = n10167 | n10174 ;
  assign n10176 = x99 & n10175 ;
  assign n10177 = x99 | n10175 ;
  assign n22128 = ~n9755 ;
  assign n10178 = n22128 & n9756 ;
  assign n10179 = n146 & n10178 ;
  assign n10180 = n9761 & n10179 ;
  assign n10181 = n9761 | n10179 ;
  assign n22129 = ~n10180 ;
  assign n10182 = n22129 & n10181 ;
  assign n22130 = ~n10182 ;
  assign n10183 = n10177 & n22130 ;
  assign n10184 = n10176 | n10183 ;
  assign n10185 = x100 & n10184 ;
  assign n10186 = x100 | n10184 ;
  assign n22131 = ~n9764 ;
  assign n10187 = n22131 & n9765 ;
  assign n10188 = n146 & n10187 ;
  assign n10189 = n9770 & n10188 ;
  assign n10190 = n9770 | n10188 ;
  assign n22132 = ~n10189 ;
  assign n10191 = n22132 & n10190 ;
  assign n22133 = ~n10191 ;
  assign n10192 = n10186 & n22133 ;
  assign n10193 = n10185 | n10192 ;
  assign n10194 = x101 & n10193 ;
  assign n10195 = x101 | n10193 ;
  assign n22134 = ~n9773 ;
  assign n10196 = n22134 & n9774 ;
  assign n10197 = n146 & n10196 ;
  assign n10198 = n9779 & n10197 ;
  assign n10199 = n9779 | n10197 ;
  assign n22135 = ~n10198 ;
  assign n10200 = n22135 & n10199 ;
  assign n22136 = ~n10200 ;
  assign n10201 = n10195 & n22136 ;
  assign n10202 = n10194 | n10201 ;
  assign n10203 = x102 & n10202 ;
  assign n10204 = x102 | n10202 ;
  assign n22137 = ~n9782 ;
  assign n10205 = n22137 & n9783 ;
  assign n10206 = n146 & n10205 ;
  assign n10207 = n9788 & n10206 ;
  assign n10208 = n9788 | n10206 ;
  assign n22138 = ~n10207 ;
  assign n10209 = n22138 & n10208 ;
  assign n22139 = ~n10209 ;
  assign n10210 = n10204 & n22139 ;
  assign n10211 = n10203 | n10210 ;
  assign n10212 = x103 & n10211 ;
  assign n10213 = x103 | n10211 ;
  assign n22140 = ~n9791 ;
  assign n10214 = n22140 & n9792 ;
  assign n10215 = n146 & n10214 ;
  assign n10216 = n22002 & n10215 ;
  assign n22141 = ~n10215 ;
  assign n10217 = n9797 & n22141 ;
  assign n10218 = n10216 | n10217 ;
  assign n22142 = ~n10218 ;
  assign n10219 = n10213 & n22142 ;
  assign n10220 = n10212 | n10219 ;
  assign n10221 = x104 & n10220 ;
  assign n10222 = x104 | n10220 ;
  assign n22143 = ~n9800 ;
  assign n10223 = n22143 & n9801 ;
  assign n10224 = n146 & n10223 ;
  assign n10225 = n9806 & n10224 ;
  assign n10226 = n9806 | n10224 ;
  assign n22144 = ~n10225 ;
  assign n10227 = n22144 & n10226 ;
  assign n22145 = ~n10227 ;
  assign n10228 = n10222 & n22145 ;
  assign n10229 = n10221 | n10228 ;
  assign n10230 = x105 & n10229 ;
  assign n10231 = x105 | n10229 ;
  assign n22146 = ~n9809 ;
  assign n10232 = n22146 & n9810 ;
  assign n10233 = n146 & n10232 ;
  assign n10234 = n9815 & n10233 ;
  assign n10235 = n9815 | n10233 ;
  assign n22147 = ~n10234 ;
  assign n10236 = n22147 & n10235 ;
  assign n22148 = ~n10236 ;
  assign n10237 = n10231 & n22148 ;
  assign n10238 = n10230 | n10237 ;
  assign n10239 = x106 & n10238 ;
  assign n10240 = x106 | n10238 ;
  assign n22149 = ~n9818 ;
  assign n10241 = n22149 & n9819 ;
  assign n10242 = n146 & n10241 ;
  assign n10243 = n9824 & n10242 ;
  assign n10244 = n9824 | n10242 ;
  assign n22150 = ~n10243 ;
  assign n10245 = n22150 & n10244 ;
  assign n22151 = ~n10245 ;
  assign n10246 = n10240 & n22151 ;
  assign n10247 = n10239 | n10246 ;
  assign n10248 = x107 & n10247 ;
  assign n10249 = x107 | n10247 ;
  assign n22152 = ~n9827 ;
  assign n10250 = n22152 & n9828 ;
  assign n10251 = n146 & n10250 ;
  assign n10252 = n9833 & n10251 ;
  assign n10253 = n9833 | n10251 ;
  assign n22153 = ~n10252 ;
  assign n10254 = n22153 & n10253 ;
  assign n22154 = ~n10254 ;
  assign n10255 = n10249 & n22154 ;
  assign n10256 = n10248 | n10255 ;
  assign n10257 = x108 & n10256 ;
  assign n10258 = x108 | n10256 ;
  assign n22155 = ~n9836 ;
  assign n10259 = n22155 & n9837 ;
  assign n10260 = n146 & n10259 ;
  assign n10261 = n22017 & n10260 ;
  assign n22156 = ~n10260 ;
  assign n10262 = n9842 & n22156 ;
  assign n10263 = n10261 | n10262 ;
  assign n22157 = ~n10263 ;
  assign n10264 = n10258 & n22157 ;
  assign n10265 = n10257 | n10264 ;
  assign n10266 = x109 & n10265 ;
  assign n10267 = x109 | n10265 ;
  assign n22158 = ~n9845 ;
  assign n10268 = n22158 & n9846 ;
  assign n10269 = n146 & n10268 ;
  assign n10270 = n9851 & n10269 ;
  assign n10271 = n9851 | n10269 ;
  assign n22159 = ~n10270 ;
  assign n10272 = n22159 & n10271 ;
  assign n22160 = ~n10272 ;
  assign n10273 = n10267 & n22160 ;
  assign n10274 = n10266 | n10273 ;
  assign n10275 = x110 & n10274 ;
  assign n10276 = x110 | n10274 ;
  assign n22161 = ~n9870 ;
  assign n10277 = n22161 & n10276 ;
  assign n10278 = n10275 | n10277 ;
  assign n10280 = x111 & n10278 ;
  assign n10281 = n18338 | n10280 ;
  assign n10279 = x111 | n10278 ;
  assign n9864 = n9457 | n9861 ;
  assign n10282 = n18348 & n9054 ;
  assign n10283 = n9864 & n10282 ;
  assign n10284 = n21884 | n10283 ;
  assign n22162 = ~n10284 ;
  assign n10285 = n10279 & n22162 ;
  assign n10286 = n10281 | n10285 ;
  assign n22163 = ~n10275 ;
  assign n10287 = n22163 & n10276 ;
  assign n145 = ~n10286 ;
  assign n10288 = n145 & n10287 ;
  assign n10289 = n9870 & n10288 ;
  assign n10290 = n9870 | n10288 ;
  assign n22165 = ~n10289 ;
  assign n10291 = n22165 & n10290 ;
  assign n22166 = ~x15 ;
  assign n10292 = n22166 & x64 ;
  assign n10293 = x65 | n10292 ;
  assign n10294 = x65 & n10292 ;
  assign n10295 = x64 & n145 ;
  assign n10296 = x16 & n10295 ;
  assign n10297 = x16 | n10295 ;
  assign n22167 = ~n10296 ;
  assign n10298 = n22167 & n10297 ;
  assign n22168 = ~n10294 ;
  assign n10299 = n22168 & n10298 ;
  assign n22169 = ~n10299 ;
  assign n10300 = n10293 & n22169 ;
  assign n10302 = x66 & n10300 ;
  assign n10301 = x66 | n10300 ;
  assign n10303 = n9872 & n22028 ;
  assign n10304 = n145 & n10303 ;
  assign n22170 = ~n9875 ;
  assign n10305 = n22170 & n10304 ;
  assign n22171 = ~n10304 ;
  assign n10306 = n9875 & n22171 ;
  assign n10307 = n10305 | n10306 ;
  assign n22172 = ~n10307 ;
  assign n10308 = n10301 & n22172 ;
  assign n10309 = n10302 | n10308 ;
  assign n10310 = x67 & n10309 ;
  assign n10311 = x67 | n10309 ;
  assign n22173 = ~n9877 ;
  assign n9879 = x66 & n22173 ;
  assign n10312 = n18580 & n9877 ;
  assign n10313 = n9879 | n10312 ;
  assign n10314 = n145 & n10313 ;
  assign n10315 = n9885 & n10314 ;
  assign n10316 = n9885 | n10314 ;
  assign n22174 = ~n10315 ;
  assign n10317 = n22174 & n10316 ;
  assign n22175 = ~n10317 ;
  assign n10318 = n10311 & n22175 ;
  assign n10319 = n10310 | n10318 ;
  assign n10320 = x68 & n10319 ;
  assign n10321 = x68 | n10319 ;
  assign n22176 = ~n9888 ;
  assign n10322 = n22176 & n9889 ;
  assign n10323 = n145 & n10322 ;
  assign n10324 = n9894 & n10323 ;
  assign n10325 = n9894 | n10323 ;
  assign n22177 = ~n10324 ;
  assign n10326 = n22177 & n10325 ;
  assign n22178 = ~n10326 ;
  assign n10327 = n10321 & n22178 ;
  assign n10328 = n10320 | n10327 ;
  assign n10329 = x69 & n10328 ;
  assign n10330 = x69 | n10328 ;
  assign n22179 = ~n9897 ;
  assign n10331 = n22179 & n9898 ;
  assign n10332 = n145 & n10331 ;
  assign n10333 = n22037 & n10332 ;
  assign n22180 = ~n10332 ;
  assign n10334 = n9903 & n22180 ;
  assign n10335 = n10333 | n10334 ;
  assign n22181 = ~n10335 ;
  assign n10336 = n10330 & n22181 ;
  assign n10337 = n10329 | n10336 ;
  assign n10338 = x70 & n10337 ;
  assign n10339 = x70 | n10337 ;
  assign n22182 = ~n9906 ;
  assign n10340 = n22182 & n9907 ;
  assign n10341 = n145 & n10340 ;
  assign n10342 = n9912 & n10341 ;
  assign n10343 = n9912 | n10341 ;
  assign n22183 = ~n10342 ;
  assign n10344 = n22183 & n10343 ;
  assign n22184 = ~n10344 ;
  assign n10345 = n10339 & n22184 ;
  assign n10346 = n10338 | n10345 ;
  assign n10347 = x71 & n10346 ;
  assign n10348 = x71 | n10346 ;
  assign n22185 = ~n9915 ;
  assign n10349 = n22185 & n9916 ;
  assign n10350 = n145 & n10349 ;
  assign n10351 = n22043 & n10350 ;
  assign n22186 = ~n10350 ;
  assign n10352 = n9921 & n22186 ;
  assign n10353 = n10351 | n10352 ;
  assign n22187 = ~n10353 ;
  assign n10354 = n10348 & n22187 ;
  assign n10355 = n10347 | n10354 ;
  assign n10356 = x72 & n10355 ;
  assign n10357 = x72 | n10355 ;
  assign n22188 = ~n9924 ;
  assign n10358 = n22188 & n9925 ;
  assign n10359 = n145 & n10358 ;
  assign n10360 = n9930 & n10359 ;
  assign n10361 = n9930 | n10359 ;
  assign n22189 = ~n10360 ;
  assign n10362 = n22189 & n10361 ;
  assign n22190 = ~n10362 ;
  assign n10363 = n10357 & n22190 ;
  assign n10364 = n10356 | n10363 ;
  assign n10365 = x73 & n10364 ;
  assign n10366 = x73 | n10364 ;
  assign n22191 = ~n9933 ;
  assign n10367 = n22191 & n9934 ;
  assign n10368 = n145 & n10367 ;
  assign n10369 = n22049 & n10368 ;
  assign n22192 = ~n10368 ;
  assign n10370 = n9939 & n22192 ;
  assign n10371 = n10369 | n10370 ;
  assign n22193 = ~n10371 ;
  assign n10372 = n10366 & n22193 ;
  assign n10373 = n10365 | n10372 ;
  assign n10374 = x74 & n10373 ;
  assign n10375 = x74 | n10373 ;
  assign n22194 = ~n9942 ;
  assign n10376 = n22194 & n9943 ;
  assign n10377 = n145 & n10376 ;
  assign n10378 = n9948 & n10377 ;
  assign n10379 = n9948 | n10377 ;
  assign n22195 = ~n10378 ;
  assign n10380 = n22195 & n10379 ;
  assign n22196 = ~n10380 ;
  assign n10381 = n10375 & n22196 ;
  assign n10382 = n10374 | n10381 ;
  assign n10383 = x75 & n10382 ;
  assign n10384 = x75 | n10382 ;
  assign n22197 = ~n9951 ;
  assign n10385 = n22197 & n9952 ;
  assign n10386 = n145 & n10385 ;
  assign n10387 = n9957 & n10386 ;
  assign n10388 = n9957 | n10386 ;
  assign n22198 = ~n10387 ;
  assign n10389 = n22198 & n10388 ;
  assign n22199 = ~n10389 ;
  assign n10390 = n10384 & n22199 ;
  assign n10391 = n10383 | n10390 ;
  assign n10392 = x76 & n10391 ;
  assign n10393 = x76 | n10391 ;
  assign n22200 = ~n9960 ;
  assign n10394 = n22200 & n9961 ;
  assign n10395 = n145 & n10394 ;
  assign n10396 = n22058 & n10395 ;
  assign n22201 = ~n10395 ;
  assign n10397 = n9966 & n22201 ;
  assign n10398 = n10396 | n10397 ;
  assign n22202 = ~n10398 ;
  assign n10399 = n10393 & n22202 ;
  assign n10400 = n10392 | n10399 ;
  assign n10401 = x77 & n10400 ;
  assign n10402 = x77 | n10400 ;
  assign n22203 = ~n9969 ;
  assign n10403 = n22203 & n9970 ;
  assign n10404 = n145 & n10403 ;
  assign n10405 = n22061 & n10404 ;
  assign n22204 = ~n10404 ;
  assign n10406 = n9975 & n22204 ;
  assign n10407 = n10405 | n10406 ;
  assign n22205 = ~n10407 ;
  assign n10408 = n10402 & n22205 ;
  assign n10409 = n10401 | n10408 ;
  assign n10410 = x78 & n10409 ;
  assign n10411 = x78 | n10409 ;
  assign n22206 = ~n9978 ;
  assign n10412 = n22206 & n9979 ;
  assign n10413 = n145 & n10412 ;
  assign n10414 = n9984 & n10413 ;
  assign n10415 = n9984 | n10413 ;
  assign n22207 = ~n10414 ;
  assign n10416 = n22207 & n10415 ;
  assign n22208 = ~n10416 ;
  assign n10417 = n10411 & n22208 ;
  assign n10418 = n10410 | n10417 ;
  assign n10419 = x79 & n10418 ;
  assign n10420 = x79 | n10418 ;
  assign n22209 = ~n9987 ;
  assign n10421 = n22209 & n9988 ;
  assign n10422 = n145 & n10421 ;
  assign n10423 = n22067 & n10422 ;
  assign n22210 = ~n10422 ;
  assign n10424 = n9993 & n22210 ;
  assign n10425 = n10423 | n10424 ;
  assign n22211 = ~n10425 ;
  assign n10426 = n10420 & n22211 ;
  assign n10427 = n10419 | n10426 ;
  assign n10428 = x80 & n10427 ;
  assign n10429 = x80 | n10427 ;
  assign n22212 = ~n9996 ;
  assign n10430 = n22212 & n9997 ;
  assign n10431 = n145 & n10430 ;
  assign n10432 = n22070 & n10431 ;
  assign n22213 = ~n10431 ;
  assign n10433 = n10002 & n22213 ;
  assign n10434 = n10432 | n10433 ;
  assign n22214 = ~n10434 ;
  assign n10435 = n10429 & n22214 ;
  assign n10436 = n10428 | n10435 ;
  assign n10437 = x81 & n10436 ;
  assign n10438 = x81 | n10436 ;
  assign n22215 = ~n10005 ;
  assign n10439 = n22215 & n10006 ;
  assign n10440 = n145 & n10439 ;
  assign n10441 = n10011 & n10440 ;
  assign n10442 = n10011 | n10440 ;
  assign n22216 = ~n10441 ;
  assign n10443 = n22216 & n10442 ;
  assign n22217 = ~n10443 ;
  assign n10444 = n10438 & n22217 ;
  assign n10445 = n10437 | n10444 ;
  assign n10446 = x82 & n10445 ;
  assign n10447 = x82 | n10445 ;
  assign n22218 = ~n10014 ;
  assign n10448 = n22218 & n10015 ;
  assign n10449 = n145 & n10448 ;
  assign n10450 = n22076 & n10449 ;
  assign n22219 = ~n10449 ;
  assign n10451 = n10020 & n22219 ;
  assign n10452 = n10450 | n10451 ;
  assign n22220 = ~n10452 ;
  assign n10453 = n10447 & n22220 ;
  assign n10454 = n10446 | n10453 ;
  assign n10455 = x83 & n10454 ;
  assign n10456 = x83 | n10454 ;
  assign n22221 = ~n10023 ;
  assign n10457 = n22221 & n10024 ;
  assign n10458 = n145 & n10457 ;
  assign n10459 = n10029 & n10458 ;
  assign n10460 = n10029 | n10458 ;
  assign n22222 = ~n10459 ;
  assign n10461 = n22222 & n10460 ;
  assign n22223 = ~n10461 ;
  assign n10462 = n10456 & n22223 ;
  assign n10463 = n10455 | n10462 ;
  assign n10464 = x84 & n10463 ;
  assign n10465 = x84 | n10463 ;
  assign n22224 = ~n10032 ;
  assign n10466 = n22224 & n10033 ;
  assign n10467 = n145 & n10466 ;
  assign n10468 = n10038 & n10467 ;
  assign n10469 = n10038 | n10467 ;
  assign n22225 = ~n10468 ;
  assign n10470 = n22225 & n10469 ;
  assign n22226 = ~n10470 ;
  assign n10471 = n10465 & n22226 ;
  assign n10472 = n10464 | n10471 ;
  assign n10473 = x85 & n10472 ;
  assign n10474 = x85 | n10472 ;
  assign n22227 = ~n10041 ;
  assign n10475 = n22227 & n10042 ;
  assign n10476 = n145 & n10475 ;
  assign n10477 = n10047 & n10476 ;
  assign n10478 = n10047 | n10476 ;
  assign n22228 = ~n10477 ;
  assign n10479 = n22228 & n10478 ;
  assign n22229 = ~n10479 ;
  assign n10480 = n10474 & n22229 ;
  assign n10481 = n10473 | n10480 ;
  assign n10482 = x86 & n10481 ;
  assign n10483 = x86 | n10481 ;
  assign n22230 = ~n10050 ;
  assign n10484 = n22230 & n10051 ;
  assign n10485 = n145 & n10484 ;
  assign n10486 = n10056 & n10485 ;
  assign n10487 = n10056 | n10485 ;
  assign n22231 = ~n10486 ;
  assign n10488 = n22231 & n10487 ;
  assign n22232 = ~n10488 ;
  assign n10489 = n10483 & n22232 ;
  assign n10490 = n10482 | n10489 ;
  assign n10491 = x87 & n10490 ;
  assign n10492 = x87 | n10490 ;
  assign n22233 = ~n10059 ;
  assign n10493 = n22233 & n10060 ;
  assign n10494 = n145 & n10493 ;
  assign n10495 = n10065 & n10494 ;
  assign n10496 = n10065 | n10494 ;
  assign n22234 = ~n10495 ;
  assign n10497 = n22234 & n10496 ;
  assign n22235 = ~n10497 ;
  assign n10498 = n10492 & n22235 ;
  assign n10499 = n10491 | n10498 ;
  assign n10500 = x88 & n10499 ;
  assign n10501 = x88 | n10499 ;
  assign n22236 = ~n10068 ;
  assign n10502 = n22236 & n10069 ;
  assign n10503 = n145 & n10502 ;
  assign n10504 = n10074 & n10503 ;
  assign n10505 = n10074 | n10503 ;
  assign n22237 = ~n10504 ;
  assign n10506 = n22237 & n10505 ;
  assign n22238 = ~n10506 ;
  assign n10507 = n10501 & n22238 ;
  assign n10508 = n10500 | n10507 ;
  assign n10509 = x89 & n10508 ;
  assign n10510 = x89 | n10508 ;
  assign n22239 = ~n10077 ;
  assign n10511 = n22239 & n10078 ;
  assign n10512 = n145 & n10511 ;
  assign n10513 = n10083 & n10512 ;
  assign n10514 = n10083 | n10512 ;
  assign n22240 = ~n10513 ;
  assign n10515 = n22240 & n10514 ;
  assign n22241 = ~n10515 ;
  assign n10516 = n10510 & n22241 ;
  assign n10517 = n10509 | n10516 ;
  assign n10518 = x90 & n10517 ;
  assign n10519 = x90 | n10517 ;
  assign n22242 = ~n10086 ;
  assign n10520 = n22242 & n10087 ;
  assign n10521 = n145 & n10520 ;
  assign n10522 = n10092 & n10521 ;
  assign n10523 = n10092 | n10521 ;
  assign n22243 = ~n10522 ;
  assign n10524 = n22243 & n10523 ;
  assign n22244 = ~n10524 ;
  assign n10525 = n10519 & n22244 ;
  assign n10526 = n10518 | n10525 ;
  assign n10527 = x91 & n10526 ;
  assign n10528 = x91 | n10526 ;
  assign n22245 = ~n10095 ;
  assign n10529 = n22245 & n10096 ;
  assign n10530 = n145 & n10529 ;
  assign n10531 = n22103 & n10530 ;
  assign n22246 = ~n10530 ;
  assign n10532 = n10101 & n22246 ;
  assign n10533 = n10531 | n10532 ;
  assign n22247 = ~n10533 ;
  assign n10534 = n10528 & n22247 ;
  assign n10535 = n10527 | n10534 ;
  assign n10536 = x92 & n10535 ;
  assign n10537 = x92 | n10535 ;
  assign n22248 = ~n10104 ;
  assign n10538 = n22248 & n10105 ;
  assign n10539 = n145 & n10538 ;
  assign n10540 = n22106 & n10539 ;
  assign n22249 = ~n10539 ;
  assign n10541 = n10110 & n22249 ;
  assign n10542 = n10540 | n10541 ;
  assign n22250 = ~n10542 ;
  assign n10543 = n10537 & n22250 ;
  assign n10544 = n10536 | n10543 ;
  assign n10545 = x93 & n10544 ;
  assign n10546 = x93 | n10544 ;
  assign n22251 = ~n10113 ;
  assign n10547 = n22251 & n10114 ;
  assign n10548 = n145 & n10547 ;
  assign n10549 = n22109 & n10548 ;
  assign n22252 = ~n10548 ;
  assign n10550 = n10119 & n22252 ;
  assign n10551 = n10549 | n10550 ;
  assign n22253 = ~n10551 ;
  assign n10552 = n10546 & n22253 ;
  assign n10553 = n10545 | n10552 ;
  assign n10554 = x94 & n10553 ;
  assign n10555 = x94 | n10553 ;
  assign n22254 = ~n10122 ;
  assign n10556 = n22254 & n10123 ;
  assign n10557 = n145 & n10556 ;
  assign n10558 = n22112 & n10557 ;
  assign n22255 = ~n10557 ;
  assign n10559 = n10128 & n22255 ;
  assign n10560 = n10558 | n10559 ;
  assign n22256 = ~n10560 ;
  assign n10561 = n10555 & n22256 ;
  assign n10562 = n10554 | n10561 ;
  assign n10563 = x95 & n10562 ;
  assign n10564 = x95 | n10562 ;
  assign n22257 = ~n10131 ;
  assign n10565 = n22257 & n10132 ;
  assign n10566 = n145 & n10565 ;
  assign n10567 = n10137 & n10566 ;
  assign n10568 = n10137 | n10566 ;
  assign n22258 = ~n10567 ;
  assign n10569 = n22258 & n10568 ;
  assign n22259 = ~n10569 ;
  assign n10570 = n10564 & n22259 ;
  assign n10571 = n10563 | n10570 ;
  assign n10572 = x96 & n10571 ;
  assign n10573 = x96 | n10571 ;
  assign n22260 = ~n10140 ;
  assign n10574 = n22260 & n10141 ;
  assign n10575 = n145 & n10574 ;
  assign n10576 = n10146 & n10575 ;
  assign n10577 = n10146 | n10575 ;
  assign n22261 = ~n10576 ;
  assign n10578 = n22261 & n10577 ;
  assign n22262 = ~n10578 ;
  assign n10579 = n10573 & n22262 ;
  assign n10580 = n10572 | n10579 ;
  assign n10581 = x97 & n10580 ;
  assign n10582 = x97 | n10580 ;
  assign n22263 = ~n10149 ;
  assign n10583 = n22263 & n10150 ;
  assign n10584 = n145 & n10583 ;
  assign n10585 = n10155 & n10584 ;
  assign n10586 = n10155 | n10584 ;
  assign n22264 = ~n10585 ;
  assign n10587 = n22264 & n10586 ;
  assign n22265 = ~n10587 ;
  assign n10588 = n10582 & n22265 ;
  assign n10589 = n10581 | n10588 ;
  assign n10590 = x98 & n10589 ;
  assign n10591 = x98 | n10589 ;
  assign n22266 = ~n10158 ;
  assign n10592 = n22266 & n10159 ;
  assign n10593 = n145 & n10592 ;
  assign n10594 = n10164 & n10593 ;
  assign n10595 = n10164 | n10593 ;
  assign n22267 = ~n10594 ;
  assign n10596 = n22267 & n10595 ;
  assign n22268 = ~n10596 ;
  assign n10597 = n10591 & n22268 ;
  assign n10598 = n10590 | n10597 ;
  assign n10599 = x99 & n10598 ;
  assign n10600 = x99 | n10598 ;
  assign n22269 = ~n10167 ;
  assign n10601 = n22269 & n10168 ;
  assign n10602 = n145 & n10601 ;
  assign n10603 = n10173 & n10602 ;
  assign n10604 = n10173 | n10602 ;
  assign n22270 = ~n10603 ;
  assign n10605 = n22270 & n10604 ;
  assign n22271 = ~n10605 ;
  assign n10606 = n10600 & n22271 ;
  assign n10607 = n10599 | n10606 ;
  assign n10608 = x100 & n10607 ;
  assign n10609 = x100 | n10607 ;
  assign n22272 = ~n10176 ;
  assign n10610 = n22272 & n10177 ;
  assign n10611 = n145 & n10610 ;
  assign n10612 = n10182 & n10611 ;
  assign n10613 = n10182 | n10611 ;
  assign n22273 = ~n10612 ;
  assign n10614 = n22273 & n10613 ;
  assign n22274 = ~n10614 ;
  assign n10615 = n10609 & n22274 ;
  assign n10616 = n10608 | n10615 ;
  assign n10617 = x101 & n10616 ;
  assign n10618 = x101 | n10616 ;
  assign n22275 = ~n10185 ;
  assign n10619 = n22275 & n10186 ;
  assign n10620 = n145 & n10619 ;
  assign n10621 = n10191 & n10620 ;
  assign n10622 = n10191 | n10620 ;
  assign n22276 = ~n10621 ;
  assign n10623 = n22276 & n10622 ;
  assign n22277 = ~n10623 ;
  assign n10624 = n10618 & n22277 ;
  assign n10625 = n10617 | n10624 ;
  assign n10626 = x102 & n10625 ;
  assign n10627 = x102 | n10625 ;
  assign n22278 = ~n10194 ;
  assign n10628 = n22278 & n10195 ;
  assign n10629 = n145 & n10628 ;
  assign n10630 = n10200 & n10629 ;
  assign n10631 = n10200 | n10629 ;
  assign n22279 = ~n10630 ;
  assign n10632 = n22279 & n10631 ;
  assign n22280 = ~n10632 ;
  assign n10633 = n10627 & n22280 ;
  assign n10634 = n10626 | n10633 ;
  assign n10635 = x103 & n10634 ;
  assign n10636 = x103 | n10634 ;
  assign n22281 = ~n10203 ;
  assign n10637 = n22281 & n10204 ;
  assign n10638 = n145 & n10637 ;
  assign n10639 = n10209 & n10638 ;
  assign n10640 = n10209 | n10638 ;
  assign n22282 = ~n10639 ;
  assign n10641 = n22282 & n10640 ;
  assign n22283 = ~n10641 ;
  assign n10642 = n10636 & n22283 ;
  assign n10643 = n10635 | n10642 ;
  assign n10644 = x104 & n10643 ;
  assign n10645 = x104 | n10643 ;
  assign n22284 = ~n10212 ;
  assign n10646 = n22284 & n10213 ;
  assign n10647 = n145 & n10646 ;
  assign n10648 = n10218 & n10647 ;
  assign n10649 = n10218 | n10647 ;
  assign n22285 = ~n10648 ;
  assign n10650 = n22285 & n10649 ;
  assign n22286 = ~n10650 ;
  assign n10651 = n10645 & n22286 ;
  assign n10652 = n10644 | n10651 ;
  assign n10653 = x105 & n10652 ;
  assign n10654 = x105 | n10652 ;
  assign n22287 = ~n10221 ;
  assign n10655 = n22287 & n10222 ;
  assign n10656 = n145 & n10655 ;
  assign n10657 = n10227 & n10656 ;
  assign n10658 = n10227 | n10656 ;
  assign n22288 = ~n10657 ;
  assign n10659 = n22288 & n10658 ;
  assign n22289 = ~n10659 ;
  assign n10660 = n10654 & n22289 ;
  assign n10661 = n10653 | n10660 ;
  assign n10662 = x106 & n10661 ;
  assign n10663 = x106 | n10661 ;
  assign n22290 = ~n10230 ;
  assign n10664 = n22290 & n10231 ;
  assign n10665 = n145 & n10664 ;
  assign n10666 = n10236 & n10665 ;
  assign n10667 = n10236 | n10665 ;
  assign n22291 = ~n10666 ;
  assign n10668 = n22291 & n10667 ;
  assign n22292 = ~n10668 ;
  assign n10669 = n10663 & n22292 ;
  assign n10670 = n10662 | n10669 ;
  assign n10671 = x107 & n10670 ;
  assign n10672 = x107 | n10670 ;
  assign n22293 = ~n10239 ;
  assign n10673 = n22293 & n10240 ;
  assign n10674 = n145 & n10673 ;
  assign n10675 = n10245 & n10674 ;
  assign n10676 = n10245 | n10674 ;
  assign n22294 = ~n10675 ;
  assign n10677 = n22294 & n10676 ;
  assign n22295 = ~n10677 ;
  assign n10678 = n10672 & n22295 ;
  assign n10679 = n10671 | n10678 ;
  assign n10680 = x108 & n10679 ;
  assign n10681 = x108 | n10679 ;
  assign n22296 = ~n10248 ;
  assign n10682 = n22296 & n10249 ;
  assign n10683 = n145 & n10682 ;
  assign n10684 = n10254 & n10683 ;
  assign n10685 = n10254 | n10683 ;
  assign n22297 = ~n10684 ;
  assign n10686 = n22297 & n10685 ;
  assign n22298 = ~n10686 ;
  assign n10687 = n10681 & n22298 ;
  assign n10688 = n10680 | n10687 ;
  assign n10689 = x109 & n10688 ;
  assign n10690 = x109 | n10688 ;
  assign n22299 = ~n10257 ;
  assign n10691 = n22299 & n10258 ;
  assign n10692 = n145 & n10691 ;
  assign n10693 = n10263 & n10692 ;
  assign n10694 = n10263 | n10692 ;
  assign n22300 = ~n10693 ;
  assign n10695 = n22300 & n10694 ;
  assign n22301 = ~n10695 ;
  assign n10696 = n10690 & n22301 ;
  assign n10697 = n10689 | n10696 ;
  assign n10698 = x110 & n10697 ;
  assign n10699 = x110 | n10697 ;
  assign n22302 = ~n10266 ;
  assign n10700 = n22302 & n10267 ;
  assign n10701 = n145 & n10700 ;
  assign n10702 = n10272 & n10701 ;
  assign n10703 = n10272 | n10701 ;
  assign n22303 = ~n10702 ;
  assign n10704 = n22303 & n10703 ;
  assign n22304 = ~n10704 ;
  assign n10705 = n10699 & n22304 ;
  assign n10706 = n10698 | n10705 ;
  assign n10707 = x111 & n10706 ;
  assign n10708 = x111 | n10706 ;
  assign n22305 = ~n10291 ;
  assign n10709 = n22305 & n10708 ;
  assign n10710 = n10707 | n10709 ;
  assign n22306 = ~n10281 ;
  assign n10711 = n10279 & n22306 ;
  assign n22307 = ~n10711 ;
  assign n10712 = n10284 & n22307 ;
  assign n22308 = ~x112 ;
  assign n10713 = n22308 & n10712 ;
  assign n22309 = ~n10713 ;
  assign n10714 = n10710 & n22309 ;
  assign n22310 = ~n10712 ;
  assign n10715 = x112 & n22310 ;
  assign n10716 = n18333 | n10715 ;
  assign n10717 = n10714 | n10716 ;
  assign n22311 = ~n10707 ;
  assign n10718 = n22311 & n10708 ;
  assign n144 = ~n10717 ;
  assign n10719 = n144 & n10718 ;
  assign n10720 = n10291 & n10719 ;
  assign n10721 = n10291 | n10719 ;
  assign n22313 = ~n10720 ;
  assign n10722 = n22313 & n10721 ;
  assign n10723 = x112 & n10710 ;
  assign n10724 = x112 | n10710 ;
  assign n22314 = ~n18333 ;
  assign n10725 = n22314 & n10724 ;
  assign n22315 = ~n10723 ;
  assign n10726 = n22315 & n10725 ;
  assign n22316 = ~n10726 ;
  assign n10727 = n10712 & n22316 ;
  assign n10728 = n22314 & n10727 ;
  assign n22317 = ~x14 ;
  assign n10729 = n22317 & x64 ;
  assign n10730 = x65 | n10729 ;
  assign n10731 = x65 & n10729 ;
  assign n10732 = x64 & n144 ;
  assign n10733 = x15 & n10732 ;
  assign n10734 = x15 | n10732 ;
  assign n22318 = ~n10733 ;
  assign n10735 = n22318 & n10734 ;
  assign n22319 = ~n10731 ;
  assign n10736 = n22319 & n10735 ;
  assign n22320 = ~n10736 ;
  assign n10737 = n10730 & n22320 ;
  assign n10739 = x66 | n10737 ;
  assign n10738 = x66 & n10737 ;
  assign n10740 = n10293 & n22168 ;
  assign n10741 = n144 & n10740 ;
  assign n22321 = ~n10298 ;
  assign n10742 = n22321 & n10741 ;
  assign n22322 = ~n10741 ;
  assign n10743 = n10298 & n22322 ;
  assign n10744 = n10742 | n10743 ;
  assign n22323 = ~n10738 ;
  assign n10745 = n22323 & n10744 ;
  assign n22324 = ~n10745 ;
  assign n10746 = n10739 & n22324 ;
  assign n10747 = x67 | n10746 ;
  assign n10748 = x67 & n10746 ;
  assign n10749 = n10302 | n10717 ;
  assign n22325 = ~n10749 ;
  assign n10750 = n10308 & n22325 ;
  assign n10751 = n10301 & n22325 ;
  assign n22326 = ~n10751 ;
  assign n10752 = n10307 & n22326 ;
  assign n10753 = n10750 | n10752 ;
  assign n22327 = ~n10748 ;
  assign n10754 = n22327 & n10753 ;
  assign n22328 = ~n10754 ;
  assign n10755 = n10747 & n22328 ;
  assign n10756 = x68 | n10755 ;
  assign n10757 = x68 & n10755 ;
  assign n22329 = ~n10310 ;
  assign n10758 = n22329 & n10311 ;
  assign n10759 = n144 & n10758 ;
  assign n10760 = n10317 & n10759 ;
  assign n10761 = n10317 | n10759 ;
  assign n22330 = ~n10760 ;
  assign n10762 = n22330 & n10761 ;
  assign n22331 = ~n10757 ;
  assign n10763 = n22331 & n10762 ;
  assign n22332 = ~n10763 ;
  assign n10764 = n10756 & n22332 ;
  assign n10765 = x69 | n10764 ;
  assign n10766 = x69 & n10764 ;
  assign n22333 = ~n10320 ;
  assign n10767 = n22333 & n10321 ;
  assign n10768 = n144 & n10767 ;
  assign n10769 = n10326 & n10768 ;
  assign n10770 = n10326 | n10768 ;
  assign n22334 = ~n10769 ;
  assign n10771 = n22334 & n10770 ;
  assign n22335 = ~n10766 ;
  assign n10772 = n22335 & n10771 ;
  assign n22336 = ~n10772 ;
  assign n10773 = n10765 & n22336 ;
  assign n10774 = x70 | n10773 ;
  assign n10775 = x70 & n10773 ;
  assign n22337 = ~n10329 ;
  assign n10776 = n22337 & n10330 ;
  assign n10777 = n144 & n10776 ;
  assign n10778 = n10335 & n10777 ;
  assign n10779 = n10335 | n10777 ;
  assign n22338 = ~n10778 ;
  assign n10780 = n22338 & n10779 ;
  assign n22339 = ~n10775 ;
  assign n10781 = n22339 & n10780 ;
  assign n22340 = ~n10781 ;
  assign n10782 = n10774 & n22340 ;
  assign n10783 = x71 | n10782 ;
  assign n10784 = x71 & n10782 ;
  assign n22341 = ~n10338 ;
  assign n10785 = n22341 & n10339 ;
  assign n10786 = n144 & n10785 ;
  assign n10787 = n10344 & n10786 ;
  assign n10788 = n10344 | n10786 ;
  assign n22342 = ~n10787 ;
  assign n10789 = n22342 & n10788 ;
  assign n22343 = ~n10784 ;
  assign n10790 = n22343 & n10789 ;
  assign n22344 = ~n10790 ;
  assign n10791 = n10783 & n22344 ;
  assign n10792 = x72 | n10791 ;
  assign n10793 = x72 & n10791 ;
  assign n22345 = ~n10347 ;
  assign n10794 = n22345 & n10348 ;
  assign n10795 = n144 & n10794 ;
  assign n10796 = n10353 & n10795 ;
  assign n10797 = n10353 | n10795 ;
  assign n22346 = ~n10796 ;
  assign n10798 = n22346 & n10797 ;
  assign n22347 = ~n10793 ;
  assign n10799 = n22347 & n10798 ;
  assign n22348 = ~n10799 ;
  assign n10800 = n10792 & n22348 ;
  assign n10801 = x73 | n10800 ;
  assign n10802 = x73 & n10800 ;
  assign n22349 = ~n10356 ;
  assign n10803 = n22349 & n10357 ;
  assign n10804 = n144 & n10803 ;
  assign n10805 = n22190 & n10804 ;
  assign n22350 = ~n10804 ;
  assign n10806 = n10362 & n22350 ;
  assign n10807 = n10805 | n10806 ;
  assign n22351 = ~n10802 ;
  assign n10808 = n22351 & n10807 ;
  assign n22352 = ~n10808 ;
  assign n10809 = n10801 & n22352 ;
  assign n10810 = x74 | n10809 ;
  assign n10811 = x74 & n10809 ;
  assign n22353 = ~n10365 ;
  assign n10812 = n22353 & n10366 ;
  assign n10813 = n144 & n10812 ;
  assign n10814 = n22193 & n10813 ;
  assign n22354 = ~n10813 ;
  assign n10815 = n10371 & n22354 ;
  assign n10816 = n10814 | n10815 ;
  assign n22355 = ~n10811 ;
  assign n10817 = n22355 & n10816 ;
  assign n22356 = ~n10817 ;
  assign n10818 = n10810 & n22356 ;
  assign n10819 = x75 | n10818 ;
  assign n10820 = x75 & n10818 ;
  assign n22357 = ~n10374 ;
  assign n10821 = n22357 & n10375 ;
  assign n10822 = n144 & n10821 ;
  assign n10823 = n10380 & n10822 ;
  assign n10824 = n10380 | n10822 ;
  assign n22358 = ~n10823 ;
  assign n10825 = n22358 & n10824 ;
  assign n22359 = ~n10820 ;
  assign n10826 = n22359 & n10825 ;
  assign n22360 = ~n10826 ;
  assign n10827 = n10819 & n22360 ;
  assign n10828 = x76 | n10827 ;
  assign n10829 = x76 & n10827 ;
  assign n22361 = ~n10383 ;
  assign n10830 = n22361 & n10384 ;
  assign n10831 = n144 & n10830 ;
  assign n10832 = n10389 & n10831 ;
  assign n10833 = n10389 | n10831 ;
  assign n22362 = ~n10832 ;
  assign n10834 = n22362 & n10833 ;
  assign n22363 = ~n10829 ;
  assign n10835 = n22363 & n10834 ;
  assign n22364 = ~n10835 ;
  assign n10836 = n10828 & n22364 ;
  assign n10837 = x77 | n10836 ;
  assign n10838 = x77 & n10836 ;
  assign n22365 = ~n10392 ;
  assign n10839 = n22365 & n10393 ;
  assign n10840 = n144 & n10839 ;
  assign n10841 = n22202 & n10840 ;
  assign n22366 = ~n10840 ;
  assign n10842 = n10398 & n22366 ;
  assign n10843 = n10841 | n10842 ;
  assign n22367 = ~n10838 ;
  assign n10844 = n22367 & n10843 ;
  assign n22368 = ~n10844 ;
  assign n10845 = n10837 & n22368 ;
  assign n10846 = x78 | n10845 ;
  assign n10847 = x78 & n10845 ;
  assign n22369 = ~n10401 ;
  assign n10848 = n22369 & n10402 ;
  assign n10849 = n144 & n10848 ;
  assign n10850 = n10407 & n10849 ;
  assign n10851 = n10407 | n10849 ;
  assign n22370 = ~n10850 ;
  assign n10852 = n22370 & n10851 ;
  assign n22371 = ~n10847 ;
  assign n10853 = n22371 & n10852 ;
  assign n22372 = ~n10853 ;
  assign n10854 = n10846 & n22372 ;
  assign n10855 = x79 | n10854 ;
  assign n10856 = x79 & n10854 ;
  assign n22373 = ~n10410 ;
  assign n10857 = n22373 & n10411 ;
  assign n10858 = n144 & n10857 ;
  assign n10859 = n22208 & n10858 ;
  assign n22374 = ~n10858 ;
  assign n10860 = n10416 & n22374 ;
  assign n10861 = n10859 | n10860 ;
  assign n22375 = ~n10856 ;
  assign n10862 = n22375 & n10861 ;
  assign n22376 = ~n10862 ;
  assign n10863 = n10855 & n22376 ;
  assign n10864 = x80 | n10863 ;
  assign n10865 = x80 & n10863 ;
  assign n22377 = ~n10419 ;
  assign n10866 = n22377 & n10420 ;
  assign n10867 = n144 & n10866 ;
  assign n10868 = n22211 & n10867 ;
  assign n22378 = ~n10867 ;
  assign n10869 = n10425 & n22378 ;
  assign n10870 = n10868 | n10869 ;
  assign n22379 = ~n10865 ;
  assign n10871 = n22379 & n10870 ;
  assign n22380 = ~n10871 ;
  assign n10872 = n10864 & n22380 ;
  assign n10873 = x81 | n10872 ;
  assign n10874 = x81 & n10872 ;
  assign n22381 = ~n10428 ;
  assign n10875 = n22381 & n10429 ;
  assign n10876 = n144 & n10875 ;
  assign n10877 = n22214 & n10876 ;
  assign n22382 = ~n10876 ;
  assign n10878 = n10434 & n22382 ;
  assign n10879 = n10877 | n10878 ;
  assign n22383 = ~n10874 ;
  assign n10880 = n22383 & n10879 ;
  assign n22384 = ~n10880 ;
  assign n10881 = n10873 & n22384 ;
  assign n10882 = x82 | n10881 ;
  assign n10883 = x82 & n10881 ;
  assign n22385 = ~n10437 ;
  assign n10884 = n22385 & n10438 ;
  assign n10885 = n144 & n10884 ;
  assign n10886 = n10443 & n10885 ;
  assign n10887 = n10443 | n10885 ;
  assign n22386 = ~n10886 ;
  assign n10888 = n22386 & n10887 ;
  assign n22387 = ~n10883 ;
  assign n10889 = n22387 & n10888 ;
  assign n22388 = ~n10889 ;
  assign n10890 = n10882 & n22388 ;
  assign n10891 = x83 | n10890 ;
  assign n10892 = x83 & n10890 ;
  assign n22389 = ~n10446 ;
  assign n10893 = n22389 & n10447 ;
  assign n10894 = n144 & n10893 ;
  assign n10895 = n10452 & n10894 ;
  assign n10896 = n10452 | n10894 ;
  assign n22390 = ~n10895 ;
  assign n10897 = n22390 & n10896 ;
  assign n22391 = ~n10892 ;
  assign n10898 = n22391 & n10897 ;
  assign n22392 = ~n10898 ;
  assign n10899 = n10891 & n22392 ;
  assign n10900 = x84 | n10899 ;
  assign n10901 = x84 & n10899 ;
  assign n22393 = ~n10455 ;
  assign n10902 = n22393 & n10456 ;
  assign n10903 = n144 & n10902 ;
  assign n10904 = n22223 & n10903 ;
  assign n22394 = ~n10903 ;
  assign n10905 = n10461 & n22394 ;
  assign n10906 = n10904 | n10905 ;
  assign n22395 = ~n10901 ;
  assign n10907 = n22395 & n10906 ;
  assign n22396 = ~n10907 ;
  assign n10908 = n10900 & n22396 ;
  assign n10909 = x85 | n10908 ;
  assign n10910 = x85 & n10908 ;
  assign n22397 = ~n10464 ;
  assign n10911 = n22397 & n10465 ;
  assign n10912 = n144 & n10911 ;
  assign n10913 = n22226 & n10912 ;
  assign n22398 = ~n10912 ;
  assign n10914 = n10470 & n22398 ;
  assign n10915 = n10913 | n10914 ;
  assign n22399 = ~n10910 ;
  assign n10916 = n22399 & n10915 ;
  assign n22400 = ~n10916 ;
  assign n10917 = n10909 & n22400 ;
  assign n10918 = x86 | n10917 ;
  assign n10919 = x86 & n10917 ;
  assign n22401 = ~n10473 ;
  assign n10920 = n22401 & n10474 ;
  assign n10921 = n144 & n10920 ;
  assign n10922 = n10479 & n10921 ;
  assign n10923 = n10479 | n10921 ;
  assign n22402 = ~n10922 ;
  assign n10924 = n22402 & n10923 ;
  assign n22403 = ~n10919 ;
  assign n10925 = n22403 & n10924 ;
  assign n22404 = ~n10925 ;
  assign n10926 = n10918 & n22404 ;
  assign n10927 = x87 | n10926 ;
  assign n10928 = x87 & n10926 ;
  assign n22405 = ~n10482 ;
  assign n10929 = n22405 & n10483 ;
  assign n10930 = n144 & n10929 ;
  assign n10931 = n10488 & n10930 ;
  assign n10932 = n10488 | n10930 ;
  assign n22406 = ~n10931 ;
  assign n10933 = n22406 & n10932 ;
  assign n22407 = ~n10928 ;
  assign n10934 = n22407 & n10933 ;
  assign n22408 = ~n10934 ;
  assign n10935 = n10927 & n22408 ;
  assign n10936 = x88 | n10935 ;
  assign n10937 = x88 & n10935 ;
  assign n22409 = ~n10491 ;
  assign n10938 = n22409 & n10492 ;
  assign n10939 = n144 & n10938 ;
  assign n10940 = n10497 & n10939 ;
  assign n10941 = n10497 | n10939 ;
  assign n22410 = ~n10940 ;
  assign n10942 = n22410 & n10941 ;
  assign n22411 = ~n10937 ;
  assign n10943 = n22411 & n10942 ;
  assign n22412 = ~n10943 ;
  assign n10944 = n10936 & n22412 ;
  assign n10945 = x89 | n10944 ;
  assign n10946 = x89 & n10944 ;
  assign n22413 = ~n10500 ;
  assign n10947 = n22413 & n10501 ;
  assign n10948 = n144 & n10947 ;
  assign n10949 = n10506 & n10948 ;
  assign n10950 = n10506 | n10948 ;
  assign n22414 = ~n10949 ;
  assign n10951 = n22414 & n10950 ;
  assign n22415 = ~n10946 ;
  assign n10952 = n22415 & n10951 ;
  assign n22416 = ~n10952 ;
  assign n10953 = n10945 & n22416 ;
  assign n10954 = x90 | n10953 ;
  assign n10955 = x90 & n10953 ;
  assign n22417 = ~n10509 ;
  assign n10956 = n22417 & n10510 ;
  assign n10957 = n144 & n10956 ;
  assign n10958 = n10515 & n10957 ;
  assign n10959 = n10515 | n10957 ;
  assign n22418 = ~n10958 ;
  assign n10960 = n22418 & n10959 ;
  assign n22419 = ~n10955 ;
  assign n10961 = n22419 & n10960 ;
  assign n22420 = ~n10961 ;
  assign n10962 = n10954 & n22420 ;
  assign n10963 = x91 | n10962 ;
  assign n10964 = x91 & n10962 ;
  assign n22421 = ~n10518 ;
  assign n10965 = n22421 & n10519 ;
  assign n10966 = n144 & n10965 ;
  assign n10967 = n10524 & n10966 ;
  assign n10968 = n10524 | n10966 ;
  assign n22422 = ~n10967 ;
  assign n10969 = n22422 & n10968 ;
  assign n22423 = ~n10964 ;
  assign n10970 = n22423 & n10969 ;
  assign n22424 = ~n10970 ;
  assign n10971 = n10963 & n22424 ;
  assign n10972 = x92 | n10971 ;
  assign n10973 = x92 & n10971 ;
  assign n22425 = ~n10527 ;
  assign n10974 = n22425 & n10528 ;
  assign n10975 = n144 & n10974 ;
  assign n10976 = n10533 & n10975 ;
  assign n10977 = n10533 | n10975 ;
  assign n22426 = ~n10976 ;
  assign n10978 = n22426 & n10977 ;
  assign n22427 = ~n10973 ;
  assign n10979 = n22427 & n10978 ;
  assign n22428 = ~n10979 ;
  assign n10980 = n10972 & n22428 ;
  assign n10981 = x93 | n10980 ;
  assign n10982 = x93 & n10980 ;
  assign n22429 = ~n10536 ;
  assign n10983 = n22429 & n10537 ;
  assign n10984 = n144 & n10983 ;
  assign n10985 = n22250 & n10984 ;
  assign n22430 = ~n10984 ;
  assign n10986 = n10542 & n22430 ;
  assign n10987 = n10985 | n10986 ;
  assign n22431 = ~n10982 ;
  assign n10988 = n22431 & n10987 ;
  assign n22432 = ~n10988 ;
  assign n10989 = n10981 & n22432 ;
  assign n10990 = x94 | n10989 ;
  assign n10991 = x94 & n10989 ;
  assign n22433 = ~n10545 ;
  assign n10992 = n22433 & n10546 ;
  assign n10993 = n144 & n10992 ;
  assign n10994 = n22253 & n10993 ;
  assign n22434 = ~n10993 ;
  assign n10995 = n10551 & n22434 ;
  assign n10996 = n10994 | n10995 ;
  assign n22435 = ~n10991 ;
  assign n10997 = n22435 & n10996 ;
  assign n22436 = ~n10997 ;
  assign n10998 = n10990 & n22436 ;
  assign n10999 = x95 | n10998 ;
  assign n11000 = x95 & n10998 ;
  assign n22437 = ~n10554 ;
  assign n11001 = n22437 & n10555 ;
  assign n11002 = n144 & n11001 ;
  assign n11003 = n10560 & n11002 ;
  assign n11004 = n10560 | n11002 ;
  assign n22438 = ~n11003 ;
  assign n11005 = n22438 & n11004 ;
  assign n22439 = ~n11000 ;
  assign n11006 = n22439 & n11005 ;
  assign n22440 = ~n11006 ;
  assign n11007 = n10999 & n22440 ;
  assign n11008 = x96 | n11007 ;
  assign n11009 = x96 & n11007 ;
  assign n22441 = ~n10563 ;
  assign n11010 = n22441 & n10564 ;
  assign n11011 = n144 & n11010 ;
  assign n11012 = n10569 & n11011 ;
  assign n11013 = n10569 | n11011 ;
  assign n22442 = ~n11012 ;
  assign n11014 = n22442 & n11013 ;
  assign n22443 = ~n11009 ;
  assign n11015 = n22443 & n11014 ;
  assign n22444 = ~n11015 ;
  assign n11016 = n11008 & n22444 ;
  assign n11017 = x97 | n11016 ;
  assign n11018 = x97 & n11016 ;
  assign n22445 = ~n10572 ;
  assign n11019 = n22445 & n10573 ;
  assign n11020 = n144 & n11019 ;
  assign n11021 = n10578 & n11020 ;
  assign n11022 = n10578 | n11020 ;
  assign n22446 = ~n11021 ;
  assign n11023 = n22446 & n11022 ;
  assign n22447 = ~n11018 ;
  assign n11024 = n22447 & n11023 ;
  assign n22448 = ~n11024 ;
  assign n11025 = n11017 & n22448 ;
  assign n11026 = x98 | n11025 ;
  assign n11027 = x98 & n11025 ;
  assign n22449 = ~n10581 ;
  assign n11028 = n22449 & n10582 ;
  assign n11029 = n144 & n11028 ;
  assign n11030 = n22265 & n11029 ;
  assign n22450 = ~n11029 ;
  assign n11031 = n10587 & n22450 ;
  assign n11032 = n11030 | n11031 ;
  assign n22451 = ~n11027 ;
  assign n11033 = n22451 & n11032 ;
  assign n22452 = ~n11033 ;
  assign n11034 = n11026 & n22452 ;
  assign n11035 = x99 | n11034 ;
  assign n11036 = x99 & n11034 ;
  assign n22453 = ~n10590 ;
  assign n11037 = n22453 & n10591 ;
  assign n11038 = n144 & n11037 ;
  assign n11039 = n10596 & n11038 ;
  assign n11040 = n10596 | n11038 ;
  assign n22454 = ~n11039 ;
  assign n11041 = n22454 & n11040 ;
  assign n22455 = ~n11036 ;
  assign n11042 = n22455 & n11041 ;
  assign n22456 = ~n11042 ;
  assign n11043 = n11035 & n22456 ;
  assign n11044 = x100 | n11043 ;
  assign n11045 = x100 & n11043 ;
  assign n22457 = ~n10599 ;
  assign n11046 = n22457 & n10600 ;
  assign n11047 = n144 & n11046 ;
  assign n11048 = n10605 & n11047 ;
  assign n11049 = n10605 | n11047 ;
  assign n22458 = ~n11048 ;
  assign n11050 = n22458 & n11049 ;
  assign n22459 = ~n11045 ;
  assign n11051 = n22459 & n11050 ;
  assign n22460 = ~n11051 ;
  assign n11052 = n11044 & n22460 ;
  assign n11053 = x101 | n11052 ;
  assign n11054 = x101 & n11052 ;
  assign n22461 = ~n10608 ;
  assign n11055 = n22461 & n10609 ;
  assign n11056 = n144 & n11055 ;
  assign n11057 = n22274 & n11056 ;
  assign n22462 = ~n11056 ;
  assign n11058 = n10614 & n22462 ;
  assign n11059 = n11057 | n11058 ;
  assign n22463 = ~n11054 ;
  assign n11060 = n22463 & n11059 ;
  assign n22464 = ~n11060 ;
  assign n11061 = n11053 & n22464 ;
  assign n11062 = x102 | n11061 ;
  assign n11063 = x102 & n11061 ;
  assign n22465 = ~n10617 ;
  assign n11064 = n22465 & n10618 ;
  assign n11065 = n144 & n11064 ;
  assign n11066 = n10623 & n11065 ;
  assign n11067 = n10623 | n11065 ;
  assign n22466 = ~n11066 ;
  assign n11068 = n22466 & n11067 ;
  assign n22467 = ~n11063 ;
  assign n11069 = n22467 & n11068 ;
  assign n22468 = ~n11069 ;
  assign n11070 = n11062 & n22468 ;
  assign n11071 = x103 | n11070 ;
  assign n11072 = x103 & n11070 ;
  assign n22469 = ~n10626 ;
  assign n11073 = n22469 & n10627 ;
  assign n11074 = n144 & n11073 ;
  assign n11075 = n10632 & n11074 ;
  assign n11076 = n10632 | n11074 ;
  assign n22470 = ~n11075 ;
  assign n11077 = n22470 & n11076 ;
  assign n22471 = ~n11072 ;
  assign n11078 = n22471 & n11077 ;
  assign n22472 = ~n11078 ;
  assign n11079 = n11071 & n22472 ;
  assign n11080 = x104 | n11079 ;
  assign n11081 = x104 & n11079 ;
  assign n22473 = ~n10635 ;
  assign n11082 = n22473 & n10636 ;
  assign n11083 = n144 & n11082 ;
  assign n11084 = n10641 & n11083 ;
  assign n11085 = n10641 | n11083 ;
  assign n22474 = ~n11084 ;
  assign n11086 = n22474 & n11085 ;
  assign n22475 = ~n11081 ;
  assign n11087 = n22475 & n11086 ;
  assign n22476 = ~n11087 ;
  assign n11088 = n11080 & n22476 ;
  assign n11089 = x105 | n11088 ;
  assign n11090 = x105 & n11088 ;
  assign n22477 = ~n10644 ;
  assign n11091 = n22477 & n10645 ;
  assign n11092 = n144 & n11091 ;
  assign n11093 = n10650 & n11092 ;
  assign n11094 = n10650 | n11092 ;
  assign n22478 = ~n11093 ;
  assign n11095 = n22478 & n11094 ;
  assign n22479 = ~n11090 ;
  assign n11096 = n22479 & n11095 ;
  assign n22480 = ~n11096 ;
  assign n11097 = n11089 & n22480 ;
  assign n11098 = x106 | n11097 ;
  assign n11099 = x106 & n11097 ;
  assign n22481 = ~n10653 ;
  assign n11100 = n22481 & n10654 ;
  assign n11101 = n144 & n11100 ;
  assign n11102 = n10659 & n11101 ;
  assign n11103 = n10659 | n11101 ;
  assign n22482 = ~n11102 ;
  assign n11104 = n22482 & n11103 ;
  assign n22483 = ~n11099 ;
  assign n11105 = n22483 & n11104 ;
  assign n22484 = ~n11105 ;
  assign n11106 = n11098 & n22484 ;
  assign n11107 = x107 | n11106 ;
  assign n11108 = x107 & n11106 ;
  assign n22485 = ~n10662 ;
  assign n11109 = n22485 & n10663 ;
  assign n11110 = n144 & n11109 ;
  assign n11111 = n22292 & n11110 ;
  assign n22486 = ~n11110 ;
  assign n11112 = n10668 & n22486 ;
  assign n11113 = n11111 | n11112 ;
  assign n22487 = ~n11108 ;
  assign n11114 = n22487 & n11113 ;
  assign n22488 = ~n11114 ;
  assign n11115 = n11107 & n22488 ;
  assign n11116 = x108 | n11115 ;
  assign n11117 = x108 & n11115 ;
  assign n22489 = ~n10671 ;
  assign n11118 = n22489 & n10672 ;
  assign n11119 = n144 & n11118 ;
  assign n11120 = n22295 & n11119 ;
  assign n22490 = ~n11119 ;
  assign n11121 = n10677 & n22490 ;
  assign n11122 = n11120 | n11121 ;
  assign n22491 = ~n11117 ;
  assign n11123 = n22491 & n11122 ;
  assign n22492 = ~n11123 ;
  assign n11124 = n11116 & n22492 ;
  assign n11125 = x109 | n11124 ;
  assign n11126 = x109 & n11124 ;
  assign n22493 = ~n10680 ;
  assign n11127 = n22493 & n10681 ;
  assign n11128 = n144 & n11127 ;
  assign n11129 = n22298 & n11128 ;
  assign n22494 = ~n11128 ;
  assign n11130 = n10686 & n22494 ;
  assign n11131 = n11129 | n11130 ;
  assign n22495 = ~n11126 ;
  assign n11132 = n22495 & n11131 ;
  assign n22496 = ~n11132 ;
  assign n11133 = n11125 & n22496 ;
  assign n11134 = x110 | n11133 ;
  assign n11135 = x110 & n11133 ;
  assign n22497 = ~n10689 ;
  assign n11136 = n22497 & n10690 ;
  assign n11137 = n144 & n11136 ;
  assign n11138 = n10695 & n11137 ;
  assign n11139 = n10695 | n11137 ;
  assign n22498 = ~n11138 ;
  assign n11140 = n22498 & n11139 ;
  assign n22499 = ~n11135 ;
  assign n11141 = n22499 & n11140 ;
  assign n22500 = ~n11141 ;
  assign n11142 = n11134 & n22500 ;
  assign n11143 = x111 | n11142 ;
  assign n11144 = x111 & n11142 ;
  assign n22501 = ~n10698 ;
  assign n11145 = n22501 & n10699 ;
  assign n11146 = n144 & n11145 ;
  assign n11147 = n22304 & n11146 ;
  assign n22502 = ~n11146 ;
  assign n11148 = n10704 & n22502 ;
  assign n11149 = n11147 | n11148 ;
  assign n22503 = ~n11144 ;
  assign n11150 = n22503 & n11149 ;
  assign n22504 = ~n11150 ;
  assign n11151 = n11143 & n22504 ;
  assign n11153 = x112 | n11151 ;
  assign n22505 = ~n10722 ;
  assign n11154 = n22505 & n11153 ;
  assign n11152 = x112 & n11151 ;
  assign n11155 = x113 & n22310 ;
  assign n11156 = n18328 | n11155 ;
  assign n22506 = ~x113 ;
  assign n11157 = n22506 & n10727 ;
  assign n11158 = n11156 | n11157 ;
  assign n11159 = n11152 | n11158 ;
  assign n11160 = n11154 | n11159 ;
  assign n22507 = ~n10728 ;
  assign n11161 = n22507 & n11160 ;
  assign n22508 = ~n11152 ;
  assign n11162 = n22508 & n11153 ;
  assign n143 = ~n11161 ;
  assign n11163 = n143 & n11162 ;
  assign n11164 = n22505 & n11163 ;
  assign n22510 = ~n11163 ;
  assign n11165 = n10722 & n22510 ;
  assign n11166 = n11164 | n11165 ;
  assign n22511 = ~x13 ;
  assign n11167 = n22511 & x64 ;
  assign n11168 = x65 | n11167 ;
  assign n11169 = x64 & n143 ;
  assign n22512 = ~n11169 ;
  assign n11170 = x14 & n22512 ;
  assign n11171 = n10729 & n143 ;
  assign n11172 = n11170 | n11171 ;
  assign n11173 = x65 & n11167 ;
  assign n22513 = ~n11173 ;
  assign n11174 = n11172 & n22513 ;
  assign n22514 = ~n11174 ;
  assign n11175 = n11168 & n22514 ;
  assign n11176 = x66 & n11175 ;
  assign n11177 = n10730 & n22319 ;
  assign n11178 = n143 & n11177 ;
  assign n11179 = n10735 & n11178 ;
  assign n11180 = n10735 | n11178 ;
  assign n22515 = ~n11179 ;
  assign n11181 = n22515 & n11180 ;
  assign n11182 = x66 | n11175 ;
  assign n22516 = ~n11181 ;
  assign n11183 = n22516 & n11182 ;
  assign n11184 = n11176 | n11183 ;
  assign n11185 = x67 & n11184 ;
  assign n11186 = x67 | n11184 ;
  assign n11187 = n10739 & n143 ;
  assign n11188 = n10745 & n11187 ;
  assign n11189 = n22323 & n11187 ;
  assign n11190 = n10744 | n11189 ;
  assign n22517 = ~n11188 ;
  assign n11191 = n22517 & n11190 ;
  assign n22518 = ~n11191 ;
  assign n11192 = n11186 & n22518 ;
  assign n11193 = n11185 | n11192 ;
  assign n11194 = x68 & n11193 ;
  assign n11195 = x68 | n11193 ;
  assign n11196 = n10747 & n22327 ;
  assign n11197 = n143 & n11196 ;
  assign n22519 = ~n10753 ;
  assign n11198 = n22519 & n11197 ;
  assign n22520 = ~n11197 ;
  assign n11199 = n10753 & n22520 ;
  assign n11200 = n11198 | n11199 ;
  assign n22521 = ~n11200 ;
  assign n11201 = n11195 & n22521 ;
  assign n11202 = n11194 | n11201 ;
  assign n11203 = x69 & n11202 ;
  assign n11204 = x69 | n11202 ;
  assign n11205 = n10756 & n22331 ;
  assign n11206 = n143 & n11205 ;
  assign n22522 = ~n10762 ;
  assign n11207 = n22522 & n11206 ;
  assign n22523 = ~n11206 ;
  assign n11208 = n10762 & n22523 ;
  assign n11209 = n11207 | n11208 ;
  assign n22524 = ~n11209 ;
  assign n11210 = n11204 & n22524 ;
  assign n11211 = n11203 | n11210 ;
  assign n11212 = x70 & n11211 ;
  assign n11213 = x70 | n11211 ;
  assign n11214 = n10765 & n22335 ;
  assign n11215 = n143 & n11214 ;
  assign n11216 = n10771 & n11215 ;
  assign n11217 = n10771 | n11215 ;
  assign n22525 = ~n11216 ;
  assign n11218 = n22525 & n11217 ;
  assign n22526 = ~n11218 ;
  assign n11219 = n11213 & n22526 ;
  assign n11220 = n11212 | n11219 ;
  assign n11221 = x71 & n11220 ;
  assign n11222 = x71 | n11220 ;
  assign n11223 = n10774 & n22339 ;
  assign n11224 = n143 & n11223 ;
  assign n11225 = n10780 & n11224 ;
  assign n11226 = n10780 | n11224 ;
  assign n22527 = ~n11225 ;
  assign n11227 = n22527 & n11226 ;
  assign n22528 = ~n11227 ;
  assign n11228 = n11222 & n22528 ;
  assign n11229 = n11221 | n11228 ;
  assign n11230 = x72 & n11229 ;
  assign n11231 = x72 | n11229 ;
  assign n11232 = n10783 & n22343 ;
  assign n11233 = n143 & n11232 ;
  assign n22529 = ~n10789 ;
  assign n11234 = n22529 & n11233 ;
  assign n22530 = ~n11233 ;
  assign n11235 = n10789 & n22530 ;
  assign n11236 = n11234 | n11235 ;
  assign n22531 = ~n11236 ;
  assign n11237 = n11231 & n22531 ;
  assign n11238 = n11230 | n11237 ;
  assign n11239 = x73 & n11238 ;
  assign n11240 = x73 | n11238 ;
  assign n11241 = n10792 & n22347 ;
  assign n11242 = n143 & n11241 ;
  assign n11243 = n10798 & n11242 ;
  assign n11244 = n10798 | n11242 ;
  assign n22532 = ~n11243 ;
  assign n11245 = n22532 & n11244 ;
  assign n22533 = ~n11245 ;
  assign n11246 = n11240 & n22533 ;
  assign n11247 = n11239 | n11246 ;
  assign n11248 = x74 & n11247 ;
  assign n11249 = x74 | n11247 ;
  assign n11250 = n10801 & n22351 ;
  assign n11251 = n143 & n11250 ;
  assign n22534 = ~n10807 ;
  assign n11252 = n22534 & n11251 ;
  assign n22535 = ~n11251 ;
  assign n11253 = n10807 & n22535 ;
  assign n11254 = n11252 | n11253 ;
  assign n22536 = ~n11254 ;
  assign n11255 = n11249 & n22536 ;
  assign n11256 = n11248 | n11255 ;
  assign n11257 = x75 & n11256 ;
  assign n11258 = x75 | n11256 ;
  assign n11259 = n10810 & n22355 ;
  assign n11260 = n143 & n11259 ;
  assign n22537 = ~n10816 ;
  assign n11261 = n22537 & n11260 ;
  assign n22538 = ~n11260 ;
  assign n11262 = n10816 & n22538 ;
  assign n11263 = n11261 | n11262 ;
  assign n22539 = ~n11263 ;
  assign n11264 = n11258 & n22539 ;
  assign n11265 = n11257 | n11264 ;
  assign n11266 = x76 & n11265 ;
  assign n11267 = x76 | n11265 ;
  assign n11268 = n10819 & n22359 ;
  assign n11269 = n143 & n11268 ;
  assign n11270 = n10825 & n11269 ;
  assign n11271 = n10825 | n11269 ;
  assign n22540 = ~n11270 ;
  assign n11272 = n22540 & n11271 ;
  assign n22541 = ~n11272 ;
  assign n11273 = n11267 & n22541 ;
  assign n11274 = n11266 | n11273 ;
  assign n11275 = x77 & n11274 ;
  assign n11276 = x77 | n11274 ;
  assign n11277 = n10828 & n22363 ;
  assign n11278 = n143 & n11277 ;
  assign n11279 = n10834 & n11278 ;
  assign n11280 = n10834 | n11278 ;
  assign n22542 = ~n11279 ;
  assign n11281 = n22542 & n11280 ;
  assign n22543 = ~n11281 ;
  assign n11282 = n11276 & n22543 ;
  assign n11283 = n11275 | n11282 ;
  assign n11284 = x78 & n11283 ;
  assign n11285 = x78 | n11283 ;
  assign n11286 = n10837 & n22367 ;
  assign n11287 = n143 & n11286 ;
  assign n22544 = ~n10843 ;
  assign n11288 = n22544 & n11287 ;
  assign n22545 = ~n11287 ;
  assign n11289 = n10843 & n22545 ;
  assign n11290 = n11288 | n11289 ;
  assign n22546 = ~n11290 ;
  assign n11291 = n11285 & n22546 ;
  assign n11292 = n11284 | n11291 ;
  assign n11293 = x79 & n11292 ;
  assign n11294 = x79 | n11292 ;
  assign n11295 = n10846 & n22371 ;
  assign n11296 = n143 & n11295 ;
  assign n11297 = n10852 & n11296 ;
  assign n11298 = n10852 | n11296 ;
  assign n22547 = ~n11297 ;
  assign n11299 = n22547 & n11298 ;
  assign n22548 = ~n11299 ;
  assign n11300 = n11294 & n22548 ;
  assign n11301 = n11293 | n11300 ;
  assign n11302 = x80 & n11301 ;
  assign n11303 = x80 | n11301 ;
  assign n11304 = n10855 & n22375 ;
  assign n11305 = n143 & n11304 ;
  assign n22549 = ~n10861 ;
  assign n11306 = n22549 & n11305 ;
  assign n22550 = ~n11305 ;
  assign n11307 = n10861 & n22550 ;
  assign n11308 = n11306 | n11307 ;
  assign n22551 = ~n11308 ;
  assign n11309 = n11303 & n22551 ;
  assign n11310 = n11302 | n11309 ;
  assign n11311 = x81 & n11310 ;
  assign n11312 = x81 | n11310 ;
  assign n11313 = n10864 & n22379 ;
  assign n11314 = n143 & n11313 ;
  assign n22552 = ~n10870 ;
  assign n11315 = n22552 & n11314 ;
  assign n22553 = ~n11314 ;
  assign n11316 = n10870 & n22553 ;
  assign n11317 = n11315 | n11316 ;
  assign n22554 = ~n11317 ;
  assign n11318 = n11312 & n22554 ;
  assign n11319 = n11311 | n11318 ;
  assign n11320 = x82 & n11319 ;
  assign n11321 = x82 | n11319 ;
  assign n11322 = n10873 & n22383 ;
  assign n11323 = n143 & n11322 ;
  assign n22555 = ~n10879 ;
  assign n11324 = n22555 & n11323 ;
  assign n22556 = ~n11323 ;
  assign n11325 = n10879 & n22556 ;
  assign n11326 = n11324 | n11325 ;
  assign n22557 = ~n11326 ;
  assign n11327 = n11321 & n22557 ;
  assign n11328 = n11320 | n11327 ;
  assign n11329 = x83 & n11328 ;
  assign n11330 = x83 | n11328 ;
  assign n11331 = n10882 & n22387 ;
  assign n11332 = n143 & n11331 ;
  assign n11333 = n10888 & n11332 ;
  assign n11334 = n10888 | n11332 ;
  assign n22558 = ~n11333 ;
  assign n11335 = n22558 & n11334 ;
  assign n22559 = ~n11335 ;
  assign n11336 = n11330 & n22559 ;
  assign n11337 = n11329 | n11336 ;
  assign n11338 = x84 & n11337 ;
  assign n11339 = x84 | n11337 ;
  assign n11340 = n10891 & n22391 ;
  assign n11341 = n143 & n11340 ;
  assign n11342 = n10897 & n11341 ;
  assign n11343 = n10897 | n11341 ;
  assign n22560 = ~n11342 ;
  assign n11344 = n22560 & n11343 ;
  assign n22561 = ~n11344 ;
  assign n11345 = n11339 & n22561 ;
  assign n11346 = n11338 | n11345 ;
  assign n11347 = x85 & n11346 ;
  assign n11348 = x85 | n11346 ;
  assign n11349 = n10900 & n22395 ;
  assign n11350 = n143 & n11349 ;
  assign n22562 = ~n10906 ;
  assign n11351 = n22562 & n11350 ;
  assign n22563 = ~n11350 ;
  assign n11352 = n10906 & n22563 ;
  assign n11353 = n11351 | n11352 ;
  assign n22564 = ~n11353 ;
  assign n11354 = n11348 & n22564 ;
  assign n11355 = n11347 | n11354 ;
  assign n11356 = x86 & n11355 ;
  assign n11357 = x86 | n11355 ;
  assign n11358 = n10909 & n22399 ;
  assign n11359 = n143 & n11358 ;
  assign n22565 = ~n10915 ;
  assign n11360 = n22565 & n11359 ;
  assign n22566 = ~n11359 ;
  assign n11361 = n10915 & n22566 ;
  assign n11362 = n11360 | n11361 ;
  assign n22567 = ~n11362 ;
  assign n11363 = n11357 & n22567 ;
  assign n11364 = n11356 | n11363 ;
  assign n11365 = x87 & n11364 ;
  assign n11366 = x87 | n11364 ;
  assign n11367 = n10918 & n22403 ;
  assign n11368 = n143 & n11367 ;
  assign n22568 = ~n10924 ;
  assign n11369 = n22568 & n11368 ;
  assign n22569 = ~n11368 ;
  assign n11370 = n10924 & n22569 ;
  assign n11371 = n11369 | n11370 ;
  assign n22570 = ~n11371 ;
  assign n11372 = n11366 & n22570 ;
  assign n11373 = n11365 | n11372 ;
  assign n11374 = x88 & n11373 ;
  assign n11375 = x88 | n11373 ;
  assign n11376 = n10927 & n22407 ;
  assign n11377 = n143 & n11376 ;
  assign n11378 = n10933 & n11377 ;
  assign n11379 = n10933 | n11377 ;
  assign n22571 = ~n11378 ;
  assign n11380 = n22571 & n11379 ;
  assign n22572 = ~n11380 ;
  assign n11381 = n11375 & n22572 ;
  assign n11382 = n11374 | n11381 ;
  assign n11383 = x89 & n11382 ;
  assign n11384 = x89 | n11382 ;
  assign n11385 = n10936 & n22411 ;
  assign n11386 = n143 & n11385 ;
  assign n22573 = ~n10942 ;
  assign n11387 = n22573 & n11386 ;
  assign n22574 = ~n11386 ;
  assign n11388 = n10942 & n22574 ;
  assign n11389 = n11387 | n11388 ;
  assign n22575 = ~n11389 ;
  assign n11390 = n11384 & n22575 ;
  assign n11391 = n11383 | n11390 ;
  assign n11392 = x90 & n11391 ;
  assign n11393 = x90 | n11391 ;
  assign n11394 = n10945 & n22415 ;
  assign n11395 = n143 & n11394 ;
  assign n11396 = n10951 & n11395 ;
  assign n11397 = n10951 | n11395 ;
  assign n22576 = ~n11396 ;
  assign n11398 = n22576 & n11397 ;
  assign n22577 = ~n11398 ;
  assign n11399 = n11393 & n22577 ;
  assign n11400 = n11392 | n11399 ;
  assign n11401 = x91 & n11400 ;
  assign n11402 = x91 | n11400 ;
  assign n11403 = n10954 & n22419 ;
  assign n11404 = n143 & n11403 ;
  assign n22578 = ~n10960 ;
  assign n11405 = n22578 & n11404 ;
  assign n22579 = ~n11404 ;
  assign n11406 = n10960 & n22579 ;
  assign n11407 = n11405 | n11406 ;
  assign n22580 = ~n11407 ;
  assign n11408 = n11402 & n22580 ;
  assign n11409 = n11401 | n11408 ;
  assign n11410 = x92 & n11409 ;
  assign n11411 = x92 | n11409 ;
  assign n11412 = n10963 & n22423 ;
  assign n11413 = n143 & n11412 ;
  assign n11414 = n10969 & n11413 ;
  assign n11415 = n10969 | n11413 ;
  assign n22581 = ~n11414 ;
  assign n11416 = n22581 & n11415 ;
  assign n22582 = ~n11416 ;
  assign n11417 = n11411 & n22582 ;
  assign n11418 = n11410 | n11417 ;
  assign n11419 = x93 & n11418 ;
  assign n11420 = x93 | n11418 ;
  assign n11421 = n10972 & n22427 ;
  assign n11422 = n143 & n11421 ;
  assign n11423 = n10978 & n11422 ;
  assign n11424 = n10978 | n11422 ;
  assign n22583 = ~n11423 ;
  assign n11425 = n22583 & n11424 ;
  assign n22584 = ~n11425 ;
  assign n11426 = n11420 & n22584 ;
  assign n11427 = n11419 | n11426 ;
  assign n11428 = x94 & n11427 ;
  assign n11429 = x94 | n11427 ;
  assign n11430 = n10981 & n22431 ;
  assign n11431 = n143 & n11430 ;
  assign n22585 = ~n10987 ;
  assign n11432 = n22585 & n11431 ;
  assign n22586 = ~n11431 ;
  assign n11433 = n10987 & n22586 ;
  assign n11434 = n11432 | n11433 ;
  assign n22587 = ~n11434 ;
  assign n11435 = n11429 & n22587 ;
  assign n11436 = n11428 | n11435 ;
  assign n11437 = x95 & n11436 ;
  assign n11438 = x95 | n11436 ;
  assign n11439 = n10990 & n22435 ;
  assign n11440 = n143 & n11439 ;
  assign n22588 = ~n10996 ;
  assign n11441 = n22588 & n11440 ;
  assign n22589 = ~n11440 ;
  assign n11442 = n10996 & n22589 ;
  assign n11443 = n11441 | n11442 ;
  assign n22590 = ~n11443 ;
  assign n11444 = n11438 & n22590 ;
  assign n11445 = n11437 | n11444 ;
  assign n11446 = x96 & n11445 ;
  assign n11447 = x96 | n11445 ;
  assign n11448 = n10999 & n22439 ;
  assign n11449 = n143 & n11448 ;
  assign n11450 = n11005 & n11449 ;
  assign n11451 = n11005 | n11449 ;
  assign n22591 = ~n11450 ;
  assign n11452 = n22591 & n11451 ;
  assign n22592 = ~n11452 ;
  assign n11453 = n11447 & n22592 ;
  assign n11454 = n11446 | n11453 ;
  assign n11455 = x97 & n11454 ;
  assign n11456 = x97 | n11454 ;
  assign n11457 = n11008 & n22443 ;
  assign n11458 = n143 & n11457 ;
  assign n11459 = n11014 & n11458 ;
  assign n11460 = n11014 | n11458 ;
  assign n22593 = ~n11459 ;
  assign n11461 = n22593 & n11460 ;
  assign n22594 = ~n11461 ;
  assign n11462 = n11456 & n22594 ;
  assign n11463 = n11455 | n11462 ;
  assign n11464 = x98 & n11463 ;
  assign n11465 = x98 | n11463 ;
  assign n11466 = n11017 & n22447 ;
  assign n11467 = n143 & n11466 ;
  assign n22595 = ~n11023 ;
  assign n11468 = n22595 & n11467 ;
  assign n22596 = ~n11467 ;
  assign n11469 = n11023 & n22596 ;
  assign n11470 = n11468 | n11469 ;
  assign n22597 = ~n11470 ;
  assign n11471 = n11465 & n22597 ;
  assign n11472 = n11464 | n11471 ;
  assign n11473 = x99 & n11472 ;
  assign n11474 = x99 | n11472 ;
  assign n11475 = n11026 & n22451 ;
  assign n11476 = n143 & n11475 ;
  assign n22598 = ~n11032 ;
  assign n11477 = n22598 & n11476 ;
  assign n22599 = ~n11476 ;
  assign n11478 = n11032 & n22599 ;
  assign n11479 = n11477 | n11478 ;
  assign n22600 = ~n11479 ;
  assign n11480 = n11474 & n22600 ;
  assign n11481 = n11473 | n11480 ;
  assign n11482 = x100 & n11481 ;
  assign n11483 = x100 | n11481 ;
  assign n11484 = n11035 & n22455 ;
  assign n11485 = n143 & n11484 ;
  assign n11486 = n11041 & n11485 ;
  assign n11487 = n11041 | n11485 ;
  assign n22601 = ~n11486 ;
  assign n11488 = n22601 & n11487 ;
  assign n22602 = ~n11488 ;
  assign n11489 = n11483 & n22602 ;
  assign n11490 = n11482 | n11489 ;
  assign n11491 = x101 & n11490 ;
  assign n11492 = x101 | n11490 ;
  assign n11493 = n11044 & n22459 ;
  assign n11494 = n143 & n11493 ;
  assign n22603 = ~n11050 ;
  assign n11495 = n22603 & n11494 ;
  assign n22604 = ~n11494 ;
  assign n11496 = n11050 & n22604 ;
  assign n11497 = n11495 | n11496 ;
  assign n22605 = ~n11497 ;
  assign n11498 = n11492 & n22605 ;
  assign n11499 = n11491 | n11498 ;
  assign n11500 = x102 & n11499 ;
  assign n11501 = x102 | n11499 ;
  assign n11502 = n11053 & n22463 ;
  assign n11503 = n143 & n11502 ;
  assign n22606 = ~n11059 ;
  assign n11504 = n22606 & n11503 ;
  assign n22607 = ~n11503 ;
  assign n11505 = n11059 & n22607 ;
  assign n11506 = n11504 | n11505 ;
  assign n22608 = ~n11506 ;
  assign n11507 = n11501 & n22608 ;
  assign n11508 = n11500 | n11507 ;
  assign n11509 = x103 & n11508 ;
  assign n11510 = x103 | n11508 ;
  assign n11511 = n11062 & n22467 ;
  assign n11512 = n143 & n11511 ;
  assign n11513 = n11068 & n11512 ;
  assign n11514 = n11068 | n11512 ;
  assign n22609 = ~n11513 ;
  assign n11515 = n22609 & n11514 ;
  assign n22610 = ~n11515 ;
  assign n11516 = n11510 & n22610 ;
  assign n11517 = n11509 | n11516 ;
  assign n11518 = x104 & n11517 ;
  assign n11519 = x104 | n11517 ;
  assign n11520 = n11071 & n22471 ;
  assign n11521 = n143 & n11520 ;
  assign n22611 = ~n11077 ;
  assign n11522 = n22611 & n11521 ;
  assign n22612 = ~n11521 ;
  assign n11523 = n11077 & n22612 ;
  assign n11524 = n11522 | n11523 ;
  assign n22613 = ~n11524 ;
  assign n11525 = n11519 & n22613 ;
  assign n11526 = n11518 | n11525 ;
  assign n11527 = x105 & n11526 ;
  assign n11528 = x105 | n11526 ;
  assign n11529 = n11080 & n22475 ;
  assign n11530 = n143 & n11529 ;
  assign n22614 = ~n11086 ;
  assign n11531 = n22614 & n11530 ;
  assign n22615 = ~n11530 ;
  assign n11532 = n11086 & n22615 ;
  assign n11533 = n11531 | n11532 ;
  assign n22616 = ~n11533 ;
  assign n11534 = n11528 & n22616 ;
  assign n11535 = n11527 | n11534 ;
  assign n11536 = x106 & n11535 ;
  assign n11537 = x106 | n11535 ;
  assign n11538 = n11089 & n22479 ;
  assign n11539 = n143 & n11538 ;
  assign n11540 = n11095 & n11539 ;
  assign n11541 = n11095 | n11539 ;
  assign n22617 = ~n11540 ;
  assign n11542 = n22617 & n11541 ;
  assign n22618 = ~n11542 ;
  assign n11543 = n11537 & n22618 ;
  assign n11544 = n11536 | n11543 ;
  assign n11545 = x107 & n11544 ;
  assign n11546 = x107 | n11544 ;
  assign n11547 = n11098 & n22483 ;
  assign n11548 = n143 & n11547 ;
  assign n22619 = ~n11104 ;
  assign n11549 = n22619 & n11548 ;
  assign n22620 = ~n11548 ;
  assign n11550 = n11104 & n22620 ;
  assign n11551 = n11549 | n11550 ;
  assign n22621 = ~n11551 ;
  assign n11552 = n11546 & n22621 ;
  assign n11553 = n11545 | n11552 ;
  assign n11554 = x108 & n11553 ;
  assign n11555 = x108 | n11553 ;
  assign n11556 = n11107 & n22487 ;
  assign n11557 = n143 & n11556 ;
  assign n22622 = ~n11113 ;
  assign n11558 = n22622 & n11557 ;
  assign n22623 = ~n11557 ;
  assign n11559 = n11113 & n22623 ;
  assign n11560 = n11558 | n11559 ;
  assign n22624 = ~n11560 ;
  assign n11561 = n11555 & n22624 ;
  assign n11562 = n11554 | n11561 ;
  assign n11563 = x109 & n11562 ;
  assign n11564 = x109 | n11562 ;
  assign n11565 = n11116 & n22491 ;
  assign n11566 = n143 & n11565 ;
  assign n22625 = ~n11122 ;
  assign n11567 = n22625 & n11566 ;
  assign n22626 = ~n11566 ;
  assign n11568 = n11122 & n22626 ;
  assign n11569 = n11567 | n11568 ;
  assign n22627 = ~n11569 ;
  assign n11570 = n11564 & n22627 ;
  assign n11571 = n11563 | n11570 ;
  assign n11572 = x110 & n11571 ;
  assign n11573 = x110 | n11571 ;
  assign n11574 = n11125 & n22495 ;
  assign n11575 = n143 & n11574 ;
  assign n22628 = ~n11131 ;
  assign n11576 = n22628 & n11575 ;
  assign n22629 = ~n11575 ;
  assign n11577 = n11131 & n22629 ;
  assign n11578 = n11576 | n11577 ;
  assign n22630 = ~n11578 ;
  assign n11579 = n11573 & n22630 ;
  assign n11580 = n11572 | n11579 ;
  assign n11581 = x111 & n11580 ;
  assign n11582 = x111 | n11580 ;
  assign n11583 = n11134 & n22499 ;
  assign n11584 = n143 & n11583 ;
  assign n11585 = n11140 & n11584 ;
  assign n11586 = n11140 | n11584 ;
  assign n22631 = ~n11585 ;
  assign n11587 = n22631 & n11586 ;
  assign n22632 = ~n11587 ;
  assign n11588 = n11582 & n22632 ;
  assign n11589 = n11581 | n11588 ;
  assign n11590 = x112 & n11589 ;
  assign n11591 = x112 | n11589 ;
  assign n11592 = n11143 & n22503 ;
  assign n11593 = n143 & n11592 ;
  assign n22633 = ~n11149 ;
  assign n11594 = n22633 & n11593 ;
  assign n22634 = ~n11593 ;
  assign n11595 = n11149 & n22634 ;
  assign n11596 = n11594 | n11595 ;
  assign n22635 = ~n11596 ;
  assign n11597 = n11591 & n22635 ;
  assign n11598 = n11590 | n11597 ;
  assign n11599 = x113 & n11598 ;
  assign n11600 = x113 | n11598 ;
  assign n22636 = ~n11166 ;
  assign n11601 = n22636 & n11600 ;
  assign n11602 = n11599 | n11601 ;
  assign n11604 = x114 & n11602 ;
  assign n11605 = n18323 | n11604 ;
  assign n11603 = x114 | n11602 ;
  assign n11606 = n18333 & n10712 ;
  assign n11607 = n11160 & n11606 ;
  assign n11608 = n21884 | n11607 ;
  assign n22637 = ~n11608 ;
  assign n11609 = n11603 & n22637 ;
  assign n11610 = n11605 | n11609 ;
  assign n22638 = ~n11599 ;
  assign n11611 = n22638 & n11600 ;
  assign n142 = ~n11610 ;
  assign n11612 = n142 & n11611 ;
  assign n11613 = n22636 & n11612 ;
  assign n22640 = ~n11612 ;
  assign n11614 = n11166 & n22640 ;
  assign n11615 = n11613 | n11614 ;
  assign n22641 = ~x12 ;
  assign n11616 = n22641 & x64 ;
  assign n11618 = x65 | n11616 ;
  assign n11617 = x65 & n11616 ;
  assign n11619 = x64 & n142 ;
  assign n11620 = x13 & n11619 ;
  assign n11621 = x13 | n11619 ;
  assign n22642 = ~n11620 ;
  assign n11622 = n22642 & n11621 ;
  assign n22643 = ~n11617 ;
  assign n11623 = n22643 & n11622 ;
  assign n22644 = ~n11623 ;
  assign n11624 = n11618 & n22644 ;
  assign n11625 = x66 | n11624 ;
  assign n11626 = x66 & n11624 ;
  assign n11627 = n11168 & n142 ;
  assign n11628 = n22513 & n11627 ;
  assign n11629 = n11172 | n11628 ;
  assign n11630 = n11174 & n11627 ;
  assign n22645 = ~n11630 ;
  assign n11631 = n11629 & n22645 ;
  assign n22646 = ~n11626 ;
  assign n11632 = n22646 & n11631 ;
  assign n22647 = ~n11632 ;
  assign n11633 = n11625 & n22647 ;
  assign n11634 = x67 | n11633 ;
  assign n11635 = x67 & n11633 ;
  assign n22648 = ~n11176 ;
  assign n11636 = n22648 & n11182 ;
  assign n11637 = n142 & n11636 ;
  assign n11638 = n11181 & n11637 ;
  assign n11639 = n11181 | n11637 ;
  assign n22649 = ~n11638 ;
  assign n11640 = n22649 & n11639 ;
  assign n22650 = ~n11635 ;
  assign n11641 = n22650 & n11640 ;
  assign n22651 = ~n11641 ;
  assign n11642 = n11634 & n22651 ;
  assign n11643 = x68 | n11642 ;
  assign n11644 = x68 & n11642 ;
  assign n22652 = ~n11185 ;
  assign n11645 = n22652 & n11186 ;
  assign n11646 = n142 & n11645 ;
  assign n11647 = n11191 & n11646 ;
  assign n11648 = n11191 | n11646 ;
  assign n22653 = ~n11647 ;
  assign n11649 = n22653 & n11648 ;
  assign n22654 = ~n11644 ;
  assign n11650 = n22654 & n11649 ;
  assign n22655 = ~n11650 ;
  assign n11651 = n11643 & n22655 ;
  assign n11652 = x69 | n11651 ;
  assign n11653 = x69 & n11651 ;
  assign n22656 = ~n11194 ;
  assign n11654 = n22656 & n11195 ;
  assign n11655 = n142 & n11654 ;
  assign n11656 = n22521 & n11655 ;
  assign n22657 = ~n11655 ;
  assign n11657 = n11200 & n22657 ;
  assign n11658 = n11656 | n11657 ;
  assign n22658 = ~n11653 ;
  assign n11659 = n22658 & n11658 ;
  assign n22659 = ~n11659 ;
  assign n11660 = n11652 & n22659 ;
  assign n11661 = x70 | n11660 ;
  assign n11662 = x70 & n11660 ;
  assign n22660 = ~n11203 ;
  assign n11663 = n22660 & n11204 ;
  assign n11664 = n142 & n11663 ;
  assign n11665 = n11209 & n11664 ;
  assign n11666 = n11209 | n11664 ;
  assign n22661 = ~n11665 ;
  assign n11667 = n22661 & n11666 ;
  assign n22662 = ~n11662 ;
  assign n11668 = n22662 & n11667 ;
  assign n22663 = ~n11668 ;
  assign n11669 = n11661 & n22663 ;
  assign n11670 = x71 | n11669 ;
  assign n11671 = x71 & n11669 ;
  assign n22664 = ~n11212 ;
  assign n11672 = n22664 & n11213 ;
  assign n11673 = n142 & n11672 ;
  assign n11674 = n11218 & n11673 ;
  assign n11675 = n11218 | n11673 ;
  assign n22665 = ~n11674 ;
  assign n11676 = n22665 & n11675 ;
  assign n22666 = ~n11671 ;
  assign n11677 = n22666 & n11676 ;
  assign n22667 = ~n11677 ;
  assign n11678 = n11670 & n22667 ;
  assign n11679 = x72 | n11678 ;
  assign n11680 = x72 & n11678 ;
  assign n22668 = ~n11221 ;
  assign n11681 = n22668 & n11222 ;
  assign n11682 = n142 & n11681 ;
  assign n11683 = n11227 & n11682 ;
  assign n11684 = n11227 | n11682 ;
  assign n22669 = ~n11683 ;
  assign n11685 = n22669 & n11684 ;
  assign n22670 = ~n11680 ;
  assign n11686 = n22670 & n11685 ;
  assign n22671 = ~n11686 ;
  assign n11687 = n11679 & n22671 ;
  assign n11688 = x73 | n11687 ;
  assign n11689 = x73 & n11687 ;
  assign n22672 = ~n11230 ;
  assign n11690 = n22672 & n11231 ;
  assign n11691 = n142 & n11690 ;
  assign n11692 = n22531 & n11691 ;
  assign n22673 = ~n11691 ;
  assign n11693 = n11236 & n22673 ;
  assign n11694 = n11692 | n11693 ;
  assign n22674 = ~n11689 ;
  assign n11695 = n22674 & n11694 ;
  assign n22675 = ~n11695 ;
  assign n11696 = n11688 & n22675 ;
  assign n11697 = x74 | n11696 ;
  assign n11698 = x74 & n11696 ;
  assign n22676 = ~n11239 ;
  assign n11699 = n22676 & n11240 ;
  assign n11700 = n142 & n11699 ;
  assign n11701 = n11245 & n11700 ;
  assign n11702 = n11245 | n11700 ;
  assign n22677 = ~n11701 ;
  assign n11703 = n22677 & n11702 ;
  assign n22678 = ~n11698 ;
  assign n11704 = n22678 & n11703 ;
  assign n22679 = ~n11704 ;
  assign n11705 = n11697 & n22679 ;
  assign n11706 = x75 | n11705 ;
  assign n11707 = x75 & n11705 ;
  assign n22680 = ~n11248 ;
  assign n11708 = n22680 & n11249 ;
  assign n11709 = n142 & n11708 ;
  assign n11710 = n22536 & n11709 ;
  assign n22681 = ~n11709 ;
  assign n11711 = n11254 & n22681 ;
  assign n11712 = n11710 | n11711 ;
  assign n22682 = ~n11707 ;
  assign n11713 = n22682 & n11712 ;
  assign n22683 = ~n11713 ;
  assign n11714 = n11706 & n22683 ;
  assign n11715 = x76 | n11714 ;
  assign n11716 = x76 & n11714 ;
  assign n22684 = ~n11257 ;
  assign n11717 = n22684 & n11258 ;
  assign n11718 = n142 & n11717 ;
  assign n11719 = n11263 & n11718 ;
  assign n11720 = n11263 | n11718 ;
  assign n22685 = ~n11719 ;
  assign n11721 = n22685 & n11720 ;
  assign n22686 = ~n11716 ;
  assign n11722 = n22686 & n11721 ;
  assign n22687 = ~n11722 ;
  assign n11723 = n11715 & n22687 ;
  assign n11724 = x77 | n11723 ;
  assign n11725 = x77 & n11723 ;
  assign n22688 = ~n11266 ;
  assign n11726 = n22688 & n11267 ;
  assign n11727 = n142 & n11726 ;
  assign n11728 = n11272 & n11727 ;
  assign n11729 = n11272 | n11727 ;
  assign n22689 = ~n11728 ;
  assign n11730 = n22689 & n11729 ;
  assign n22690 = ~n11725 ;
  assign n11731 = n22690 & n11730 ;
  assign n22691 = ~n11731 ;
  assign n11732 = n11724 & n22691 ;
  assign n11733 = x78 | n11732 ;
  assign n11734 = x78 & n11732 ;
  assign n22692 = ~n11275 ;
  assign n11735 = n22692 & n11276 ;
  assign n11736 = n142 & n11735 ;
  assign n11737 = n11281 & n11736 ;
  assign n11738 = n11281 | n11736 ;
  assign n22693 = ~n11737 ;
  assign n11739 = n22693 & n11738 ;
  assign n22694 = ~n11734 ;
  assign n11740 = n22694 & n11739 ;
  assign n22695 = ~n11740 ;
  assign n11741 = n11733 & n22695 ;
  assign n11742 = x79 | n11741 ;
  assign n11743 = x79 & n11741 ;
  assign n22696 = ~n11284 ;
  assign n11744 = n22696 & n11285 ;
  assign n11745 = n142 & n11744 ;
  assign n11746 = n11290 & n11745 ;
  assign n11747 = n11290 | n11745 ;
  assign n22697 = ~n11746 ;
  assign n11748 = n22697 & n11747 ;
  assign n22698 = ~n11743 ;
  assign n11749 = n22698 & n11748 ;
  assign n22699 = ~n11749 ;
  assign n11750 = n11742 & n22699 ;
  assign n11751 = x80 | n11750 ;
  assign n11752 = x80 & n11750 ;
  assign n22700 = ~n11293 ;
  assign n11753 = n22700 & n11294 ;
  assign n11754 = n142 & n11753 ;
  assign n11755 = n11299 & n11754 ;
  assign n11756 = n11299 | n11754 ;
  assign n22701 = ~n11755 ;
  assign n11757 = n22701 & n11756 ;
  assign n22702 = ~n11752 ;
  assign n11758 = n22702 & n11757 ;
  assign n22703 = ~n11758 ;
  assign n11759 = n11751 & n22703 ;
  assign n11760 = x81 | n11759 ;
  assign n11761 = x81 & n11759 ;
  assign n22704 = ~n11302 ;
  assign n11762 = n22704 & n11303 ;
  assign n11763 = n142 & n11762 ;
  assign n11764 = n11308 & n11763 ;
  assign n11765 = n11308 | n11763 ;
  assign n22705 = ~n11764 ;
  assign n11766 = n22705 & n11765 ;
  assign n22706 = ~n11761 ;
  assign n11767 = n22706 & n11766 ;
  assign n22707 = ~n11767 ;
  assign n11768 = n11760 & n22707 ;
  assign n11769 = x82 | n11768 ;
  assign n11770 = x82 & n11768 ;
  assign n22708 = ~n11311 ;
  assign n11771 = n22708 & n11312 ;
  assign n11772 = n142 & n11771 ;
  assign n11773 = n11317 & n11772 ;
  assign n11774 = n11317 | n11772 ;
  assign n22709 = ~n11773 ;
  assign n11775 = n22709 & n11774 ;
  assign n22710 = ~n11770 ;
  assign n11776 = n22710 & n11775 ;
  assign n22711 = ~n11776 ;
  assign n11777 = n11769 & n22711 ;
  assign n11778 = x83 | n11777 ;
  assign n11779 = x83 & n11777 ;
  assign n22712 = ~n11320 ;
  assign n11780 = n22712 & n11321 ;
  assign n11781 = n142 & n11780 ;
  assign n11782 = n22557 & n11781 ;
  assign n22713 = ~n11781 ;
  assign n11783 = n11326 & n22713 ;
  assign n11784 = n11782 | n11783 ;
  assign n22714 = ~n11779 ;
  assign n11785 = n22714 & n11784 ;
  assign n22715 = ~n11785 ;
  assign n11786 = n11778 & n22715 ;
  assign n11787 = x84 | n11786 ;
  assign n11788 = x84 & n11786 ;
  assign n22716 = ~n11329 ;
  assign n11789 = n22716 & n11330 ;
  assign n11790 = n142 & n11789 ;
  assign n11791 = n11335 & n11790 ;
  assign n11792 = n11335 | n11790 ;
  assign n22717 = ~n11791 ;
  assign n11793 = n22717 & n11792 ;
  assign n22718 = ~n11788 ;
  assign n11794 = n22718 & n11793 ;
  assign n22719 = ~n11794 ;
  assign n11795 = n11787 & n22719 ;
  assign n11796 = x85 | n11795 ;
  assign n11797 = x85 & n11795 ;
  assign n22720 = ~n11338 ;
  assign n11798 = n22720 & n11339 ;
  assign n11799 = n142 & n11798 ;
  assign n11800 = n11344 & n11799 ;
  assign n11801 = n11344 | n11799 ;
  assign n22721 = ~n11800 ;
  assign n11802 = n22721 & n11801 ;
  assign n22722 = ~n11797 ;
  assign n11803 = n22722 & n11802 ;
  assign n22723 = ~n11803 ;
  assign n11804 = n11796 & n22723 ;
  assign n11805 = x86 | n11804 ;
  assign n11806 = x86 & n11804 ;
  assign n22724 = ~n11347 ;
  assign n11807 = n22724 & n11348 ;
  assign n11808 = n142 & n11807 ;
  assign n11809 = n11353 & n11808 ;
  assign n11810 = n11353 | n11808 ;
  assign n22725 = ~n11809 ;
  assign n11811 = n22725 & n11810 ;
  assign n22726 = ~n11806 ;
  assign n11812 = n22726 & n11811 ;
  assign n22727 = ~n11812 ;
  assign n11813 = n11805 & n22727 ;
  assign n11814 = x87 | n11813 ;
  assign n11815 = x87 & n11813 ;
  assign n22728 = ~n11356 ;
  assign n11816 = n22728 & n11357 ;
  assign n11817 = n142 & n11816 ;
  assign n11818 = n11362 & n11817 ;
  assign n11819 = n11362 | n11817 ;
  assign n22729 = ~n11818 ;
  assign n11820 = n22729 & n11819 ;
  assign n22730 = ~n11815 ;
  assign n11821 = n22730 & n11820 ;
  assign n22731 = ~n11821 ;
  assign n11822 = n11814 & n22731 ;
  assign n11823 = x88 | n11822 ;
  assign n11824 = x88 & n11822 ;
  assign n22732 = ~n11365 ;
  assign n11825 = n22732 & n11366 ;
  assign n11826 = n142 & n11825 ;
  assign n11827 = n22570 & n11826 ;
  assign n22733 = ~n11826 ;
  assign n11828 = n11371 & n22733 ;
  assign n11829 = n11827 | n11828 ;
  assign n22734 = ~n11824 ;
  assign n11830 = n22734 & n11829 ;
  assign n22735 = ~n11830 ;
  assign n11831 = n11823 & n22735 ;
  assign n11832 = x89 | n11831 ;
  assign n11833 = x89 & n11831 ;
  assign n22736 = ~n11374 ;
  assign n11834 = n22736 & n11375 ;
  assign n11835 = n142 & n11834 ;
  assign n11836 = n11380 & n11835 ;
  assign n11837 = n11380 | n11835 ;
  assign n22737 = ~n11836 ;
  assign n11838 = n22737 & n11837 ;
  assign n22738 = ~n11833 ;
  assign n11839 = n22738 & n11838 ;
  assign n22739 = ~n11839 ;
  assign n11840 = n11832 & n22739 ;
  assign n11841 = x90 | n11840 ;
  assign n11842 = x90 & n11840 ;
  assign n22740 = ~n11383 ;
  assign n11843 = n22740 & n11384 ;
  assign n11844 = n142 & n11843 ;
  assign n11845 = n22575 & n11844 ;
  assign n22741 = ~n11844 ;
  assign n11846 = n11389 & n22741 ;
  assign n11847 = n11845 | n11846 ;
  assign n22742 = ~n11842 ;
  assign n11848 = n22742 & n11847 ;
  assign n22743 = ~n11848 ;
  assign n11849 = n11841 & n22743 ;
  assign n11850 = x91 | n11849 ;
  assign n11851 = x91 & n11849 ;
  assign n22744 = ~n11392 ;
  assign n11852 = n22744 & n11393 ;
  assign n11853 = n142 & n11852 ;
  assign n11854 = n11398 & n11853 ;
  assign n11855 = n11398 | n11853 ;
  assign n22745 = ~n11854 ;
  assign n11856 = n22745 & n11855 ;
  assign n22746 = ~n11851 ;
  assign n11857 = n22746 & n11856 ;
  assign n22747 = ~n11857 ;
  assign n11858 = n11850 & n22747 ;
  assign n11859 = x92 | n11858 ;
  assign n11860 = x92 & n11858 ;
  assign n22748 = ~n11401 ;
  assign n11861 = n22748 & n11402 ;
  assign n11862 = n142 & n11861 ;
  assign n11863 = n22580 & n11862 ;
  assign n22749 = ~n11862 ;
  assign n11864 = n11407 & n22749 ;
  assign n11865 = n11863 | n11864 ;
  assign n22750 = ~n11860 ;
  assign n11866 = n22750 & n11865 ;
  assign n22751 = ~n11866 ;
  assign n11867 = n11859 & n22751 ;
  assign n11868 = x93 | n11867 ;
  assign n11869 = x93 & n11867 ;
  assign n22752 = ~n11410 ;
  assign n11870 = n22752 & n11411 ;
  assign n11871 = n142 & n11870 ;
  assign n11872 = n11416 & n11871 ;
  assign n11873 = n11416 | n11871 ;
  assign n22753 = ~n11872 ;
  assign n11874 = n22753 & n11873 ;
  assign n22754 = ~n11869 ;
  assign n11875 = n22754 & n11874 ;
  assign n22755 = ~n11875 ;
  assign n11876 = n11868 & n22755 ;
  assign n11877 = x94 | n11876 ;
  assign n11878 = x94 & n11876 ;
  assign n22756 = ~n11419 ;
  assign n11879 = n22756 & n11420 ;
  assign n11880 = n142 & n11879 ;
  assign n11881 = n11425 & n11880 ;
  assign n11882 = n11425 | n11880 ;
  assign n22757 = ~n11881 ;
  assign n11883 = n22757 & n11882 ;
  assign n22758 = ~n11878 ;
  assign n11884 = n22758 & n11883 ;
  assign n22759 = ~n11884 ;
  assign n11885 = n11877 & n22759 ;
  assign n11886 = x95 | n11885 ;
  assign n11887 = x95 & n11885 ;
  assign n22760 = ~n11428 ;
  assign n11888 = n22760 & n11429 ;
  assign n11889 = n142 & n11888 ;
  assign n11890 = n11434 & n11889 ;
  assign n11891 = n11434 | n11889 ;
  assign n22761 = ~n11890 ;
  assign n11892 = n22761 & n11891 ;
  assign n22762 = ~n11887 ;
  assign n11893 = n22762 & n11892 ;
  assign n22763 = ~n11893 ;
  assign n11894 = n11886 & n22763 ;
  assign n11895 = x96 | n11894 ;
  assign n11896 = x96 & n11894 ;
  assign n22764 = ~n11437 ;
  assign n11897 = n22764 & n11438 ;
  assign n11898 = n142 & n11897 ;
  assign n11899 = n11443 & n11898 ;
  assign n11900 = n11443 | n11898 ;
  assign n22765 = ~n11899 ;
  assign n11901 = n22765 & n11900 ;
  assign n22766 = ~n11896 ;
  assign n11902 = n22766 & n11901 ;
  assign n22767 = ~n11902 ;
  assign n11903 = n11895 & n22767 ;
  assign n11904 = x97 | n11903 ;
  assign n11905 = x97 & n11903 ;
  assign n22768 = ~n11446 ;
  assign n11906 = n22768 & n11447 ;
  assign n11907 = n142 & n11906 ;
  assign n11908 = n11452 & n11907 ;
  assign n11909 = n11452 | n11907 ;
  assign n22769 = ~n11908 ;
  assign n11910 = n22769 & n11909 ;
  assign n22770 = ~n11905 ;
  assign n11911 = n22770 & n11910 ;
  assign n22771 = ~n11911 ;
  assign n11912 = n11904 & n22771 ;
  assign n11913 = x98 | n11912 ;
  assign n11914 = x98 & n11912 ;
  assign n22772 = ~n11455 ;
  assign n11915 = n22772 & n11456 ;
  assign n11916 = n142 & n11915 ;
  assign n11917 = n11461 & n11916 ;
  assign n11918 = n11461 | n11916 ;
  assign n22773 = ~n11917 ;
  assign n11919 = n22773 & n11918 ;
  assign n22774 = ~n11914 ;
  assign n11920 = n22774 & n11919 ;
  assign n22775 = ~n11920 ;
  assign n11921 = n11913 & n22775 ;
  assign n11922 = x99 | n11921 ;
  assign n11923 = x99 & n11921 ;
  assign n22776 = ~n11464 ;
  assign n11924 = n22776 & n11465 ;
  assign n11925 = n142 & n11924 ;
  assign n11926 = n22597 & n11925 ;
  assign n22777 = ~n11925 ;
  assign n11927 = n11470 & n22777 ;
  assign n11928 = n11926 | n11927 ;
  assign n22778 = ~n11923 ;
  assign n11929 = n22778 & n11928 ;
  assign n22779 = ~n11929 ;
  assign n11930 = n11922 & n22779 ;
  assign n11931 = x100 | n11930 ;
  assign n11932 = x100 & n11930 ;
  assign n22780 = ~n11473 ;
  assign n11933 = n22780 & n11474 ;
  assign n11934 = n142 & n11933 ;
  assign n11935 = n11479 & n11934 ;
  assign n11936 = n11479 | n11934 ;
  assign n22781 = ~n11935 ;
  assign n11937 = n22781 & n11936 ;
  assign n22782 = ~n11932 ;
  assign n11938 = n22782 & n11937 ;
  assign n22783 = ~n11938 ;
  assign n11939 = n11931 & n22783 ;
  assign n11940 = x101 | n11939 ;
  assign n11941 = x101 & n11939 ;
  assign n22784 = ~n11482 ;
  assign n11942 = n22784 & n11483 ;
  assign n11943 = n142 & n11942 ;
  assign n11944 = n11488 & n11943 ;
  assign n11945 = n11488 | n11943 ;
  assign n22785 = ~n11944 ;
  assign n11946 = n22785 & n11945 ;
  assign n22786 = ~n11941 ;
  assign n11947 = n22786 & n11946 ;
  assign n22787 = ~n11947 ;
  assign n11948 = n11940 & n22787 ;
  assign n11949 = x102 | n11948 ;
  assign n11950 = x102 & n11948 ;
  assign n22788 = ~n11491 ;
  assign n11951 = n22788 & n11492 ;
  assign n11952 = n142 & n11951 ;
  assign n11953 = n22605 & n11952 ;
  assign n22789 = ~n11952 ;
  assign n11954 = n11497 & n22789 ;
  assign n11955 = n11953 | n11954 ;
  assign n22790 = ~n11950 ;
  assign n11956 = n22790 & n11955 ;
  assign n22791 = ~n11956 ;
  assign n11957 = n11949 & n22791 ;
  assign n11958 = x103 | n11957 ;
  assign n11959 = x103 & n11957 ;
  assign n22792 = ~n11500 ;
  assign n11960 = n22792 & n11501 ;
  assign n11961 = n142 & n11960 ;
  assign n11962 = n11506 & n11961 ;
  assign n11963 = n11506 | n11961 ;
  assign n22793 = ~n11962 ;
  assign n11964 = n22793 & n11963 ;
  assign n22794 = ~n11959 ;
  assign n11965 = n22794 & n11964 ;
  assign n22795 = ~n11965 ;
  assign n11966 = n11958 & n22795 ;
  assign n11967 = x104 | n11966 ;
  assign n11968 = x104 & n11966 ;
  assign n22796 = ~n11509 ;
  assign n11969 = n22796 & n11510 ;
  assign n11970 = n142 & n11969 ;
  assign n11971 = n11515 & n11970 ;
  assign n11972 = n11515 | n11970 ;
  assign n22797 = ~n11971 ;
  assign n11973 = n22797 & n11972 ;
  assign n22798 = ~n11968 ;
  assign n11974 = n22798 & n11973 ;
  assign n22799 = ~n11974 ;
  assign n11975 = n11967 & n22799 ;
  assign n11976 = x105 | n11975 ;
  assign n11977 = x105 & n11975 ;
  assign n22800 = ~n11518 ;
  assign n11978 = n22800 & n11519 ;
  assign n11979 = n142 & n11978 ;
  assign n11980 = n22613 & n11979 ;
  assign n22801 = ~n11979 ;
  assign n11981 = n11524 & n22801 ;
  assign n11982 = n11980 | n11981 ;
  assign n22802 = ~n11977 ;
  assign n11983 = n22802 & n11982 ;
  assign n22803 = ~n11983 ;
  assign n11984 = n11976 & n22803 ;
  assign n11985 = x106 | n11984 ;
  assign n11986 = x106 & n11984 ;
  assign n22804 = ~n11527 ;
  assign n11987 = n22804 & n11528 ;
  assign n11988 = n142 & n11987 ;
  assign n11989 = n22616 & n11988 ;
  assign n22805 = ~n11988 ;
  assign n11990 = n11533 & n22805 ;
  assign n11991 = n11989 | n11990 ;
  assign n22806 = ~n11986 ;
  assign n11992 = n22806 & n11991 ;
  assign n22807 = ~n11992 ;
  assign n11993 = n11985 & n22807 ;
  assign n11994 = x107 | n11993 ;
  assign n11995 = x107 & n11993 ;
  assign n22808 = ~n11536 ;
  assign n11996 = n22808 & n11537 ;
  assign n11997 = n142 & n11996 ;
  assign n11998 = n11542 & n11997 ;
  assign n11999 = n11542 | n11997 ;
  assign n22809 = ~n11998 ;
  assign n12000 = n22809 & n11999 ;
  assign n22810 = ~n11995 ;
  assign n12001 = n22810 & n12000 ;
  assign n22811 = ~n12001 ;
  assign n12002 = n11994 & n22811 ;
  assign n12003 = x108 | n12002 ;
  assign n12004 = x108 & n12002 ;
  assign n22812 = ~n11545 ;
  assign n12005 = n22812 & n11546 ;
  assign n12006 = n142 & n12005 ;
  assign n12007 = n22621 & n12006 ;
  assign n22813 = ~n12006 ;
  assign n12008 = n11551 & n22813 ;
  assign n12009 = n12007 | n12008 ;
  assign n22814 = ~n12004 ;
  assign n12010 = n22814 & n12009 ;
  assign n22815 = ~n12010 ;
  assign n12011 = n12003 & n22815 ;
  assign n12012 = x109 | n12011 ;
  assign n12013 = x109 & n12011 ;
  assign n22816 = ~n11554 ;
  assign n12014 = n22816 & n11555 ;
  assign n12015 = n142 & n12014 ;
  assign n12016 = n11560 & n12015 ;
  assign n12017 = n11560 | n12015 ;
  assign n22817 = ~n12016 ;
  assign n12018 = n22817 & n12017 ;
  assign n22818 = ~n12013 ;
  assign n12019 = n22818 & n12018 ;
  assign n22819 = ~n12019 ;
  assign n12020 = n12012 & n22819 ;
  assign n12021 = x110 | n12020 ;
  assign n12022 = x110 & n12020 ;
  assign n22820 = ~n11563 ;
  assign n12023 = n22820 & n11564 ;
  assign n12024 = n142 & n12023 ;
  assign n12025 = n11569 & n12024 ;
  assign n12026 = n11569 | n12024 ;
  assign n22821 = ~n12025 ;
  assign n12027 = n22821 & n12026 ;
  assign n22822 = ~n12022 ;
  assign n12028 = n22822 & n12027 ;
  assign n22823 = ~n12028 ;
  assign n12029 = n12021 & n22823 ;
  assign n12030 = x111 | n12029 ;
  assign n12031 = x111 & n12029 ;
  assign n22824 = ~n11572 ;
  assign n12032 = n22824 & n11573 ;
  assign n12033 = n142 & n12032 ;
  assign n12034 = n11578 & n12033 ;
  assign n12035 = n11578 | n12033 ;
  assign n22825 = ~n12034 ;
  assign n12036 = n22825 & n12035 ;
  assign n22826 = ~n12031 ;
  assign n12037 = n22826 & n12036 ;
  assign n22827 = ~n12037 ;
  assign n12038 = n12030 & n22827 ;
  assign n12039 = x112 | n12038 ;
  assign n12040 = x112 & n12038 ;
  assign n22828 = ~n11581 ;
  assign n12041 = n22828 & n11582 ;
  assign n12042 = n142 & n12041 ;
  assign n12043 = n11587 & n12042 ;
  assign n12044 = n11587 | n12042 ;
  assign n22829 = ~n12043 ;
  assign n12045 = n22829 & n12044 ;
  assign n22830 = ~n12040 ;
  assign n12046 = n22830 & n12045 ;
  assign n22831 = ~n12046 ;
  assign n12047 = n12039 & n22831 ;
  assign n12048 = x113 | n12047 ;
  assign n12049 = x113 & n12047 ;
  assign n22832 = ~n11590 ;
  assign n12050 = n22832 & n11591 ;
  assign n12051 = n142 & n12050 ;
  assign n12052 = n11596 & n12051 ;
  assign n12053 = n11596 | n12051 ;
  assign n22833 = ~n12052 ;
  assign n12054 = n22833 & n12053 ;
  assign n22834 = ~n12049 ;
  assign n12055 = n22834 & n12054 ;
  assign n22835 = ~n12055 ;
  assign n12056 = n12048 & n22835 ;
  assign n12057 = x114 | n12056 ;
  assign n12058 = x114 & n12056 ;
  assign n22836 = ~n12058 ;
  assign n12059 = n11615 & n22836 ;
  assign n22837 = ~n12059 ;
  assign n12060 = n12057 & n22837 ;
  assign n22838 = ~n11605 ;
  assign n12061 = n11603 & n22838 ;
  assign n22839 = ~n12061 ;
  assign n12062 = n11608 & n22839 ;
  assign n22840 = ~x115 ;
  assign n12063 = n22840 & n12062 ;
  assign n22841 = ~n12063 ;
  assign n12064 = n12060 & n22841 ;
  assign n22842 = ~n12062 ;
  assign n12065 = x115 & n22842 ;
  assign n12066 = n18318 | n12065 ;
  assign n12067 = n12064 | n12066 ;
  assign n12068 = n12057 & n22836 ;
  assign n141 = ~n12067 ;
  assign n12069 = n141 & n12068 ;
  assign n12070 = n11615 & n12069 ;
  assign n12071 = n11615 | n12069 ;
  assign n22844 = ~n12070 ;
  assign n12072 = n22844 & n12071 ;
  assign n12073 = x115 & n12060 ;
  assign n12074 = x115 | n12060 ;
  assign n22845 = ~n18318 ;
  assign n12075 = n22845 & n12074 ;
  assign n22846 = ~n12073 ;
  assign n12076 = n22846 & n12075 ;
  assign n22847 = ~n12076 ;
  assign n12077 = n12062 & n22847 ;
  assign n12078 = n22845 & n12077 ;
  assign n22848 = ~x11 ;
  assign n12079 = n22848 & x64 ;
  assign n12080 = x65 | n12079 ;
  assign n12081 = x65 & n12079 ;
  assign n12082 = x64 & n141 ;
  assign n12083 = x12 & n12082 ;
  assign n12084 = x12 | n12082 ;
  assign n22849 = ~n12083 ;
  assign n12085 = n22849 & n12084 ;
  assign n22850 = ~n12081 ;
  assign n12086 = n22850 & n12085 ;
  assign n22851 = ~n12086 ;
  assign n12087 = n12080 & n22851 ;
  assign n12089 = x66 | n12087 ;
  assign n12088 = x66 & n12087 ;
  assign n12090 = n22643 & n11618 ;
  assign n12091 = n141 & n12090 ;
  assign n12092 = n11622 & n12091 ;
  assign n12093 = n11622 | n12091 ;
  assign n22852 = ~n12092 ;
  assign n12094 = n22852 & n12093 ;
  assign n22853 = ~n12088 ;
  assign n12095 = n22853 & n12094 ;
  assign n22854 = ~n12095 ;
  assign n12096 = n12089 & n22854 ;
  assign n12097 = x67 | n12096 ;
  assign n12098 = x67 & n12096 ;
  assign n12099 = n11625 & n22646 ;
  assign n12100 = n141 & n12099 ;
  assign n22855 = ~n11631 ;
  assign n12101 = n22855 & n12100 ;
  assign n22856 = ~n12100 ;
  assign n12102 = n11631 & n22856 ;
  assign n12103 = n12101 | n12102 ;
  assign n22857 = ~n12098 ;
  assign n12104 = n22857 & n12103 ;
  assign n22858 = ~n12104 ;
  assign n12105 = n12097 & n22858 ;
  assign n12106 = x68 | n12105 ;
  assign n12107 = x68 & n12105 ;
  assign n12108 = n11634 & n22650 ;
  assign n12109 = n141 & n12108 ;
  assign n22859 = ~n11640 ;
  assign n12110 = n22859 & n12109 ;
  assign n22860 = ~n12109 ;
  assign n12111 = n11640 & n22860 ;
  assign n12112 = n12110 | n12111 ;
  assign n22861 = ~n12107 ;
  assign n12113 = n22861 & n12112 ;
  assign n22862 = ~n12113 ;
  assign n12114 = n12106 & n22862 ;
  assign n12115 = x69 | n12114 ;
  assign n12116 = x69 & n12114 ;
  assign n12117 = n11643 & n22654 ;
  assign n12118 = n141 & n12117 ;
  assign n22863 = ~n11649 ;
  assign n12119 = n22863 & n12118 ;
  assign n22864 = ~n12118 ;
  assign n12120 = n11649 & n22864 ;
  assign n12121 = n12119 | n12120 ;
  assign n22865 = ~n12116 ;
  assign n12122 = n22865 & n12121 ;
  assign n22866 = ~n12122 ;
  assign n12123 = n12115 & n22866 ;
  assign n12124 = x70 | n12123 ;
  assign n12125 = x70 & n12123 ;
  assign n12126 = n11652 & n22658 ;
  assign n12127 = n141 & n12126 ;
  assign n22867 = ~n11658 ;
  assign n12128 = n22867 & n12127 ;
  assign n22868 = ~n12127 ;
  assign n12129 = n11658 & n22868 ;
  assign n12130 = n12128 | n12129 ;
  assign n22869 = ~n12125 ;
  assign n12131 = n22869 & n12130 ;
  assign n22870 = ~n12131 ;
  assign n12132 = n12124 & n22870 ;
  assign n12133 = x71 | n12132 ;
  assign n12134 = x71 & n12132 ;
  assign n12135 = n11661 & n22662 ;
  assign n12136 = n141 & n12135 ;
  assign n12137 = n11667 & n12136 ;
  assign n12138 = n11667 | n12136 ;
  assign n22871 = ~n12137 ;
  assign n12139 = n22871 & n12138 ;
  assign n22872 = ~n12134 ;
  assign n12140 = n22872 & n12139 ;
  assign n22873 = ~n12140 ;
  assign n12141 = n12133 & n22873 ;
  assign n12142 = x72 | n12141 ;
  assign n12143 = x72 & n12141 ;
  assign n12144 = n11670 & n22666 ;
  assign n12145 = n141 & n12144 ;
  assign n22874 = ~n11676 ;
  assign n12146 = n22874 & n12145 ;
  assign n22875 = ~n12145 ;
  assign n12147 = n11676 & n22875 ;
  assign n12148 = n12146 | n12147 ;
  assign n22876 = ~n12143 ;
  assign n12149 = n22876 & n12148 ;
  assign n22877 = ~n12149 ;
  assign n12150 = n12142 & n22877 ;
  assign n12151 = x73 | n12150 ;
  assign n12152 = x73 & n12150 ;
  assign n12153 = n11679 & n22670 ;
  assign n12154 = n141 & n12153 ;
  assign n22878 = ~n11685 ;
  assign n12155 = n22878 & n12154 ;
  assign n22879 = ~n12154 ;
  assign n12156 = n11685 & n22879 ;
  assign n12157 = n12155 | n12156 ;
  assign n22880 = ~n12152 ;
  assign n12158 = n22880 & n12157 ;
  assign n22881 = ~n12158 ;
  assign n12159 = n12151 & n22881 ;
  assign n12160 = x74 | n12159 ;
  assign n12161 = x74 & n12159 ;
  assign n12162 = n11688 & n22674 ;
  assign n12163 = n141 & n12162 ;
  assign n22882 = ~n11694 ;
  assign n12164 = n22882 & n12163 ;
  assign n22883 = ~n12163 ;
  assign n12165 = n11694 & n22883 ;
  assign n12166 = n12164 | n12165 ;
  assign n22884 = ~n12161 ;
  assign n12167 = n22884 & n12166 ;
  assign n22885 = ~n12167 ;
  assign n12168 = n12160 & n22885 ;
  assign n12169 = x75 | n12168 ;
  assign n12170 = x75 & n12168 ;
  assign n12171 = n11697 & n22678 ;
  assign n12172 = n141 & n12171 ;
  assign n22886 = ~n11703 ;
  assign n12173 = n22886 & n12172 ;
  assign n22887 = ~n12172 ;
  assign n12174 = n11703 & n22887 ;
  assign n12175 = n12173 | n12174 ;
  assign n22888 = ~n12170 ;
  assign n12176 = n22888 & n12175 ;
  assign n22889 = ~n12176 ;
  assign n12177 = n12169 & n22889 ;
  assign n12178 = x76 | n12177 ;
  assign n12179 = x76 & n12177 ;
  assign n12180 = n11706 & n22682 ;
  assign n12181 = n141 & n12180 ;
  assign n22890 = ~n11712 ;
  assign n12182 = n22890 & n12181 ;
  assign n22891 = ~n12181 ;
  assign n12183 = n11712 & n22891 ;
  assign n12184 = n12182 | n12183 ;
  assign n22892 = ~n12179 ;
  assign n12185 = n22892 & n12184 ;
  assign n22893 = ~n12185 ;
  assign n12186 = n12178 & n22893 ;
  assign n12187 = x77 | n12186 ;
  assign n12188 = x77 & n12186 ;
  assign n12189 = n11715 & n22686 ;
  assign n12190 = n141 & n12189 ;
  assign n12191 = n11721 & n12190 ;
  assign n12192 = n11721 | n12190 ;
  assign n22894 = ~n12191 ;
  assign n12193 = n22894 & n12192 ;
  assign n22895 = ~n12188 ;
  assign n12194 = n22895 & n12193 ;
  assign n22896 = ~n12194 ;
  assign n12195 = n12187 & n22896 ;
  assign n12196 = x78 | n12195 ;
  assign n12197 = x78 & n12195 ;
  assign n12198 = n11724 & n22690 ;
  assign n12199 = n141 & n12198 ;
  assign n22897 = ~n11730 ;
  assign n12200 = n22897 & n12199 ;
  assign n22898 = ~n12199 ;
  assign n12201 = n11730 & n22898 ;
  assign n12202 = n12200 | n12201 ;
  assign n22899 = ~n12197 ;
  assign n12203 = n22899 & n12202 ;
  assign n22900 = ~n12203 ;
  assign n12204 = n12196 & n22900 ;
  assign n12205 = x79 | n12204 ;
  assign n12206 = x79 & n12204 ;
  assign n12207 = n11733 & n22694 ;
  assign n12208 = n141 & n12207 ;
  assign n22901 = ~n11739 ;
  assign n12209 = n22901 & n12208 ;
  assign n22902 = ~n12208 ;
  assign n12210 = n11739 & n22902 ;
  assign n12211 = n12209 | n12210 ;
  assign n22903 = ~n12206 ;
  assign n12212 = n22903 & n12211 ;
  assign n22904 = ~n12212 ;
  assign n12213 = n12205 & n22904 ;
  assign n12214 = x80 | n12213 ;
  assign n12215 = x80 & n12213 ;
  assign n12216 = n11742 & n22698 ;
  assign n12217 = n141 & n12216 ;
  assign n12218 = n11748 & n12217 ;
  assign n12219 = n11748 | n12217 ;
  assign n22905 = ~n12218 ;
  assign n12220 = n22905 & n12219 ;
  assign n22906 = ~n12215 ;
  assign n12221 = n22906 & n12220 ;
  assign n22907 = ~n12221 ;
  assign n12222 = n12214 & n22907 ;
  assign n12223 = x81 | n12222 ;
  assign n12224 = x81 & n12222 ;
  assign n12225 = n11751 & n22702 ;
  assign n12226 = n141 & n12225 ;
  assign n22908 = ~n11757 ;
  assign n12227 = n22908 & n12226 ;
  assign n22909 = ~n12226 ;
  assign n12228 = n11757 & n22909 ;
  assign n12229 = n12227 | n12228 ;
  assign n22910 = ~n12224 ;
  assign n12230 = n22910 & n12229 ;
  assign n22911 = ~n12230 ;
  assign n12231 = n12223 & n22911 ;
  assign n12232 = x82 | n12231 ;
  assign n12233 = x82 & n12231 ;
  assign n12234 = n11760 & n22706 ;
  assign n12235 = n141 & n12234 ;
  assign n12236 = n11766 & n12235 ;
  assign n12237 = n11766 | n12235 ;
  assign n22912 = ~n12236 ;
  assign n12238 = n22912 & n12237 ;
  assign n22913 = ~n12233 ;
  assign n12239 = n22913 & n12238 ;
  assign n22914 = ~n12239 ;
  assign n12240 = n12232 & n22914 ;
  assign n12241 = x83 | n12240 ;
  assign n12242 = x83 & n12240 ;
  assign n12243 = n11769 & n22710 ;
  assign n12244 = n141 & n12243 ;
  assign n12245 = n11775 & n12244 ;
  assign n12246 = n11775 | n12244 ;
  assign n22915 = ~n12245 ;
  assign n12247 = n22915 & n12246 ;
  assign n22916 = ~n12242 ;
  assign n12248 = n22916 & n12247 ;
  assign n22917 = ~n12248 ;
  assign n12249 = n12241 & n22917 ;
  assign n12250 = x84 | n12249 ;
  assign n12251 = x84 & n12249 ;
  assign n12252 = n11778 & n22714 ;
  assign n12253 = n141 & n12252 ;
  assign n22918 = ~n11784 ;
  assign n12254 = n22918 & n12253 ;
  assign n22919 = ~n12253 ;
  assign n12255 = n11784 & n22919 ;
  assign n12256 = n12254 | n12255 ;
  assign n22920 = ~n12251 ;
  assign n12257 = n22920 & n12256 ;
  assign n22921 = ~n12257 ;
  assign n12258 = n12250 & n22921 ;
  assign n12259 = x85 | n12258 ;
  assign n12260 = x85 & n12258 ;
  assign n12261 = n11787 & n22718 ;
  assign n12262 = n141 & n12261 ;
  assign n22922 = ~n11793 ;
  assign n12263 = n22922 & n12262 ;
  assign n22923 = ~n12262 ;
  assign n12264 = n11793 & n22923 ;
  assign n12265 = n12263 | n12264 ;
  assign n22924 = ~n12260 ;
  assign n12266 = n22924 & n12265 ;
  assign n22925 = ~n12266 ;
  assign n12267 = n12259 & n22925 ;
  assign n12268 = x86 | n12267 ;
  assign n12269 = x86 & n12267 ;
  assign n12270 = n11796 & n22722 ;
  assign n12271 = n141 & n12270 ;
  assign n12272 = n11802 & n12271 ;
  assign n12273 = n11802 | n12271 ;
  assign n22926 = ~n12272 ;
  assign n12274 = n22926 & n12273 ;
  assign n22927 = ~n12269 ;
  assign n12275 = n22927 & n12274 ;
  assign n22928 = ~n12275 ;
  assign n12276 = n12268 & n22928 ;
  assign n12277 = x87 | n12276 ;
  assign n12278 = x87 & n12276 ;
  assign n12279 = n11805 & n22726 ;
  assign n12280 = n141 & n12279 ;
  assign n12281 = n11811 & n12280 ;
  assign n12282 = n11811 | n12280 ;
  assign n22929 = ~n12281 ;
  assign n12283 = n22929 & n12282 ;
  assign n22930 = ~n12278 ;
  assign n12284 = n22930 & n12283 ;
  assign n22931 = ~n12284 ;
  assign n12285 = n12277 & n22931 ;
  assign n12286 = x88 | n12285 ;
  assign n12287 = x88 & n12285 ;
  assign n12288 = n11814 & n22730 ;
  assign n12289 = n141 & n12288 ;
  assign n12290 = n11820 & n12289 ;
  assign n12291 = n11820 | n12289 ;
  assign n22932 = ~n12290 ;
  assign n12292 = n22932 & n12291 ;
  assign n22933 = ~n12287 ;
  assign n12293 = n22933 & n12292 ;
  assign n22934 = ~n12293 ;
  assign n12294 = n12286 & n22934 ;
  assign n12295 = x89 | n12294 ;
  assign n12296 = x89 & n12294 ;
  assign n12297 = n11823 & n22734 ;
  assign n12298 = n141 & n12297 ;
  assign n22935 = ~n11829 ;
  assign n12299 = n22935 & n12298 ;
  assign n22936 = ~n12298 ;
  assign n12300 = n11829 & n22936 ;
  assign n12301 = n12299 | n12300 ;
  assign n22937 = ~n12296 ;
  assign n12302 = n22937 & n12301 ;
  assign n22938 = ~n12302 ;
  assign n12303 = n12295 & n22938 ;
  assign n12304 = x90 | n12303 ;
  assign n12305 = x90 & n12303 ;
  assign n12306 = n11832 & n22738 ;
  assign n12307 = n141 & n12306 ;
  assign n22939 = ~n11838 ;
  assign n12308 = n22939 & n12307 ;
  assign n22940 = ~n12307 ;
  assign n12309 = n11838 & n22940 ;
  assign n12310 = n12308 | n12309 ;
  assign n22941 = ~n12305 ;
  assign n12311 = n22941 & n12310 ;
  assign n22942 = ~n12311 ;
  assign n12312 = n12304 & n22942 ;
  assign n12313 = x91 | n12312 ;
  assign n12314 = x91 & n12312 ;
  assign n12315 = n11841 & n22742 ;
  assign n12316 = n141 & n12315 ;
  assign n22943 = ~n11847 ;
  assign n12317 = n22943 & n12316 ;
  assign n22944 = ~n12316 ;
  assign n12318 = n11847 & n22944 ;
  assign n12319 = n12317 | n12318 ;
  assign n22945 = ~n12314 ;
  assign n12320 = n22945 & n12319 ;
  assign n22946 = ~n12320 ;
  assign n12321 = n12313 & n22946 ;
  assign n12322 = x92 | n12321 ;
  assign n12323 = x92 & n12321 ;
  assign n12324 = n11850 & n22746 ;
  assign n12325 = n141 & n12324 ;
  assign n22947 = ~n11856 ;
  assign n12326 = n22947 & n12325 ;
  assign n22948 = ~n12325 ;
  assign n12327 = n11856 & n22948 ;
  assign n12328 = n12326 | n12327 ;
  assign n22949 = ~n12323 ;
  assign n12329 = n22949 & n12328 ;
  assign n22950 = ~n12329 ;
  assign n12330 = n12322 & n22950 ;
  assign n12331 = x93 | n12330 ;
  assign n12332 = x93 & n12330 ;
  assign n12333 = n11859 & n22750 ;
  assign n12334 = n141 & n12333 ;
  assign n22951 = ~n11865 ;
  assign n12335 = n22951 & n12334 ;
  assign n22952 = ~n12334 ;
  assign n12336 = n11865 & n22952 ;
  assign n12337 = n12335 | n12336 ;
  assign n22953 = ~n12332 ;
  assign n12338 = n22953 & n12337 ;
  assign n22954 = ~n12338 ;
  assign n12339 = n12331 & n22954 ;
  assign n12340 = x94 | n12339 ;
  assign n12341 = x94 & n12339 ;
  assign n12342 = n11868 & n22754 ;
  assign n12343 = n141 & n12342 ;
  assign n22955 = ~n11874 ;
  assign n12344 = n22955 & n12343 ;
  assign n22956 = ~n12343 ;
  assign n12345 = n11874 & n22956 ;
  assign n12346 = n12344 | n12345 ;
  assign n22957 = ~n12341 ;
  assign n12347 = n22957 & n12346 ;
  assign n22958 = ~n12347 ;
  assign n12348 = n12340 & n22958 ;
  assign n12349 = x95 | n12348 ;
  assign n12350 = x95 & n12348 ;
  assign n12351 = n11877 & n22758 ;
  assign n12352 = n141 & n12351 ;
  assign n22959 = ~n11883 ;
  assign n12353 = n22959 & n12352 ;
  assign n22960 = ~n12352 ;
  assign n12354 = n11883 & n22960 ;
  assign n12355 = n12353 | n12354 ;
  assign n22961 = ~n12350 ;
  assign n12356 = n22961 & n12355 ;
  assign n22962 = ~n12356 ;
  assign n12357 = n12349 & n22962 ;
  assign n12358 = x96 | n12357 ;
  assign n12359 = x96 & n12357 ;
  assign n12360 = n11886 & n22762 ;
  assign n12361 = n141 & n12360 ;
  assign n12362 = n11892 & n12361 ;
  assign n12363 = n11892 | n12361 ;
  assign n22963 = ~n12362 ;
  assign n12364 = n22963 & n12363 ;
  assign n22964 = ~n12359 ;
  assign n12365 = n22964 & n12364 ;
  assign n22965 = ~n12365 ;
  assign n12366 = n12358 & n22965 ;
  assign n12367 = x97 | n12366 ;
  assign n12368 = x97 & n12366 ;
  assign n12369 = n11895 & n22766 ;
  assign n12370 = n141 & n12369 ;
  assign n12371 = n11901 & n12370 ;
  assign n12372 = n11901 | n12370 ;
  assign n22966 = ~n12371 ;
  assign n12373 = n22966 & n12372 ;
  assign n22967 = ~n12368 ;
  assign n12374 = n22967 & n12373 ;
  assign n22968 = ~n12374 ;
  assign n12375 = n12367 & n22968 ;
  assign n12376 = x98 | n12375 ;
  assign n12377 = x98 & n12375 ;
  assign n12378 = n11904 & n22770 ;
  assign n12379 = n141 & n12378 ;
  assign n22969 = ~n11910 ;
  assign n12380 = n22969 & n12379 ;
  assign n22970 = ~n12379 ;
  assign n12381 = n11910 & n22970 ;
  assign n12382 = n12380 | n12381 ;
  assign n22971 = ~n12377 ;
  assign n12383 = n22971 & n12382 ;
  assign n22972 = ~n12383 ;
  assign n12384 = n12376 & n22972 ;
  assign n12385 = x99 | n12384 ;
  assign n12386 = x99 & n12384 ;
  assign n12387 = n11913 & n22774 ;
  assign n12388 = n141 & n12387 ;
  assign n22973 = ~n11919 ;
  assign n12389 = n22973 & n12388 ;
  assign n22974 = ~n12388 ;
  assign n12390 = n11919 & n22974 ;
  assign n12391 = n12389 | n12390 ;
  assign n22975 = ~n12386 ;
  assign n12392 = n22975 & n12391 ;
  assign n22976 = ~n12392 ;
  assign n12393 = n12385 & n22976 ;
  assign n12394 = x100 | n12393 ;
  assign n12395 = x100 & n12393 ;
  assign n12396 = n11922 & n22778 ;
  assign n12397 = n141 & n12396 ;
  assign n22977 = ~n11928 ;
  assign n12398 = n22977 & n12397 ;
  assign n22978 = ~n12397 ;
  assign n12399 = n11928 & n22978 ;
  assign n12400 = n12398 | n12399 ;
  assign n22979 = ~n12395 ;
  assign n12401 = n22979 & n12400 ;
  assign n22980 = ~n12401 ;
  assign n12402 = n12394 & n22980 ;
  assign n12403 = x101 | n12402 ;
  assign n12404 = x101 & n12402 ;
  assign n12405 = n11931 & n22782 ;
  assign n12406 = n141 & n12405 ;
  assign n12407 = n11937 & n12406 ;
  assign n12408 = n11937 | n12406 ;
  assign n22981 = ~n12407 ;
  assign n12409 = n22981 & n12408 ;
  assign n22982 = ~n12404 ;
  assign n12410 = n22982 & n12409 ;
  assign n22983 = ~n12410 ;
  assign n12411 = n12403 & n22983 ;
  assign n12412 = x102 | n12411 ;
  assign n12413 = x102 & n12411 ;
  assign n12414 = n11940 & n22786 ;
  assign n12415 = n141 & n12414 ;
  assign n22984 = ~n11946 ;
  assign n12416 = n22984 & n12415 ;
  assign n22985 = ~n12415 ;
  assign n12417 = n11946 & n22985 ;
  assign n12418 = n12416 | n12417 ;
  assign n22986 = ~n12413 ;
  assign n12419 = n22986 & n12418 ;
  assign n22987 = ~n12419 ;
  assign n12420 = n12412 & n22987 ;
  assign n12421 = x103 | n12420 ;
  assign n12422 = x103 & n12420 ;
  assign n12423 = n11949 & n22790 ;
  assign n12424 = n141 & n12423 ;
  assign n22988 = ~n11955 ;
  assign n12425 = n22988 & n12424 ;
  assign n22989 = ~n12424 ;
  assign n12426 = n11955 & n22989 ;
  assign n12427 = n12425 | n12426 ;
  assign n22990 = ~n12422 ;
  assign n12428 = n22990 & n12427 ;
  assign n22991 = ~n12428 ;
  assign n12429 = n12421 & n22991 ;
  assign n12430 = x104 | n12429 ;
  assign n12431 = x104 & n12429 ;
  assign n12432 = n11958 & n22794 ;
  assign n12433 = n141 & n12432 ;
  assign n12434 = n11964 & n12433 ;
  assign n12435 = n11964 | n12433 ;
  assign n22992 = ~n12434 ;
  assign n12436 = n22992 & n12435 ;
  assign n22993 = ~n12431 ;
  assign n12437 = n22993 & n12436 ;
  assign n22994 = ~n12437 ;
  assign n12438 = n12430 & n22994 ;
  assign n12439 = x105 | n12438 ;
  assign n12440 = x105 & n12438 ;
  assign n12441 = n11967 & n22798 ;
  assign n12442 = n141 & n12441 ;
  assign n22995 = ~n11973 ;
  assign n12443 = n22995 & n12442 ;
  assign n22996 = ~n12442 ;
  assign n12444 = n11973 & n22996 ;
  assign n12445 = n12443 | n12444 ;
  assign n22997 = ~n12440 ;
  assign n12446 = n22997 & n12445 ;
  assign n22998 = ~n12446 ;
  assign n12447 = n12439 & n22998 ;
  assign n12448 = x106 | n12447 ;
  assign n12449 = x106 & n12447 ;
  assign n12450 = n11976 & n22802 ;
  assign n12451 = n141 & n12450 ;
  assign n22999 = ~n11982 ;
  assign n12452 = n22999 & n12451 ;
  assign n23000 = ~n12451 ;
  assign n12453 = n11982 & n23000 ;
  assign n12454 = n12452 | n12453 ;
  assign n23001 = ~n12449 ;
  assign n12455 = n23001 & n12454 ;
  assign n23002 = ~n12455 ;
  assign n12456 = n12448 & n23002 ;
  assign n12457 = x107 | n12456 ;
  assign n12458 = x107 & n12456 ;
  assign n12459 = n11985 & n22806 ;
  assign n12460 = n141 & n12459 ;
  assign n23003 = ~n11991 ;
  assign n12461 = n23003 & n12460 ;
  assign n23004 = ~n12460 ;
  assign n12462 = n11991 & n23004 ;
  assign n12463 = n12461 | n12462 ;
  assign n23005 = ~n12458 ;
  assign n12464 = n23005 & n12463 ;
  assign n23006 = ~n12464 ;
  assign n12465 = n12457 & n23006 ;
  assign n12466 = x108 | n12465 ;
  assign n12467 = x108 & n12465 ;
  assign n12468 = n11994 & n22810 ;
  assign n12469 = n141 & n12468 ;
  assign n23007 = ~n12000 ;
  assign n12470 = n23007 & n12469 ;
  assign n23008 = ~n12469 ;
  assign n12471 = n12000 & n23008 ;
  assign n12472 = n12470 | n12471 ;
  assign n23009 = ~n12467 ;
  assign n12473 = n23009 & n12472 ;
  assign n23010 = ~n12473 ;
  assign n12474 = n12466 & n23010 ;
  assign n12475 = x109 | n12474 ;
  assign n12476 = x109 & n12474 ;
  assign n12477 = n12003 & n22814 ;
  assign n12478 = n141 & n12477 ;
  assign n23011 = ~n12009 ;
  assign n12479 = n23011 & n12478 ;
  assign n23012 = ~n12478 ;
  assign n12480 = n12009 & n23012 ;
  assign n12481 = n12479 | n12480 ;
  assign n23013 = ~n12476 ;
  assign n12482 = n23013 & n12481 ;
  assign n23014 = ~n12482 ;
  assign n12483 = n12475 & n23014 ;
  assign n12484 = x110 | n12483 ;
  assign n12485 = x110 & n12483 ;
  assign n12486 = n12012 & n22818 ;
  assign n12487 = n141 & n12486 ;
  assign n12488 = n12018 & n12487 ;
  assign n12489 = n12018 | n12487 ;
  assign n23015 = ~n12488 ;
  assign n12490 = n23015 & n12489 ;
  assign n23016 = ~n12485 ;
  assign n12491 = n23016 & n12490 ;
  assign n23017 = ~n12491 ;
  assign n12492 = n12484 & n23017 ;
  assign n12493 = x111 | n12492 ;
  assign n12494 = x111 & n12492 ;
  assign n12495 = n12021 & n22822 ;
  assign n12496 = n141 & n12495 ;
  assign n12497 = n12027 & n12496 ;
  assign n12498 = n12027 | n12496 ;
  assign n23018 = ~n12497 ;
  assign n12499 = n23018 & n12498 ;
  assign n23019 = ~n12494 ;
  assign n12500 = n23019 & n12499 ;
  assign n23020 = ~n12500 ;
  assign n12501 = n12493 & n23020 ;
  assign n12502 = x112 | n12501 ;
  assign n12503 = x112 & n12501 ;
  assign n12504 = n12030 & n22826 ;
  assign n12505 = n141 & n12504 ;
  assign n12506 = n12036 & n12505 ;
  assign n12507 = n12036 | n12505 ;
  assign n23021 = ~n12506 ;
  assign n12508 = n23021 & n12507 ;
  assign n23022 = ~n12503 ;
  assign n12509 = n23022 & n12508 ;
  assign n23023 = ~n12509 ;
  assign n12510 = n12502 & n23023 ;
  assign n12511 = x113 | n12510 ;
  assign n12512 = x113 & n12510 ;
  assign n12513 = n12039 & n22830 ;
  assign n12514 = n141 & n12513 ;
  assign n23024 = ~n12045 ;
  assign n12515 = n23024 & n12514 ;
  assign n23025 = ~n12514 ;
  assign n12516 = n12045 & n23025 ;
  assign n12517 = n12515 | n12516 ;
  assign n23026 = ~n12512 ;
  assign n12518 = n23026 & n12517 ;
  assign n23027 = ~n12518 ;
  assign n12519 = n12511 & n23027 ;
  assign n12520 = x114 | n12519 ;
  assign n12521 = x114 & n12519 ;
  assign n12522 = n12048 & n22834 ;
  assign n12523 = n141 & n12522 ;
  assign n12524 = n12054 & n12523 ;
  assign n12525 = n12054 | n12523 ;
  assign n23028 = ~n12524 ;
  assign n12526 = n23028 & n12525 ;
  assign n23029 = ~n12521 ;
  assign n12527 = n23029 & n12526 ;
  assign n23030 = ~n12527 ;
  assign n12528 = n12520 & n23030 ;
  assign n12530 = x115 | n12528 ;
  assign n23031 = ~n12072 ;
  assign n12531 = n23031 & n12530 ;
  assign n12529 = x115 & n12528 ;
  assign n12532 = x116 & n22842 ;
  assign n12533 = n18313 | n12532 ;
  assign n23032 = ~x116 ;
  assign n12534 = n23032 & n12077 ;
  assign n12535 = n12533 | n12534 ;
  assign n12536 = n12529 | n12535 ;
  assign n12537 = n12531 | n12536 ;
  assign n23033 = ~n12078 ;
  assign n12538 = n23033 & n12537 ;
  assign n23034 = ~n12529 ;
  assign n12539 = n23034 & n12530 ;
  assign n140 = ~n12538 ;
  assign n12540 = n140 & n12539 ;
  assign n12541 = n12072 & n12540 ;
  assign n12542 = n12072 | n12540 ;
  assign n23036 = ~n12541 ;
  assign n12543 = n23036 & n12542 ;
  assign n23037 = ~x10 ;
  assign n12544 = n23037 & x64 ;
  assign n12545 = x65 | n12544 ;
  assign n12546 = x64 & n140 ;
  assign n23038 = ~n12546 ;
  assign n12547 = x11 & n23038 ;
  assign n12548 = n12079 & n140 ;
  assign n12549 = n12547 | n12548 ;
  assign n12550 = x65 & n12544 ;
  assign n23039 = ~n12550 ;
  assign n12551 = n12549 & n23039 ;
  assign n23040 = ~n12551 ;
  assign n12552 = n12545 & n23040 ;
  assign n12554 = x66 & n12552 ;
  assign n12553 = x66 | n12552 ;
  assign n12555 = n12080 & n22850 ;
  assign n12556 = n140 & n12555 ;
  assign n12557 = n12085 & n12556 ;
  assign n12558 = n12085 | n12556 ;
  assign n23041 = ~n12557 ;
  assign n12559 = n23041 & n12558 ;
  assign n23042 = ~n12559 ;
  assign n12560 = n12553 & n23042 ;
  assign n12561 = n12554 | n12560 ;
  assign n12562 = x67 & n12561 ;
  assign n12563 = x67 | n12561 ;
  assign n12564 = n12089 & n140 ;
  assign n12565 = n12095 & n12564 ;
  assign n12566 = n22853 & n12564 ;
  assign n12567 = n12094 | n12566 ;
  assign n23043 = ~n12565 ;
  assign n12568 = n23043 & n12567 ;
  assign n23044 = ~n12568 ;
  assign n12569 = n12563 & n23044 ;
  assign n12570 = n12562 | n12569 ;
  assign n12571 = x68 & n12570 ;
  assign n12572 = x68 | n12570 ;
  assign n12573 = n12097 & n140 ;
  assign n12574 = n12104 & n12573 ;
  assign n12575 = n22857 & n12573 ;
  assign n12576 = n12103 | n12575 ;
  assign n23045 = ~n12574 ;
  assign n12577 = n23045 & n12576 ;
  assign n23046 = ~n12577 ;
  assign n12578 = n12572 & n23046 ;
  assign n12579 = n12571 | n12578 ;
  assign n12580 = x69 & n12579 ;
  assign n12581 = x69 | n12579 ;
  assign n12582 = n12106 & n22861 ;
  assign n12583 = n140 & n12582 ;
  assign n23047 = ~n12112 ;
  assign n12584 = n23047 & n12583 ;
  assign n23048 = ~n12583 ;
  assign n12585 = n12112 & n23048 ;
  assign n12586 = n12584 | n12585 ;
  assign n23049 = ~n12586 ;
  assign n12587 = n12581 & n23049 ;
  assign n12588 = n12580 | n12587 ;
  assign n12589 = x70 & n12588 ;
  assign n12590 = x70 | n12588 ;
  assign n12591 = n12115 & n22865 ;
  assign n12592 = n140 & n12591 ;
  assign n23050 = ~n12121 ;
  assign n12593 = n23050 & n12592 ;
  assign n23051 = ~n12592 ;
  assign n12594 = n12121 & n23051 ;
  assign n12595 = n12593 | n12594 ;
  assign n23052 = ~n12595 ;
  assign n12596 = n12590 & n23052 ;
  assign n12597 = n12589 | n12596 ;
  assign n12598 = x71 & n12597 ;
  assign n12599 = x71 | n12597 ;
  assign n12600 = n12124 & n22869 ;
  assign n12601 = n140 & n12600 ;
  assign n23053 = ~n12130 ;
  assign n12602 = n23053 & n12601 ;
  assign n23054 = ~n12601 ;
  assign n12603 = n12130 & n23054 ;
  assign n12604 = n12602 | n12603 ;
  assign n23055 = ~n12604 ;
  assign n12605 = n12599 & n23055 ;
  assign n12606 = n12598 | n12605 ;
  assign n12607 = x72 & n12606 ;
  assign n12608 = x72 | n12606 ;
  assign n12609 = n12133 & n22872 ;
  assign n12610 = n140 & n12609 ;
  assign n23056 = ~n12139 ;
  assign n12611 = n23056 & n12610 ;
  assign n23057 = ~n12610 ;
  assign n12612 = n12139 & n23057 ;
  assign n12613 = n12611 | n12612 ;
  assign n23058 = ~n12613 ;
  assign n12614 = n12608 & n23058 ;
  assign n12615 = n12607 | n12614 ;
  assign n12616 = x73 & n12615 ;
  assign n12617 = x73 | n12615 ;
  assign n12618 = n12142 & n22876 ;
  assign n12619 = n140 & n12618 ;
  assign n23059 = ~n12148 ;
  assign n12620 = n23059 & n12619 ;
  assign n23060 = ~n12619 ;
  assign n12621 = n12148 & n23060 ;
  assign n12622 = n12620 | n12621 ;
  assign n23061 = ~n12622 ;
  assign n12623 = n12617 & n23061 ;
  assign n12624 = n12616 | n12623 ;
  assign n12625 = x74 & n12624 ;
  assign n12626 = x74 | n12624 ;
  assign n12627 = n12151 & n22880 ;
  assign n12628 = n140 & n12627 ;
  assign n23062 = ~n12157 ;
  assign n12629 = n23062 & n12628 ;
  assign n23063 = ~n12628 ;
  assign n12630 = n12157 & n23063 ;
  assign n12631 = n12629 | n12630 ;
  assign n23064 = ~n12631 ;
  assign n12632 = n12626 & n23064 ;
  assign n12633 = n12625 | n12632 ;
  assign n12634 = x75 & n12633 ;
  assign n12635 = x75 | n12633 ;
  assign n12636 = n12160 & n22884 ;
  assign n12637 = n140 & n12636 ;
  assign n23065 = ~n12166 ;
  assign n12638 = n23065 & n12637 ;
  assign n23066 = ~n12637 ;
  assign n12639 = n12166 & n23066 ;
  assign n12640 = n12638 | n12639 ;
  assign n23067 = ~n12640 ;
  assign n12641 = n12635 & n23067 ;
  assign n12642 = n12634 | n12641 ;
  assign n12643 = x76 & n12642 ;
  assign n12644 = x76 | n12642 ;
  assign n12645 = n12169 & n22888 ;
  assign n12646 = n140 & n12645 ;
  assign n23068 = ~n12175 ;
  assign n12647 = n23068 & n12646 ;
  assign n23069 = ~n12646 ;
  assign n12648 = n12175 & n23069 ;
  assign n12649 = n12647 | n12648 ;
  assign n23070 = ~n12649 ;
  assign n12650 = n12644 & n23070 ;
  assign n12651 = n12643 | n12650 ;
  assign n12652 = x77 & n12651 ;
  assign n12653 = x77 | n12651 ;
  assign n12654 = n12178 & n22892 ;
  assign n12655 = n140 & n12654 ;
  assign n23071 = ~n12184 ;
  assign n12656 = n23071 & n12655 ;
  assign n23072 = ~n12655 ;
  assign n12657 = n12184 & n23072 ;
  assign n12658 = n12656 | n12657 ;
  assign n23073 = ~n12658 ;
  assign n12659 = n12653 & n23073 ;
  assign n12660 = n12652 | n12659 ;
  assign n12661 = x78 & n12660 ;
  assign n12662 = x78 | n12660 ;
  assign n12663 = n12187 & n22895 ;
  assign n12664 = n140 & n12663 ;
  assign n23074 = ~n12193 ;
  assign n12665 = n23074 & n12664 ;
  assign n23075 = ~n12664 ;
  assign n12666 = n12193 & n23075 ;
  assign n12667 = n12665 | n12666 ;
  assign n23076 = ~n12667 ;
  assign n12668 = n12662 & n23076 ;
  assign n12669 = n12661 | n12668 ;
  assign n12670 = x79 & n12669 ;
  assign n12671 = x79 | n12669 ;
  assign n12672 = n12196 & n22899 ;
  assign n12673 = n140 & n12672 ;
  assign n23077 = ~n12202 ;
  assign n12674 = n23077 & n12673 ;
  assign n23078 = ~n12673 ;
  assign n12675 = n12202 & n23078 ;
  assign n12676 = n12674 | n12675 ;
  assign n23079 = ~n12676 ;
  assign n12677 = n12671 & n23079 ;
  assign n12678 = n12670 | n12677 ;
  assign n12679 = x80 & n12678 ;
  assign n12680 = x80 | n12678 ;
  assign n12681 = n12205 & n22903 ;
  assign n12682 = n140 & n12681 ;
  assign n23080 = ~n12211 ;
  assign n12683 = n23080 & n12682 ;
  assign n23081 = ~n12682 ;
  assign n12684 = n12211 & n23081 ;
  assign n12685 = n12683 | n12684 ;
  assign n23082 = ~n12685 ;
  assign n12686 = n12680 & n23082 ;
  assign n12687 = n12679 | n12686 ;
  assign n12688 = x81 & n12687 ;
  assign n12689 = x81 | n12687 ;
  assign n12690 = n12214 & n22906 ;
  assign n12691 = n140 & n12690 ;
  assign n23083 = ~n12220 ;
  assign n12692 = n23083 & n12691 ;
  assign n23084 = ~n12691 ;
  assign n12693 = n12220 & n23084 ;
  assign n12694 = n12692 | n12693 ;
  assign n23085 = ~n12694 ;
  assign n12695 = n12689 & n23085 ;
  assign n12696 = n12688 | n12695 ;
  assign n12697 = x82 & n12696 ;
  assign n12698 = x82 | n12696 ;
  assign n12699 = n12223 & n22910 ;
  assign n12700 = n140 & n12699 ;
  assign n23086 = ~n12229 ;
  assign n12701 = n23086 & n12700 ;
  assign n23087 = ~n12700 ;
  assign n12702 = n12229 & n23087 ;
  assign n12703 = n12701 | n12702 ;
  assign n23088 = ~n12703 ;
  assign n12704 = n12698 & n23088 ;
  assign n12705 = n12697 | n12704 ;
  assign n12706 = x83 & n12705 ;
  assign n12707 = x83 | n12705 ;
  assign n12708 = n12232 & n22913 ;
  assign n12709 = n140 & n12708 ;
  assign n12710 = n12238 & n12709 ;
  assign n12711 = n12238 | n12709 ;
  assign n23089 = ~n12710 ;
  assign n12712 = n23089 & n12711 ;
  assign n23090 = ~n12712 ;
  assign n12713 = n12707 & n23090 ;
  assign n12714 = n12706 | n12713 ;
  assign n12715 = x84 & n12714 ;
  assign n12716 = x84 | n12714 ;
  assign n12717 = n12241 & n22916 ;
  assign n12718 = n140 & n12717 ;
  assign n23091 = ~n12247 ;
  assign n12719 = n23091 & n12718 ;
  assign n23092 = ~n12718 ;
  assign n12720 = n12247 & n23092 ;
  assign n12721 = n12719 | n12720 ;
  assign n23093 = ~n12721 ;
  assign n12722 = n12716 & n23093 ;
  assign n12723 = n12715 | n12722 ;
  assign n12724 = x85 & n12723 ;
  assign n12725 = x85 | n12723 ;
  assign n12726 = n12250 & n22920 ;
  assign n12727 = n140 & n12726 ;
  assign n12728 = n12256 & n12727 ;
  assign n12729 = n12256 | n12727 ;
  assign n23094 = ~n12728 ;
  assign n12730 = n23094 & n12729 ;
  assign n23095 = ~n12730 ;
  assign n12731 = n12725 & n23095 ;
  assign n12732 = n12724 | n12731 ;
  assign n12733 = x86 & n12732 ;
  assign n12734 = x86 | n12732 ;
  assign n12735 = n12259 & n22924 ;
  assign n12736 = n140 & n12735 ;
  assign n23096 = ~n12265 ;
  assign n12737 = n23096 & n12736 ;
  assign n23097 = ~n12736 ;
  assign n12738 = n12265 & n23097 ;
  assign n12739 = n12737 | n12738 ;
  assign n23098 = ~n12739 ;
  assign n12740 = n12734 & n23098 ;
  assign n12741 = n12733 | n12740 ;
  assign n12742 = x87 & n12741 ;
  assign n12743 = x87 | n12741 ;
  assign n12744 = n12268 & n22927 ;
  assign n12745 = n140 & n12744 ;
  assign n12746 = n12274 & n12745 ;
  assign n12747 = n12274 | n12745 ;
  assign n23099 = ~n12746 ;
  assign n12748 = n23099 & n12747 ;
  assign n23100 = ~n12748 ;
  assign n12749 = n12743 & n23100 ;
  assign n12750 = n12742 | n12749 ;
  assign n12751 = x88 & n12750 ;
  assign n12752 = x88 | n12750 ;
  assign n12753 = n12277 & n22930 ;
  assign n12754 = n140 & n12753 ;
  assign n12755 = n12283 & n12754 ;
  assign n12756 = n12283 | n12754 ;
  assign n23101 = ~n12755 ;
  assign n12757 = n23101 & n12756 ;
  assign n23102 = ~n12757 ;
  assign n12758 = n12752 & n23102 ;
  assign n12759 = n12751 | n12758 ;
  assign n12760 = x89 & n12759 ;
  assign n12761 = x89 | n12759 ;
  assign n12762 = n12286 & n22933 ;
  assign n12763 = n140 & n12762 ;
  assign n12764 = n12292 & n12763 ;
  assign n12765 = n12292 | n12763 ;
  assign n23103 = ~n12764 ;
  assign n12766 = n23103 & n12765 ;
  assign n23104 = ~n12766 ;
  assign n12767 = n12761 & n23104 ;
  assign n12768 = n12760 | n12767 ;
  assign n12769 = x90 & n12768 ;
  assign n12770 = x90 | n12768 ;
  assign n12771 = n12295 & n22937 ;
  assign n12772 = n140 & n12771 ;
  assign n23105 = ~n12301 ;
  assign n12773 = n23105 & n12772 ;
  assign n23106 = ~n12772 ;
  assign n12774 = n12301 & n23106 ;
  assign n12775 = n12773 | n12774 ;
  assign n23107 = ~n12775 ;
  assign n12776 = n12770 & n23107 ;
  assign n12777 = n12769 | n12776 ;
  assign n12778 = x91 & n12777 ;
  assign n12779 = x91 | n12777 ;
  assign n12780 = n12304 & n22941 ;
  assign n12781 = n140 & n12780 ;
  assign n23108 = ~n12310 ;
  assign n12782 = n23108 & n12781 ;
  assign n23109 = ~n12781 ;
  assign n12783 = n12310 & n23109 ;
  assign n12784 = n12782 | n12783 ;
  assign n23110 = ~n12784 ;
  assign n12785 = n12779 & n23110 ;
  assign n12786 = n12778 | n12785 ;
  assign n12787 = x92 & n12786 ;
  assign n12788 = x92 | n12786 ;
  assign n12789 = n12313 & n22945 ;
  assign n12790 = n140 & n12789 ;
  assign n23111 = ~n12319 ;
  assign n12791 = n23111 & n12790 ;
  assign n23112 = ~n12790 ;
  assign n12792 = n12319 & n23112 ;
  assign n12793 = n12791 | n12792 ;
  assign n23113 = ~n12793 ;
  assign n12794 = n12788 & n23113 ;
  assign n12795 = n12787 | n12794 ;
  assign n12796 = x93 & n12795 ;
  assign n12797 = x93 | n12795 ;
  assign n12798 = n12322 & n22949 ;
  assign n12799 = n140 & n12798 ;
  assign n23114 = ~n12328 ;
  assign n12800 = n23114 & n12799 ;
  assign n23115 = ~n12799 ;
  assign n12801 = n12328 & n23115 ;
  assign n12802 = n12800 | n12801 ;
  assign n23116 = ~n12802 ;
  assign n12803 = n12797 & n23116 ;
  assign n12804 = n12796 | n12803 ;
  assign n12805 = x94 & n12804 ;
  assign n12806 = x94 | n12804 ;
  assign n12807 = n12331 & n22953 ;
  assign n12808 = n140 & n12807 ;
  assign n12809 = n12337 & n12808 ;
  assign n12810 = n12337 | n12808 ;
  assign n23117 = ~n12809 ;
  assign n12811 = n23117 & n12810 ;
  assign n23118 = ~n12811 ;
  assign n12812 = n12806 & n23118 ;
  assign n12813 = n12805 | n12812 ;
  assign n12814 = x95 & n12813 ;
  assign n12815 = x95 | n12813 ;
  assign n12816 = n12340 & n22957 ;
  assign n12817 = n140 & n12816 ;
  assign n23119 = ~n12346 ;
  assign n12818 = n23119 & n12817 ;
  assign n23120 = ~n12817 ;
  assign n12819 = n12346 & n23120 ;
  assign n12820 = n12818 | n12819 ;
  assign n23121 = ~n12820 ;
  assign n12821 = n12815 & n23121 ;
  assign n12822 = n12814 | n12821 ;
  assign n12823 = x96 & n12822 ;
  assign n12824 = x96 | n12822 ;
  assign n12825 = n12349 & n22961 ;
  assign n12826 = n140 & n12825 ;
  assign n23122 = ~n12355 ;
  assign n12827 = n23122 & n12826 ;
  assign n23123 = ~n12826 ;
  assign n12828 = n12355 & n23123 ;
  assign n12829 = n12827 | n12828 ;
  assign n23124 = ~n12829 ;
  assign n12830 = n12824 & n23124 ;
  assign n12831 = n12823 | n12830 ;
  assign n12832 = x97 & n12831 ;
  assign n12833 = x97 | n12831 ;
  assign n12834 = n12358 & n22964 ;
  assign n12835 = n140 & n12834 ;
  assign n23125 = ~n12364 ;
  assign n12836 = n23125 & n12835 ;
  assign n23126 = ~n12835 ;
  assign n12837 = n12364 & n23126 ;
  assign n12838 = n12836 | n12837 ;
  assign n23127 = ~n12838 ;
  assign n12839 = n12833 & n23127 ;
  assign n12840 = n12832 | n12839 ;
  assign n12841 = x98 & n12840 ;
  assign n12842 = x98 | n12840 ;
  assign n12843 = n12367 & n22967 ;
  assign n12844 = n140 & n12843 ;
  assign n23128 = ~n12373 ;
  assign n12845 = n23128 & n12844 ;
  assign n23129 = ~n12844 ;
  assign n12846 = n12373 & n23129 ;
  assign n12847 = n12845 | n12846 ;
  assign n23130 = ~n12847 ;
  assign n12848 = n12842 & n23130 ;
  assign n12849 = n12841 | n12848 ;
  assign n12850 = x99 & n12849 ;
  assign n12851 = x99 | n12849 ;
  assign n12852 = n12376 & n22971 ;
  assign n12853 = n140 & n12852 ;
  assign n23131 = ~n12382 ;
  assign n12854 = n23131 & n12853 ;
  assign n23132 = ~n12853 ;
  assign n12855 = n12382 & n23132 ;
  assign n12856 = n12854 | n12855 ;
  assign n23133 = ~n12856 ;
  assign n12857 = n12851 & n23133 ;
  assign n12858 = n12850 | n12857 ;
  assign n12859 = x100 & n12858 ;
  assign n12860 = x100 | n12858 ;
  assign n12861 = n12385 & n22975 ;
  assign n12862 = n140 & n12861 ;
  assign n23134 = ~n12391 ;
  assign n12863 = n23134 & n12862 ;
  assign n23135 = ~n12862 ;
  assign n12864 = n12391 & n23135 ;
  assign n12865 = n12863 | n12864 ;
  assign n23136 = ~n12865 ;
  assign n12866 = n12860 & n23136 ;
  assign n12867 = n12859 | n12866 ;
  assign n12868 = x101 & n12867 ;
  assign n12869 = x101 | n12867 ;
  assign n12870 = n12394 & n22979 ;
  assign n12871 = n140 & n12870 ;
  assign n23137 = ~n12400 ;
  assign n12872 = n23137 & n12871 ;
  assign n23138 = ~n12871 ;
  assign n12873 = n12400 & n23138 ;
  assign n12874 = n12872 | n12873 ;
  assign n23139 = ~n12874 ;
  assign n12875 = n12869 & n23139 ;
  assign n12876 = n12868 | n12875 ;
  assign n12877 = x102 & n12876 ;
  assign n12878 = x102 | n12876 ;
  assign n12879 = n12403 & n22982 ;
  assign n12880 = n140 & n12879 ;
  assign n12881 = n12409 & n12880 ;
  assign n12882 = n12409 | n12880 ;
  assign n23140 = ~n12881 ;
  assign n12883 = n23140 & n12882 ;
  assign n23141 = ~n12883 ;
  assign n12884 = n12878 & n23141 ;
  assign n12885 = n12877 | n12884 ;
  assign n12886 = x103 & n12885 ;
  assign n12887 = x103 | n12885 ;
  assign n12888 = n12412 & n22986 ;
  assign n12889 = n140 & n12888 ;
  assign n23142 = ~n12418 ;
  assign n12890 = n23142 & n12889 ;
  assign n23143 = ~n12889 ;
  assign n12891 = n12418 & n23143 ;
  assign n12892 = n12890 | n12891 ;
  assign n23144 = ~n12892 ;
  assign n12893 = n12887 & n23144 ;
  assign n12894 = n12886 | n12893 ;
  assign n12895 = x104 & n12894 ;
  assign n12896 = x104 | n12894 ;
  assign n12897 = n12421 & n22990 ;
  assign n12898 = n140 & n12897 ;
  assign n23145 = ~n12427 ;
  assign n12899 = n23145 & n12898 ;
  assign n23146 = ~n12898 ;
  assign n12900 = n12427 & n23146 ;
  assign n12901 = n12899 | n12900 ;
  assign n23147 = ~n12901 ;
  assign n12902 = n12896 & n23147 ;
  assign n12903 = n12895 | n12902 ;
  assign n12904 = x105 & n12903 ;
  assign n12905 = x105 | n12903 ;
  assign n12906 = n12430 & n22993 ;
  assign n12907 = n140 & n12906 ;
  assign n12908 = n12436 & n12907 ;
  assign n12909 = n12436 | n12907 ;
  assign n23148 = ~n12908 ;
  assign n12910 = n23148 & n12909 ;
  assign n23149 = ~n12910 ;
  assign n12911 = n12905 & n23149 ;
  assign n12912 = n12904 | n12911 ;
  assign n12913 = x106 & n12912 ;
  assign n12914 = x106 | n12912 ;
  assign n12915 = n12439 & n22997 ;
  assign n12916 = n140 & n12915 ;
  assign n23150 = ~n12445 ;
  assign n12917 = n23150 & n12916 ;
  assign n23151 = ~n12916 ;
  assign n12918 = n12445 & n23151 ;
  assign n12919 = n12917 | n12918 ;
  assign n23152 = ~n12919 ;
  assign n12920 = n12914 & n23152 ;
  assign n12921 = n12913 | n12920 ;
  assign n12922 = x107 & n12921 ;
  assign n12923 = x107 | n12921 ;
  assign n12924 = n12448 & n23001 ;
  assign n12925 = n140 & n12924 ;
  assign n23153 = ~n12454 ;
  assign n12926 = n23153 & n12925 ;
  assign n23154 = ~n12925 ;
  assign n12927 = n12454 & n23154 ;
  assign n12928 = n12926 | n12927 ;
  assign n23155 = ~n12928 ;
  assign n12929 = n12923 & n23155 ;
  assign n12930 = n12922 | n12929 ;
  assign n12931 = x108 & n12930 ;
  assign n12932 = x108 | n12930 ;
  assign n12933 = n12457 & n23005 ;
  assign n12934 = n140 & n12933 ;
  assign n23156 = ~n12463 ;
  assign n12935 = n23156 & n12934 ;
  assign n23157 = ~n12934 ;
  assign n12936 = n12463 & n23157 ;
  assign n12937 = n12935 | n12936 ;
  assign n23158 = ~n12937 ;
  assign n12938 = n12932 & n23158 ;
  assign n12939 = n12931 | n12938 ;
  assign n12940 = x109 & n12939 ;
  assign n12941 = x109 | n12939 ;
  assign n12942 = n12466 & n23009 ;
  assign n12943 = n140 & n12942 ;
  assign n23159 = ~n12472 ;
  assign n12944 = n23159 & n12943 ;
  assign n23160 = ~n12943 ;
  assign n12945 = n12472 & n23160 ;
  assign n12946 = n12944 | n12945 ;
  assign n23161 = ~n12946 ;
  assign n12947 = n12941 & n23161 ;
  assign n12948 = n12940 | n12947 ;
  assign n12949 = x110 & n12948 ;
  assign n12950 = x110 | n12948 ;
  assign n12951 = n12475 & n23013 ;
  assign n12952 = n140 & n12951 ;
  assign n23162 = ~n12481 ;
  assign n12953 = n23162 & n12952 ;
  assign n23163 = ~n12952 ;
  assign n12954 = n12481 & n23163 ;
  assign n12955 = n12953 | n12954 ;
  assign n23164 = ~n12955 ;
  assign n12956 = n12950 & n23164 ;
  assign n12957 = n12949 | n12956 ;
  assign n12958 = x111 & n12957 ;
  assign n12959 = x111 | n12957 ;
  assign n12960 = n12484 & n23016 ;
  assign n12961 = n140 & n12960 ;
  assign n12962 = n12490 & n12961 ;
  assign n12963 = n12490 | n12961 ;
  assign n23165 = ~n12962 ;
  assign n12964 = n23165 & n12963 ;
  assign n23166 = ~n12964 ;
  assign n12965 = n12959 & n23166 ;
  assign n12966 = n12958 | n12965 ;
  assign n12967 = x112 & n12966 ;
  assign n12968 = x112 | n12966 ;
  assign n12969 = n12493 & n23019 ;
  assign n12970 = n140 & n12969 ;
  assign n12971 = n12499 & n12970 ;
  assign n12972 = n12499 | n12970 ;
  assign n23167 = ~n12971 ;
  assign n12973 = n23167 & n12972 ;
  assign n23168 = ~n12973 ;
  assign n12974 = n12968 & n23168 ;
  assign n12975 = n12967 | n12974 ;
  assign n12976 = x113 & n12975 ;
  assign n12977 = x113 | n12975 ;
  assign n12978 = n12502 & n23022 ;
  assign n12979 = n140 & n12978 ;
  assign n12980 = n12508 & n12979 ;
  assign n12981 = n12508 | n12979 ;
  assign n23169 = ~n12980 ;
  assign n12982 = n23169 & n12981 ;
  assign n23170 = ~n12982 ;
  assign n12983 = n12977 & n23170 ;
  assign n12984 = n12976 | n12983 ;
  assign n12985 = x114 & n12984 ;
  assign n12986 = x114 | n12984 ;
  assign n12987 = n12511 & n23026 ;
  assign n12988 = n140 & n12987 ;
  assign n23171 = ~n12517 ;
  assign n12989 = n23171 & n12988 ;
  assign n23172 = ~n12988 ;
  assign n12990 = n12517 & n23172 ;
  assign n12991 = n12989 | n12990 ;
  assign n23173 = ~n12991 ;
  assign n12992 = n12986 & n23173 ;
  assign n12993 = n12985 | n12992 ;
  assign n12994 = x115 & n12993 ;
  assign n12995 = x115 | n12993 ;
  assign n12996 = n12520 & n23029 ;
  assign n12997 = n140 & n12996 ;
  assign n12998 = n12526 & n12997 ;
  assign n12999 = n12526 | n12997 ;
  assign n23174 = ~n12998 ;
  assign n13000 = n23174 & n12999 ;
  assign n23175 = ~n13000 ;
  assign n13001 = n12995 & n23175 ;
  assign n13002 = n12994 | n13001 ;
  assign n13003 = x116 & n13002 ;
  assign n13004 = x116 | n13002 ;
  assign n23176 = ~n12543 ;
  assign n13005 = n23176 & n13004 ;
  assign n13006 = n13003 | n13005 ;
  assign n13008 = x117 & n13006 ;
  assign n13009 = n18308 | n13008 ;
  assign n13007 = x117 | n13006 ;
  assign n13010 = n18318 & n12062 ;
  assign n13011 = n12537 & n13010 ;
  assign n13012 = n21884 | n13011 ;
  assign n23177 = ~n13012 ;
  assign n13013 = n13007 & n23177 ;
  assign n13014 = n13009 | n13013 ;
  assign n23178 = ~n13003 ;
  assign n13015 = n23178 & n13004 ;
  assign n139 = ~n13014 ;
  assign n13016 = n139 & n13015 ;
  assign n13017 = n12543 & n13016 ;
  assign n13018 = n12543 | n13016 ;
  assign n23180 = ~n13017 ;
  assign n13019 = n23180 & n13018 ;
  assign n23181 = ~x9 ;
  assign n13020 = n23181 & x64 ;
  assign n13022 = x65 | n13020 ;
  assign n13021 = x65 & n13020 ;
  assign n13023 = x64 & n139 ;
  assign n13024 = x10 & n13023 ;
  assign n13025 = x10 | n13023 ;
  assign n23182 = ~n13024 ;
  assign n13026 = n23182 & n13025 ;
  assign n23183 = ~n13021 ;
  assign n13027 = n23183 & n13026 ;
  assign n23184 = ~n13027 ;
  assign n13028 = n13022 & n23184 ;
  assign n13029 = x66 | n13028 ;
  assign n13030 = x66 & n13028 ;
  assign n13031 = n12545 & n139 ;
  assign n13032 = n23039 & n13031 ;
  assign n13033 = n12549 | n13032 ;
  assign n13034 = n12551 & n13031 ;
  assign n23185 = ~n13034 ;
  assign n13035 = n13033 & n23185 ;
  assign n23186 = ~n13030 ;
  assign n13036 = n23186 & n13035 ;
  assign n23187 = ~n13036 ;
  assign n13037 = n13029 & n23187 ;
  assign n13038 = x67 | n13037 ;
  assign n13039 = x67 & n13037 ;
  assign n23188 = ~n12554 ;
  assign n13040 = n12553 & n23188 ;
  assign n13041 = n139 & n13040 ;
  assign n13042 = n23042 & n13041 ;
  assign n23189 = ~n13041 ;
  assign n13043 = n12559 & n23189 ;
  assign n13044 = n13042 | n13043 ;
  assign n23190 = ~n13039 ;
  assign n13045 = n23190 & n13044 ;
  assign n23191 = ~n13045 ;
  assign n13046 = n13038 & n23191 ;
  assign n13047 = x68 | n13046 ;
  assign n13048 = x68 & n13046 ;
  assign n13049 = n12562 | n13014 ;
  assign n23192 = ~n13049 ;
  assign n13050 = n12569 & n23192 ;
  assign n13051 = n12563 & n23192 ;
  assign n23193 = ~n13051 ;
  assign n13052 = n12568 & n23193 ;
  assign n13053 = n13050 | n13052 ;
  assign n23194 = ~n13048 ;
  assign n13054 = n23194 & n13053 ;
  assign n23195 = ~n13054 ;
  assign n13055 = n13047 & n23195 ;
  assign n13056 = x69 | n13055 ;
  assign n13057 = x69 & n13055 ;
  assign n23196 = ~n12571 ;
  assign n13058 = n23196 & n12572 ;
  assign n13059 = n139 & n13058 ;
  assign n13060 = n12577 & n13059 ;
  assign n13061 = n12577 | n13059 ;
  assign n23197 = ~n13060 ;
  assign n13062 = n23197 & n13061 ;
  assign n23198 = ~n13057 ;
  assign n13063 = n23198 & n13062 ;
  assign n23199 = ~n13063 ;
  assign n13064 = n13056 & n23199 ;
  assign n13065 = x70 | n13064 ;
  assign n13066 = x70 & n13064 ;
  assign n23200 = ~n12580 ;
  assign n13067 = n23200 & n12581 ;
  assign n13068 = n139 & n13067 ;
  assign n13069 = n12586 & n13068 ;
  assign n13070 = n12586 | n13068 ;
  assign n23201 = ~n13069 ;
  assign n13071 = n23201 & n13070 ;
  assign n23202 = ~n13066 ;
  assign n13072 = n23202 & n13071 ;
  assign n23203 = ~n13072 ;
  assign n13073 = n13065 & n23203 ;
  assign n13074 = x71 | n13073 ;
  assign n13075 = x71 & n13073 ;
  assign n23204 = ~n12589 ;
  assign n13076 = n23204 & n12590 ;
  assign n13077 = n139 & n13076 ;
  assign n13078 = n12595 & n13077 ;
  assign n13079 = n12595 | n13077 ;
  assign n23205 = ~n13078 ;
  assign n13080 = n23205 & n13079 ;
  assign n23206 = ~n13075 ;
  assign n13081 = n23206 & n13080 ;
  assign n23207 = ~n13081 ;
  assign n13082 = n13074 & n23207 ;
  assign n13083 = x72 | n13082 ;
  assign n13084 = x72 & n13082 ;
  assign n23208 = ~n12598 ;
  assign n13085 = n23208 & n12599 ;
  assign n13086 = n139 & n13085 ;
  assign n13087 = n12604 & n13086 ;
  assign n13088 = n12604 | n13086 ;
  assign n23209 = ~n13087 ;
  assign n13089 = n23209 & n13088 ;
  assign n23210 = ~n13084 ;
  assign n13090 = n23210 & n13089 ;
  assign n23211 = ~n13090 ;
  assign n13091 = n13083 & n23211 ;
  assign n13092 = x73 | n13091 ;
  assign n13093 = x73 & n13091 ;
  assign n23212 = ~n12607 ;
  assign n13094 = n23212 & n12608 ;
  assign n13095 = n139 & n13094 ;
  assign n13096 = n23058 & n13095 ;
  assign n23213 = ~n13095 ;
  assign n13097 = n12613 & n23213 ;
  assign n13098 = n13096 | n13097 ;
  assign n23214 = ~n13093 ;
  assign n13099 = n23214 & n13098 ;
  assign n23215 = ~n13099 ;
  assign n13100 = n13092 & n23215 ;
  assign n13101 = x74 | n13100 ;
  assign n13102 = x74 & n13100 ;
  assign n23216 = ~n12616 ;
  assign n13103 = n23216 & n12617 ;
  assign n13104 = n139 & n13103 ;
  assign n13105 = n23061 & n13104 ;
  assign n23217 = ~n13104 ;
  assign n13106 = n12622 & n23217 ;
  assign n13107 = n13105 | n13106 ;
  assign n23218 = ~n13102 ;
  assign n13108 = n23218 & n13107 ;
  assign n23219 = ~n13108 ;
  assign n13109 = n13101 & n23219 ;
  assign n13110 = x75 | n13109 ;
  assign n13111 = x75 & n13109 ;
  assign n23220 = ~n12625 ;
  assign n13112 = n23220 & n12626 ;
  assign n13113 = n139 & n13112 ;
  assign n13114 = n23064 & n13113 ;
  assign n23221 = ~n13113 ;
  assign n13115 = n12631 & n23221 ;
  assign n13116 = n13114 | n13115 ;
  assign n23222 = ~n13111 ;
  assign n13117 = n23222 & n13116 ;
  assign n23223 = ~n13117 ;
  assign n13118 = n13110 & n23223 ;
  assign n13119 = x76 | n13118 ;
  assign n13120 = x76 & n13118 ;
  assign n23224 = ~n12634 ;
  assign n13121 = n23224 & n12635 ;
  assign n13122 = n139 & n13121 ;
  assign n13123 = n12640 & n13122 ;
  assign n13124 = n12640 | n13122 ;
  assign n23225 = ~n13123 ;
  assign n13125 = n23225 & n13124 ;
  assign n23226 = ~n13120 ;
  assign n13126 = n23226 & n13125 ;
  assign n23227 = ~n13126 ;
  assign n13127 = n13119 & n23227 ;
  assign n13128 = x77 | n13127 ;
  assign n13129 = x77 & n13127 ;
  assign n23228 = ~n12643 ;
  assign n13130 = n23228 & n12644 ;
  assign n13131 = n139 & n13130 ;
  assign n13132 = n23070 & n13131 ;
  assign n23229 = ~n13131 ;
  assign n13133 = n12649 & n23229 ;
  assign n13134 = n13132 | n13133 ;
  assign n23230 = ~n13129 ;
  assign n13135 = n23230 & n13134 ;
  assign n23231 = ~n13135 ;
  assign n13136 = n13128 & n23231 ;
  assign n13137 = x78 | n13136 ;
  assign n13138 = x78 & n13136 ;
  assign n23232 = ~n12652 ;
  assign n13139 = n23232 & n12653 ;
  assign n13140 = n139 & n13139 ;
  assign n13141 = n23073 & n13140 ;
  assign n23233 = ~n13140 ;
  assign n13142 = n12658 & n23233 ;
  assign n13143 = n13141 | n13142 ;
  assign n23234 = ~n13138 ;
  assign n13144 = n23234 & n13143 ;
  assign n23235 = ~n13144 ;
  assign n13145 = n13137 & n23235 ;
  assign n13146 = x79 | n13145 ;
  assign n13147 = x79 & n13145 ;
  assign n23236 = ~n12661 ;
  assign n13148 = n23236 & n12662 ;
  assign n13149 = n139 & n13148 ;
  assign n13150 = n23076 & n13149 ;
  assign n23237 = ~n13149 ;
  assign n13151 = n12667 & n23237 ;
  assign n13152 = n13150 | n13151 ;
  assign n23238 = ~n13147 ;
  assign n13153 = n23238 & n13152 ;
  assign n23239 = ~n13153 ;
  assign n13154 = n13146 & n23239 ;
  assign n13155 = x80 | n13154 ;
  assign n13156 = x80 & n13154 ;
  assign n23240 = ~n12670 ;
  assign n13157 = n23240 & n12671 ;
  assign n13158 = n139 & n13157 ;
  assign n13159 = n12676 & n13158 ;
  assign n13160 = n12676 | n13158 ;
  assign n23241 = ~n13159 ;
  assign n13161 = n23241 & n13160 ;
  assign n23242 = ~n13156 ;
  assign n13162 = n23242 & n13161 ;
  assign n23243 = ~n13162 ;
  assign n13163 = n13155 & n23243 ;
  assign n13164 = x81 | n13163 ;
  assign n13165 = x81 & n13163 ;
  assign n23244 = ~n12679 ;
  assign n13166 = n23244 & n12680 ;
  assign n13167 = n139 & n13166 ;
  assign n13168 = n23082 & n13167 ;
  assign n23245 = ~n13167 ;
  assign n13169 = n12685 & n23245 ;
  assign n13170 = n13168 | n13169 ;
  assign n23246 = ~n13165 ;
  assign n13171 = n23246 & n13170 ;
  assign n23247 = ~n13171 ;
  assign n13172 = n13164 & n23247 ;
  assign n13173 = x82 | n13172 ;
  assign n13174 = x82 & n13172 ;
  assign n23248 = ~n12688 ;
  assign n13175 = n23248 & n12689 ;
  assign n13176 = n139 & n13175 ;
  assign n13177 = n23085 & n13176 ;
  assign n23249 = ~n13176 ;
  assign n13178 = n12694 & n23249 ;
  assign n13179 = n13177 | n13178 ;
  assign n23250 = ~n13174 ;
  assign n13180 = n23250 & n13179 ;
  assign n23251 = ~n13180 ;
  assign n13181 = n13173 & n23251 ;
  assign n13182 = x83 | n13181 ;
  assign n13183 = x83 & n13181 ;
  assign n23252 = ~n12697 ;
  assign n13184 = n23252 & n12698 ;
  assign n13185 = n139 & n13184 ;
  assign n13186 = n23088 & n13185 ;
  assign n23253 = ~n13185 ;
  assign n13187 = n12703 & n23253 ;
  assign n13188 = n13186 | n13187 ;
  assign n23254 = ~n13183 ;
  assign n13189 = n23254 & n13188 ;
  assign n23255 = ~n13189 ;
  assign n13190 = n13182 & n23255 ;
  assign n13191 = x84 | n13190 ;
  assign n13192 = x84 & n13190 ;
  assign n23256 = ~n12706 ;
  assign n13193 = n23256 & n12707 ;
  assign n13194 = n139 & n13193 ;
  assign n13195 = n12712 & n13194 ;
  assign n13196 = n12712 | n13194 ;
  assign n23257 = ~n13195 ;
  assign n13197 = n23257 & n13196 ;
  assign n23258 = ~n13192 ;
  assign n13198 = n23258 & n13197 ;
  assign n23259 = ~n13198 ;
  assign n13199 = n13191 & n23259 ;
  assign n13200 = x85 | n13199 ;
  assign n13201 = x85 & n13199 ;
  assign n23260 = ~n12715 ;
  assign n13202 = n23260 & n12716 ;
  assign n13203 = n139 & n13202 ;
  assign n13204 = n23093 & n13203 ;
  assign n23261 = ~n13203 ;
  assign n13205 = n12721 & n23261 ;
  assign n13206 = n13204 | n13205 ;
  assign n23262 = ~n13201 ;
  assign n13207 = n23262 & n13206 ;
  assign n23263 = ~n13207 ;
  assign n13208 = n13200 & n23263 ;
  assign n13209 = x86 | n13208 ;
  assign n13210 = x86 & n13208 ;
  assign n23264 = ~n12724 ;
  assign n13211 = n23264 & n12725 ;
  assign n13212 = n139 & n13211 ;
  assign n13213 = n12730 & n13212 ;
  assign n13214 = n12730 | n13212 ;
  assign n23265 = ~n13213 ;
  assign n13215 = n23265 & n13214 ;
  assign n23266 = ~n13210 ;
  assign n13216 = n23266 & n13215 ;
  assign n23267 = ~n13216 ;
  assign n13217 = n13209 & n23267 ;
  assign n13218 = x87 | n13217 ;
  assign n13219 = x87 & n13217 ;
  assign n23268 = ~n12733 ;
  assign n13220 = n23268 & n12734 ;
  assign n13221 = n139 & n13220 ;
  assign n13222 = n12739 & n13221 ;
  assign n13223 = n12739 | n13221 ;
  assign n23269 = ~n13222 ;
  assign n13224 = n23269 & n13223 ;
  assign n23270 = ~n13219 ;
  assign n13225 = n23270 & n13224 ;
  assign n23271 = ~n13225 ;
  assign n13226 = n13218 & n23271 ;
  assign n13227 = x88 | n13226 ;
  assign n13228 = x88 & n13226 ;
  assign n23272 = ~n12742 ;
  assign n13229 = n23272 & n12743 ;
  assign n13230 = n139 & n13229 ;
  assign n13231 = n12748 & n13230 ;
  assign n13232 = n12748 | n13230 ;
  assign n23273 = ~n13231 ;
  assign n13233 = n23273 & n13232 ;
  assign n23274 = ~n13228 ;
  assign n13234 = n23274 & n13233 ;
  assign n23275 = ~n13234 ;
  assign n13235 = n13227 & n23275 ;
  assign n13236 = x89 | n13235 ;
  assign n13237 = x89 & n13235 ;
  assign n23276 = ~n12751 ;
  assign n13238 = n23276 & n12752 ;
  assign n13239 = n139 & n13238 ;
  assign n13240 = n12757 & n13239 ;
  assign n13241 = n12757 | n13239 ;
  assign n23277 = ~n13240 ;
  assign n13242 = n23277 & n13241 ;
  assign n23278 = ~n13237 ;
  assign n13243 = n23278 & n13242 ;
  assign n23279 = ~n13243 ;
  assign n13244 = n13236 & n23279 ;
  assign n13245 = x90 | n13244 ;
  assign n13246 = x90 & n13244 ;
  assign n23280 = ~n12760 ;
  assign n13247 = n23280 & n12761 ;
  assign n13248 = n139 & n13247 ;
  assign n13249 = n12766 & n13248 ;
  assign n13250 = n12766 | n13248 ;
  assign n23281 = ~n13249 ;
  assign n13251 = n23281 & n13250 ;
  assign n23282 = ~n13246 ;
  assign n13252 = n23282 & n13251 ;
  assign n23283 = ~n13252 ;
  assign n13253 = n13245 & n23283 ;
  assign n13254 = x91 | n13253 ;
  assign n13255 = x91 & n13253 ;
  assign n23284 = ~n12769 ;
  assign n13256 = n23284 & n12770 ;
  assign n13257 = n139 & n13256 ;
  assign n13258 = n23107 & n13257 ;
  assign n23285 = ~n13257 ;
  assign n13259 = n12775 & n23285 ;
  assign n13260 = n13258 | n13259 ;
  assign n23286 = ~n13255 ;
  assign n13261 = n23286 & n13260 ;
  assign n23287 = ~n13261 ;
  assign n13262 = n13254 & n23287 ;
  assign n13263 = x92 | n13262 ;
  assign n13264 = x92 & n13262 ;
  assign n23288 = ~n12778 ;
  assign n13265 = n23288 & n12779 ;
  assign n13266 = n139 & n13265 ;
  assign n13267 = n23110 & n13266 ;
  assign n23289 = ~n13266 ;
  assign n13268 = n12784 & n23289 ;
  assign n13269 = n13267 | n13268 ;
  assign n23290 = ~n13264 ;
  assign n13270 = n23290 & n13269 ;
  assign n23291 = ~n13270 ;
  assign n13271 = n13263 & n23291 ;
  assign n13272 = x93 | n13271 ;
  assign n13273 = x93 & n13271 ;
  assign n23292 = ~n12787 ;
  assign n13274 = n23292 & n12788 ;
  assign n13275 = n139 & n13274 ;
  assign n13276 = n12793 & n13275 ;
  assign n13277 = n12793 | n13275 ;
  assign n23293 = ~n13276 ;
  assign n13278 = n23293 & n13277 ;
  assign n23294 = ~n13273 ;
  assign n13279 = n23294 & n13278 ;
  assign n23295 = ~n13279 ;
  assign n13280 = n13272 & n23295 ;
  assign n13281 = x94 | n13280 ;
  assign n13282 = x94 & n13280 ;
  assign n23296 = ~n12796 ;
  assign n13283 = n23296 & n12797 ;
  assign n13284 = n139 & n13283 ;
  assign n13285 = n23116 & n13284 ;
  assign n23297 = ~n13284 ;
  assign n13286 = n12802 & n23297 ;
  assign n13287 = n13285 | n13286 ;
  assign n23298 = ~n13282 ;
  assign n13288 = n23298 & n13287 ;
  assign n23299 = ~n13288 ;
  assign n13289 = n13281 & n23299 ;
  assign n13290 = x95 | n13289 ;
  assign n13291 = x95 & n13289 ;
  assign n23300 = ~n12805 ;
  assign n13292 = n23300 & n12806 ;
  assign n13293 = n139 & n13292 ;
  assign n13294 = n12811 & n13293 ;
  assign n13295 = n12811 | n13293 ;
  assign n23301 = ~n13294 ;
  assign n13296 = n23301 & n13295 ;
  assign n23302 = ~n13291 ;
  assign n13297 = n23302 & n13296 ;
  assign n23303 = ~n13297 ;
  assign n13298 = n13290 & n23303 ;
  assign n13299 = x96 | n13298 ;
  assign n13300 = x96 & n13298 ;
  assign n23304 = ~n12814 ;
  assign n13301 = n23304 & n12815 ;
  assign n13302 = n139 & n13301 ;
  assign n13303 = n12820 & n13302 ;
  assign n13304 = n12820 | n13302 ;
  assign n23305 = ~n13303 ;
  assign n13305 = n23305 & n13304 ;
  assign n23306 = ~n13300 ;
  assign n13306 = n23306 & n13305 ;
  assign n23307 = ~n13306 ;
  assign n13307 = n13299 & n23307 ;
  assign n13308 = x97 | n13307 ;
  assign n13309 = x97 & n13307 ;
  assign n23308 = ~n12823 ;
  assign n13310 = n23308 & n12824 ;
  assign n13311 = n139 & n13310 ;
  assign n13312 = n23124 & n13311 ;
  assign n23309 = ~n13311 ;
  assign n13313 = n12829 & n23309 ;
  assign n13314 = n13312 | n13313 ;
  assign n23310 = ~n13309 ;
  assign n13315 = n23310 & n13314 ;
  assign n23311 = ~n13315 ;
  assign n13316 = n13308 & n23311 ;
  assign n13317 = x98 | n13316 ;
  assign n13318 = x98 & n13316 ;
  assign n23312 = ~n12832 ;
  assign n13319 = n23312 & n12833 ;
  assign n13320 = n139 & n13319 ;
  assign n13321 = n23127 & n13320 ;
  assign n23313 = ~n13320 ;
  assign n13322 = n12838 & n23313 ;
  assign n13323 = n13321 | n13322 ;
  assign n23314 = ~n13318 ;
  assign n13324 = n23314 & n13323 ;
  assign n23315 = ~n13324 ;
  assign n13325 = n13317 & n23315 ;
  assign n13326 = x99 | n13325 ;
  assign n13327 = x99 & n13325 ;
  assign n23316 = ~n12841 ;
  assign n13328 = n23316 & n12842 ;
  assign n13329 = n139 & n13328 ;
  assign n13330 = n23130 & n13329 ;
  assign n23317 = ~n13329 ;
  assign n13331 = n12847 & n23317 ;
  assign n13332 = n13330 | n13331 ;
  assign n23318 = ~n13327 ;
  assign n13333 = n23318 & n13332 ;
  assign n23319 = ~n13333 ;
  assign n13334 = n13326 & n23319 ;
  assign n13335 = x100 | n13334 ;
  assign n13336 = x100 & n13334 ;
  assign n23320 = ~n12850 ;
  assign n13337 = n23320 & n12851 ;
  assign n13338 = n139 & n13337 ;
  assign n13339 = n23133 & n13338 ;
  assign n23321 = ~n13338 ;
  assign n13340 = n12856 & n23321 ;
  assign n13341 = n13339 | n13340 ;
  assign n23322 = ~n13336 ;
  assign n13342 = n23322 & n13341 ;
  assign n23323 = ~n13342 ;
  assign n13343 = n13335 & n23323 ;
  assign n13344 = x101 | n13343 ;
  assign n13345 = x101 & n13343 ;
  assign n23324 = ~n12859 ;
  assign n13346 = n23324 & n12860 ;
  assign n13347 = n139 & n13346 ;
  assign n13348 = n23136 & n13347 ;
  assign n23325 = ~n13347 ;
  assign n13349 = n12865 & n23325 ;
  assign n13350 = n13348 | n13349 ;
  assign n23326 = ~n13345 ;
  assign n13351 = n23326 & n13350 ;
  assign n23327 = ~n13351 ;
  assign n13352 = n13344 & n23327 ;
  assign n13353 = x102 | n13352 ;
  assign n13354 = x102 & n13352 ;
  assign n23328 = ~n12868 ;
  assign n13355 = n23328 & n12869 ;
  assign n13356 = n139 & n13355 ;
  assign n13357 = n12874 & n13356 ;
  assign n13358 = n12874 | n13356 ;
  assign n23329 = ~n13357 ;
  assign n13359 = n23329 & n13358 ;
  assign n23330 = ~n13354 ;
  assign n13360 = n23330 & n13359 ;
  assign n23331 = ~n13360 ;
  assign n13361 = n13353 & n23331 ;
  assign n13362 = x103 | n13361 ;
  assign n13363 = x103 & n13361 ;
  assign n23332 = ~n12877 ;
  assign n13364 = n23332 & n12878 ;
  assign n13365 = n139 & n13364 ;
  assign n13366 = n12883 & n13365 ;
  assign n13367 = n12883 | n13365 ;
  assign n23333 = ~n13366 ;
  assign n13368 = n23333 & n13367 ;
  assign n23334 = ~n13363 ;
  assign n13369 = n23334 & n13368 ;
  assign n23335 = ~n13369 ;
  assign n13370 = n13362 & n23335 ;
  assign n13371 = x104 | n13370 ;
  assign n13372 = x104 & n13370 ;
  assign n23336 = ~n12886 ;
  assign n13373 = n23336 & n12887 ;
  assign n13374 = n139 & n13373 ;
  assign n13375 = n23144 & n13374 ;
  assign n23337 = ~n13374 ;
  assign n13376 = n12892 & n23337 ;
  assign n13377 = n13375 | n13376 ;
  assign n23338 = ~n13372 ;
  assign n13378 = n23338 & n13377 ;
  assign n23339 = ~n13378 ;
  assign n13379 = n13371 & n23339 ;
  assign n13380 = x105 | n13379 ;
  assign n13381 = x105 & n13379 ;
  assign n23340 = ~n12895 ;
  assign n13382 = n23340 & n12896 ;
  assign n13383 = n139 & n13382 ;
  assign n13384 = n23147 & n13383 ;
  assign n23341 = ~n13383 ;
  assign n13385 = n12901 & n23341 ;
  assign n13386 = n13384 | n13385 ;
  assign n23342 = ~n13381 ;
  assign n13387 = n23342 & n13386 ;
  assign n23343 = ~n13387 ;
  assign n13388 = n13380 & n23343 ;
  assign n13389 = x106 | n13388 ;
  assign n13390 = x106 & n13388 ;
  assign n23344 = ~n12904 ;
  assign n13391 = n23344 & n12905 ;
  assign n13392 = n139 & n13391 ;
  assign n13393 = n12910 & n13392 ;
  assign n13394 = n12910 | n13392 ;
  assign n23345 = ~n13393 ;
  assign n13395 = n23345 & n13394 ;
  assign n23346 = ~n13390 ;
  assign n13396 = n23346 & n13395 ;
  assign n23347 = ~n13396 ;
  assign n13397 = n13389 & n23347 ;
  assign n13398 = x107 | n13397 ;
  assign n13399 = x107 & n13397 ;
  assign n23348 = ~n12913 ;
  assign n13400 = n23348 & n12914 ;
  assign n13401 = n139 & n13400 ;
  assign n13402 = n12919 & n13401 ;
  assign n13403 = n12919 | n13401 ;
  assign n23349 = ~n13402 ;
  assign n13404 = n23349 & n13403 ;
  assign n23350 = ~n13399 ;
  assign n13405 = n23350 & n13404 ;
  assign n23351 = ~n13405 ;
  assign n13406 = n13398 & n23351 ;
  assign n13407 = x108 | n13406 ;
  assign n13408 = x108 & n13406 ;
  assign n23352 = ~n12922 ;
  assign n13409 = n23352 & n12923 ;
  assign n13410 = n139 & n13409 ;
  assign n13411 = n12928 & n13410 ;
  assign n13412 = n12928 | n13410 ;
  assign n23353 = ~n13411 ;
  assign n13413 = n23353 & n13412 ;
  assign n23354 = ~n13408 ;
  assign n13414 = n23354 & n13413 ;
  assign n23355 = ~n13414 ;
  assign n13415 = n13407 & n23355 ;
  assign n13416 = x109 | n13415 ;
  assign n13417 = x109 & n13415 ;
  assign n23356 = ~n12931 ;
  assign n13418 = n23356 & n12932 ;
  assign n13419 = n139 & n13418 ;
  assign n13420 = n12937 & n13419 ;
  assign n13421 = n12937 | n13419 ;
  assign n23357 = ~n13420 ;
  assign n13422 = n23357 & n13421 ;
  assign n23358 = ~n13417 ;
  assign n13423 = n23358 & n13422 ;
  assign n23359 = ~n13423 ;
  assign n13424 = n13416 & n23359 ;
  assign n13425 = x110 | n13424 ;
  assign n13426 = x110 & n13424 ;
  assign n23360 = ~n12940 ;
  assign n13427 = n23360 & n12941 ;
  assign n13428 = n139 & n13427 ;
  assign n13429 = n23161 & n13428 ;
  assign n23361 = ~n13428 ;
  assign n13430 = n12946 & n23361 ;
  assign n13431 = n13429 | n13430 ;
  assign n23362 = ~n13426 ;
  assign n13432 = n23362 & n13431 ;
  assign n23363 = ~n13432 ;
  assign n13433 = n13425 & n23363 ;
  assign n13434 = x111 | n13433 ;
  assign n13435 = x111 & n13433 ;
  assign n23364 = ~n12949 ;
  assign n13436 = n23364 & n12950 ;
  assign n13437 = n139 & n13436 ;
  assign n13438 = n23164 & n13437 ;
  assign n23365 = ~n13437 ;
  assign n13439 = n12955 & n23365 ;
  assign n13440 = n13438 | n13439 ;
  assign n23366 = ~n13435 ;
  assign n13441 = n23366 & n13440 ;
  assign n23367 = ~n13441 ;
  assign n13442 = n13434 & n23367 ;
  assign n13443 = x112 | n13442 ;
  assign n13444 = x112 & n13442 ;
  assign n23368 = ~n12958 ;
  assign n13445 = n23368 & n12959 ;
  assign n13446 = n139 & n13445 ;
  assign n13447 = n12964 & n13446 ;
  assign n13448 = n12964 | n13446 ;
  assign n23369 = ~n13447 ;
  assign n13449 = n23369 & n13448 ;
  assign n23370 = ~n13444 ;
  assign n13450 = n23370 & n13449 ;
  assign n23371 = ~n13450 ;
  assign n13451 = n13443 & n23371 ;
  assign n13452 = x113 | n13451 ;
  assign n13453 = x113 & n13451 ;
  assign n23372 = ~n12967 ;
  assign n13454 = n23372 & n12968 ;
  assign n13455 = n139 & n13454 ;
  assign n13456 = n12973 & n13455 ;
  assign n13457 = n12973 | n13455 ;
  assign n23373 = ~n13456 ;
  assign n13458 = n23373 & n13457 ;
  assign n23374 = ~n13453 ;
  assign n13459 = n23374 & n13458 ;
  assign n23375 = ~n13459 ;
  assign n13460 = n13452 & n23375 ;
  assign n13461 = x114 | n13460 ;
  assign n13462 = x114 & n13460 ;
  assign n23376 = ~n12976 ;
  assign n13463 = n23376 & n12977 ;
  assign n13464 = n139 & n13463 ;
  assign n13465 = n12982 & n13464 ;
  assign n13466 = n12982 | n13464 ;
  assign n23377 = ~n13465 ;
  assign n13467 = n23377 & n13466 ;
  assign n23378 = ~n13462 ;
  assign n13468 = n23378 & n13467 ;
  assign n23379 = ~n13468 ;
  assign n13469 = n13461 & n23379 ;
  assign n13470 = x115 | n13469 ;
  assign n13471 = x115 & n13469 ;
  assign n23380 = ~n12985 ;
  assign n13472 = n23380 & n12986 ;
  assign n13473 = n139 & n13472 ;
  assign n13474 = n23173 & n13473 ;
  assign n23381 = ~n13473 ;
  assign n13475 = n12991 & n23381 ;
  assign n13476 = n13474 | n13475 ;
  assign n23382 = ~n13471 ;
  assign n13477 = n23382 & n13476 ;
  assign n23383 = ~n13477 ;
  assign n13478 = n13470 & n23383 ;
  assign n13479 = x116 | n13478 ;
  assign n13480 = x116 & n13478 ;
  assign n23384 = ~n12994 ;
  assign n13481 = n23384 & n12995 ;
  assign n13482 = n139 & n13481 ;
  assign n13483 = n13000 & n13482 ;
  assign n13484 = n13000 | n13482 ;
  assign n23385 = ~n13483 ;
  assign n13485 = n23385 & n13484 ;
  assign n23386 = ~n13480 ;
  assign n13486 = n23386 & n13485 ;
  assign n23387 = ~n13486 ;
  assign n13487 = n13479 & n23387 ;
  assign n13488 = x117 | n13487 ;
  assign n13489 = x117 & n13487 ;
  assign n23388 = ~n13489 ;
  assign n13490 = n13019 & n23388 ;
  assign n23389 = ~n13490 ;
  assign n13491 = n13488 & n23389 ;
  assign n23390 = ~n13009 ;
  assign n13492 = n13007 & n23390 ;
  assign n23391 = ~n13492 ;
  assign n13493 = n13012 & n23391 ;
  assign n23392 = ~x118 ;
  assign n13494 = n23392 & n13493 ;
  assign n23393 = ~n13494 ;
  assign n13495 = n13491 & n23393 ;
  assign n23394 = ~n13493 ;
  assign n13496 = x118 & n23394 ;
  assign n13497 = n18303 | n13496 ;
  assign n13498 = n13495 | n13497 ;
  assign n13499 = n13488 & n23388 ;
  assign n138 = ~n13498 ;
  assign n13500 = n138 & n13499 ;
  assign n13501 = n13019 & n13500 ;
  assign n13502 = n13019 | n13500 ;
  assign n23396 = ~n13501 ;
  assign n13503 = n23396 & n13502 ;
  assign n23397 = ~x8 ;
  assign n13504 = n23397 & x64 ;
  assign n13506 = x65 | n13504 ;
  assign n13505 = x65 & n13504 ;
  assign n13507 = x64 & n138 ;
  assign n13508 = x9 & n13507 ;
  assign n13509 = x9 | n13507 ;
  assign n23398 = ~n13508 ;
  assign n13510 = n23398 & n13509 ;
  assign n23399 = ~n13505 ;
  assign n13511 = n23399 & n13510 ;
  assign n23400 = ~n13511 ;
  assign n13512 = n13506 & n23400 ;
  assign n13513 = x66 | n13512 ;
  assign n13514 = x66 & n13512 ;
  assign n13515 = n23183 & n13022 ;
  assign n13516 = n138 & n13515 ;
  assign n13517 = n13026 & n13516 ;
  assign n13518 = n13026 | n13516 ;
  assign n23401 = ~n13517 ;
  assign n13519 = n23401 & n13518 ;
  assign n23402 = ~n13514 ;
  assign n13520 = n23402 & n13519 ;
  assign n23403 = ~n13520 ;
  assign n13521 = n13513 & n23403 ;
  assign n13522 = x67 | n13521 ;
  assign n13523 = x67 & n13521 ;
  assign n13524 = n13029 & n23186 ;
  assign n13525 = n138 & n13524 ;
  assign n23404 = ~n13035 ;
  assign n13526 = n23404 & n13525 ;
  assign n23405 = ~n13525 ;
  assign n13527 = n13035 & n23405 ;
  assign n13528 = n13526 | n13527 ;
  assign n23406 = ~n13523 ;
  assign n13529 = n23406 & n13528 ;
  assign n23407 = ~n13529 ;
  assign n13530 = n13522 & n23407 ;
  assign n13531 = x68 | n13530 ;
  assign n13532 = x68 & n13530 ;
  assign n13533 = n13038 & n23190 ;
  assign n13534 = n138 & n13533 ;
  assign n23408 = ~n13044 ;
  assign n13535 = n23408 & n13534 ;
  assign n23409 = ~n13534 ;
  assign n13536 = n13044 & n23409 ;
  assign n13537 = n13535 | n13536 ;
  assign n23410 = ~n13532 ;
  assign n13538 = n23410 & n13537 ;
  assign n23411 = ~n13538 ;
  assign n13539 = n13531 & n23411 ;
  assign n13540 = x69 | n13539 ;
  assign n13541 = x69 & n13539 ;
  assign n13542 = n13047 & n23194 ;
  assign n13543 = n138 & n13542 ;
  assign n13544 = n13053 & n13543 ;
  assign n13545 = n13053 | n13543 ;
  assign n23412 = ~n13544 ;
  assign n13546 = n23412 & n13545 ;
  assign n23413 = ~n13541 ;
  assign n13547 = n23413 & n13546 ;
  assign n23414 = ~n13547 ;
  assign n13548 = n13540 & n23414 ;
  assign n13549 = x70 | n13548 ;
  assign n13550 = x70 & n13548 ;
  assign n13551 = n13056 & n23198 ;
  assign n13552 = n138 & n13551 ;
  assign n23415 = ~n13062 ;
  assign n13553 = n23415 & n13552 ;
  assign n23416 = ~n13552 ;
  assign n13554 = n13062 & n23416 ;
  assign n13555 = n13553 | n13554 ;
  assign n23417 = ~n13550 ;
  assign n13556 = n23417 & n13555 ;
  assign n23418 = ~n13556 ;
  assign n13557 = n13549 & n23418 ;
  assign n13558 = x71 | n13557 ;
  assign n13559 = x71 & n13557 ;
  assign n13560 = n13065 & n23202 ;
  assign n13561 = n138 & n13560 ;
  assign n13562 = n13071 & n13561 ;
  assign n13563 = n13071 | n13561 ;
  assign n23419 = ~n13562 ;
  assign n13564 = n23419 & n13563 ;
  assign n23420 = ~n13559 ;
  assign n13565 = n23420 & n13564 ;
  assign n23421 = ~n13565 ;
  assign n13566 = n13558 & n23421 ;
  assign n13567 = x72 | n13566 ;
  assign n13568 = x72 & n13566 ;
  assign n13569 = n13074 & n23206 ;
  assign n13570 = n138 & n13569 ;
  assign n13571 = n13080 & n13570 ;
  assign n13572 = n13080 | n13570 ;
  assign n23422 = ~n13571 ;
  assign n13573 = n23422 & n13572 ;
  assign n23423 = ~n13568 ;
  assign n13574 = n23423 & n13573 ;
  assign n23424 = ~n13574 ;
  assign n13575 = n13567 & n23424 ;
  assign n13576 = x73 | n13575 ;
  assign n13577 = x73 & n13575 ;
  assign n13578 = n13083 & n23210 ;
  assign n13579 = n138 & n13578 ;
  assign n13580 = n13089 & n13579 ;
  assign n13581 = n13089 | n13579 ;
  assign n23425 = ~n13580 ;
  assign n13582 = n23425 & n13581 ;
  assign n23426 = ~n13577 ;
  assign n13583 = n23426 & n13582 ;
  assign n23427 = ~n13583 ;
  assign n13584 = n13576 & n23427 ;
  assign n13585 = x74 | n13584 ;
  assign n13586 = x74 & n13584 ;
  assign n13587 = n13092 & n23214 ;
  assign n13588 = n138 & n13587 ;
  assign n23428 = ~n13098 ;
  assign n13589 = n23428 & n13588 ;
  assign n23429 = ~n13588 ;
  assign n13590 = n13098 & n23429 ;
  assign n13591 = n13589 | n13590 ;
  assign n23430 = ~n13586 ;
  assign n13592 = n23430 & n13591 ;
  assign n23431 = ~n13592 ;
  assign n13593 = n13585 & n23431 ;
  assign n13594 = x75 | n13593 ;
  assign n13595 = x75 & n13593 ;
  assign n13596 = n13101 & n23218 ;
  assign n13597 = n138 & n13596 ;
  assign n23432 = ~n13107 ;
  assign n13598 = n23432 & n13597 ;
  assign n23433 = ~n13597 ;
  assign n13599 = n13107 & n23433 ;
  assign n13600 = n13598 | n13599 ;
  assign n23434 = ~n13595 ;
  assign n13601 = n23434 & n13600 ;
  assign n23435 = ~n13601 ;
  assign n13602 = n13594 & n23435 ;
  assign n13603 = x76 | n13602 ;
  assign n13604 = x76 & n13602 ;
  assign n13605 = n13110 & n23222 ;
  assign n13606 = n138 & n13605 ;
  assign n23436 = ~n13116 ;
  assign n13607 = n23436 & n13606 ;
  assign n23437 = ~n13606 ;
  assign n13608 = n13116 & n23437 ;
  assign n13609 = n13607 | n13608 ;
  assign n23438 = ~n13604 ;
  assign n13610 = n23438 & n13609 ;
  assign n23439 = ~n13610 ;
  assign n13611 = n13603 & n23439 ;
  assign n13612 = x77 | n13611 ;
  assign n13613 = x77 & n13611 ;
  assign n13614 = n13119 & n23226 ;
  assign n13615 = n138 & n13614 ;
  assign n13616 = n13125 & n13615 ;
  assign n13617 = n13125 | n13615 ;
  assign n23440 = ~n13616 ;
  assign n13618 = n23440 & n13617 ;
  assign n23441 = ~n13613 ;
  assign n13619 = n23441 & n13618 ;
  assign n23442 = ~n13619 ;
  assign n13620 = n13612 & n23442 ;
  assign n13621 = x78 | n13620 ;
  assign n13622 = x78 & n13620 ;
  assign n13623 = n13128 & n23230 ;
  assign n13624 = n138 & n13623 ;
  assign n23443 = ~n13134 ;
  assign n13625 = n23443 & n13624 ;
  assign n23444 = ~n13624 ;
  assign n13626 = n13134 & n23444 ;
  assign n13627 = n13625 | n13626 ;
  assign n23445 = ~n13622 ;
  assign n13628 = n23445 & n13627 ;
  assign n23446 = ~n13628 ;
  assign n13629 = n13621 & n23446 ;
  assign n13630 = x79 | n13629 ;
  assign n13631 = x79 & n13629 ;
  assign n13632 = n13137 & n23234 ;
  assign n13633 = n138 & n13632 ;
  assign n23447 = ~n13143 ;
  assign n13634 = n23447 & n13633 ;
  assign n23448 = ~n13633 ;
  assign n13635 = n13143 & n23448 ;
  assign n13636 = n13634 | n13635 ;
  assign n23449 = ~n13631 ;
  assign n13637 = n23449 & n13636 ;
  assign n23450 = ~n13637 ;
  assign n13638 = n13630 & n23450 ;
  assign n13639 = x80 | n13638 ;
  assign n13640 = x80 & n13638 ;
  assign n13641 = n13146 & n23238 ;
  assign n13642 = n138 & n13641 ;
  assign n23451 = ~n13152 ;
  assign n13643 = n23451 & n13642 ;
  assign n23452 = ~n13642 ;
  assign n13644 = n13152 & n23452 ;
  assign n13645 = n13643 | n13644 ;
  assign n23453 = ~n13640 ;
  assign n13646 = n23453 & n13645 ;
  assign n23454 = ~n13646 ;
  assign n13647 = n13639 & n23454 ;
  assign n13648 = x81 | n13647 ;
  assign n13649 = x81 & n13647 ;
  assign n13650 = n13155 & n23242 ;
  assign n13651 = n138 & n13650 ;
  assign n13652 = n13161 & n13651 ;
  assign n13653 = n13161 | n13651 ;
  assign n23455 = ~n13652 ;
  assign n13654 = n23455 & n13653 ;
  assign n23456 = ~n13649 ;
  assign n13655 = n23456 & n13654 ;
  assign n23457 = ~n13655 ;
  assign n13656 = n13648 & n23457 ;
  assign n13657 = x82 | n13656 ;
  assign n13658 = x82 & n13656 ;
  assign n13659 = n13164 & n23246 ;
  assign n13660 = n138 & n13659 ;
  assign n23458 = ~n13170 ;
  assign n13661 = n23458 & n13660 ;
  assign n23459 = ~n13660 ;
  assign n13662 = n13170 & n23459 ;
  assign n13663 = n13661 | n13662 ;
  assign n23460 = ~n13658 ;
  assign n13664 = n23460 & n13663 ;
  assign n23461 = ~n13664 ;
  assign n13665 = n13657 & n23461 ;
  assign n13666 = x83 | n13665 ;
  assign n13667 = x83 & n13665 ;
  assign n13668 = n13173 & n23250 ;
  assign n13669 = n138 & n13668 ;
  assign n23462 = ~n13179 ;
  assign n13670 = n23462 & n13669 ;
  assign n23463 = ~n13669 ;
  assign n13671 = n13179 & n23463 ;
  assign n13672 = n13670 | n13671 ;
  assign n23464 = ~n13667 ;
  assign n13673 = n23464 & n13672 ;
  assign n23465 = ~n13673 ;
  assign n13674 = n13666 & n23465 ;
  assign n13675 = x84 | n13674 ;
  assign n13676 = x84 & n13674 ;
  assign n13677 = n13182 & n23254 ;
  assign n13678 = n138 & n13677 ;
  assign n23466 = ~n13188 ;
  assign n13679 = n23466 & n13678 ;
  assign n23467 = ~n13678 ;
  assign n13680 = n13188 & n23467 ;
  assign n13681 = n13679 | n13680 ;
  assign n23468 = ~n13676 ;
  assign n13682 = n23468 & n13681 ;
  assign n23469 = ~n13682 ;
  assign n13683 = n13675 & n23469 ;
  assign n13684 = x85 | n13683 ;
  assign n13685 = x85 & n13683 ;
  assign n13686 = n13191 & n23258 ;
  assign n13687 = n138 & n13686 ;
  assign n23470 = ~n13197 ;
  assign n13688 = n23470 & n13687 ;
  assign n23471 = ~n13687 ;
  assign n13689 = n13197 & n23471 ;
  assign n13690 = n13688 | n13689 ;
  assign n23472 = ~n13685 ;
  assign n13691 = n23472 & n13690 ;
  assign n23473 = ~n13691 ;
  assign n13692 = n13684 & n23473 ;
  assign n13693 = x86 | n13692 ;
  assign n13694 = x86 & n13692 ;
  assign n13695 = n13200 & n23262 ;
  assign n13696 = n138 & n13695 ;
  assign n23474 = ~n13206 ;
  assign n13697 = n23474 & n13696 ;
  assign n23475 = ~n13696 ;
  assign n13698 = n13206 & n23475 ;
  assign n13699 = n13697 | n13698 ;
  assign n23476 = ~n13694 ;
  assign n13700 = n23476 & n13699 ;
  assign n23477 = ~n13700 ;
  assign n13701 = n13693 & n23477 ;
  assign n13702 = x87 | n13701 ;
  assign n13703 = x87 & n13701 ;
  assign n13704 = n13209 & n23266 ;
  assign n13705 = n138 & n13704 ;
  assign n23478 = ~n13215 ;
  assign n13706 = n23478 & n13705 ;
  assign n23479 = ~n13705 ;
  assign n13707 = n13215 & n23479 ;
  assign n13708 = n13706 | n13707 ;
  assign n23480 = ~n13703 ;
  assign n13709 = n23480 & n13708 ;
  assign n23481 = ~n13709 ;
  assign n13710 = n13702 & n23481 ;
  assign n13711 = x88 | n13710 ;
  assign n13712 = x88 & n13710 ;
  assign n13713 = n13218 & n23270 ;
  assign n13714 = n138 & n13713 ;
  assign n13715 = n13224 & n13714 ;
  assign n13716 = n13224 | n13714 ;
  assign n23482 = ~n13715 ;
  assign n13717 = n23482 & n13716 ;
  assign n23483 = ~n13712 ;
  assign n13718 = n23483 & n13717 ;
  assign n23484 = ~n13718 ;
  assign n13719 = n13711 & n23484 ;
  assign n13720 = x89 | n13719 ;
  assign n13721 = x89 & n13719 ;
  assign n13722 = n13227 & n23274 ;
  assign n13723 = n138 & n13722 ;
  assign n23485 = ~n13233 ;
  assign n13724 = n23485 & n13723 ;
  assign n23486 = ~n13723 ;
  assign n13725 = n13233 & n23486 ;
  assign n13726 = n13724 | n13725 ;
  assign n23487 = ~n13721 ;
  assign n13727 = n23487 & n13726 ;
  assign n23488 = ~n13727 ;
  assign n13728 = n13720 & n23488 ;
  assign n13729 = x90 | n13728 ;
  assign n13730 = x90 & n13728 ;
  assign n13731 = n13236 & n23278 ;
  assign n13732 = n138 & n13731 ;
  assign n23489 = ~n13242 ;
  assign n13733 = n23489 & n13732 ;
  assign n23490 = ~n13732 ;
  assign n13734 = n13242 & n23490 ;
  assign n13735 = n13733 | n13734 ;
  assign n23491 = ~n13730 ;
  assign n13736 = n23491 & n13735 ;
  assign n23492 = ~n13736 ;
  assign n13737 = n13729 & n23492 ;
  assign n13738 = x91 | n13737 ;
  assign n13739 = x91 & n13737 ;
  assign n13740 = n13245 & n23282 ;
  assign n13741 = n138 & n13740 ;
  assign n23493 = ~n13251 ;
  assign n13742 = n23493 & n13741 ;
  assign n23494 = ~n13741 ;
  assign n13743 = n13251 & n23494 ;
  assign n13744 = n13742 | n13743 ;
  assign n23495 = ~n13739 ;
  assign n13745 = n23495 & n13744 ;
  assign n23496 = ~n13745 ;
  assign n13746 = n13738 & n23496 ;
  assign n13747 = x92 | n13746 ;
  assign n13748 = x92 & n13746 ;
  assign n13749 = n13254 & n23286 ;
  assign n13750 = n138 & n13749 ;
  assign n23497 = ~n13260 ;
  assign n13751 = n23497 & n13750 ;
  assign n23498 = ~n13750 ;
  assign n13752 = n13260 & n23498 ;
  assign n13753 = n13751 | n13752 ;
  assign n23499 = ~n13748 ;
  assign n13754 = n23499 & n13753 ;
  assign n23500 = ~n13754 ;
  assign n13755 = n13747 & n23500 ;
  assign n13756 = x93 | n13755 ;
  assign n13757 = x93 & n13755 ;
  assign n13758 = n13263 & n23290 ;
  assign n13759 = n138 & n13758 ;
  assign n23501 = ~n13269 ;
  assign n13760 = n23501 & n13759 ;
  assign n23502 = ~n13759 ;
  assign n13761 = n13269 & n23502 ;
  assign n13762 = n13760 | n13761 ;
  assign n23503 = ~n13757 ;
  assign n13763 = n23503 & n13762 ;
  assign n23504 = ~n13763 ;
  assign n13764 = n13756 & n23504 ;
  assign n13765 = x94 | n13764 ;
  assign n13766 = x94 & n13764 ;
  assign n13767 = n13272 & n23294 ;
  assign n13768 = n138 & n13767 ;
  assign n13769 = n13278 & n13768 ;
  assign n13770 = n13278 | n13768 ;
  assign n23505 = ~n13769 ;
  assign n13771 = n23505 & n13770 ;
  assign n23506 = ~n13766 ;
  assign n13772 = n23506 & n13771 ;
  assign n23507 = ~n13772 ;
  assign n13773 = n13765 & n23507 ;
  assign n13774 = x95 | n13773 ;
  assign n13775 = x95 & n13773 ;
  assign n13776 = n13281 & n23298 ;
  assign n13777 = n138 & n13776 ;
  assign n23508 = ~n13287 ;
  assign n13778 = n23508 & n13777 ;
  assign n23509 = ~n13777 ;
  assign n13779 = n13287 & n23509 ;
  assign n13780 = n13778 | n13779 ;
  assign n23510 = ~n13775 ;
  assign n13781 = n23510 & n13780 ;
  assign n23511 = ~n13781 ;
  assign n13782 = n13774 & n23511 ;
  assign n13783 = x96 | n13782 ;
  assign n13784 = x96 & n13782 ;
  assign n13785 = n13290 & n23302 ;
  assign n13786 = n138 & n13785 ;
  assign n23512 = ~n13296 ;
  assign n13787 = n23512 & n13786 ;
  assign n23513 = ~n13786 ;
  assign n13788 = n13296 & n23513 ;
  assign n13789 = n13787 | n13788 ;
  assign n23514 = ~n13784 ;
  assign n13790 = n23514 & n13789 ;
  assign n23515 = ~n13790 ;
  assign n13791 = n13783 & n23515 ;
  assign n13792 = x97 | n13791 ;
  assign n13793 = x97 & n13791 ;
  assign n13794 = n13299 & n23306 ;
  assign n13795 = n138 & n13794 ;
  assign n13796 = n13305 & n13795 ;
  assign n13797 = n13305 | n13795 ;
  assign n23516 = ~n13796 ;
  assign n13798 = n23516 & n13797 ;
  assign n23517 = ~n13793 ;
  assign n13799 = n23517 & n13798 ;
  assign n23518 = ~n13799 ;
  assign n13800 = n13792 & n23518 ;
  assign n13801 = x98 | n13800 ;
  assign n13802 = x98 & n13800 ;
  assign n13803 = n13308 & n23310 ;
  assign n13804 = n138 & n13803 ;
  assign n23519 = ~n13314 ;
  assign n13805 = n23519 & n13804 ;
  assign n23520 = ~n13804 ;
  assign n13806 = n13314 & n23520 ;
  assign n13807 = n13805 | n13806 ;
  assign n23521 = ~n13802 ;
  assign n13808 = n23521 & n13807 ;
  assign n23522 = ~n13808 ;
  assign n13809 = n13801 & n23522 ;
  assign n13810 = x99 | n13809 ;
  assign n13811 = x99 & n13809 ;
  assign n13812 = n13317 & n23314 ;
  assign n13813 = n138 & n13812 ;
  assign n23523 = ~n13323 ;
  assign n13814 = n23523 & n13813 ;
  assign n23524 = ~n13813 ;
  assign n13815 = n13323 & n23524 ;
  assign n13816 = n13814 | n13815 ;
  assign n23525 = ~n13811 ;
  assign n13817 = n23525 & n13816 ;
  assign n23526 = ~n13817 ;
  assign n13818 = n13810 & n23526 ;
  assign n13819 = x100 | n13818 ;
  assign n13820 = x100 & n13818 ;
  assign n13821 = n13326 & n23318 ;
  assign n13822 = n138 & n13821 ;
  assign n23527 = ~n13332 ;
  assign n13823 = n23527 & n13822 ;
  assign n23528 = ~n13822 ;
  assign n13824 = n13332 & n23528 ;
  assign n13825 = n13823 | n13824 ;
  assign n23529 = ~n13820 ;
  assign n13826 = n23529 & n13825 ;
  assign n23530 = ~n13826 ;
  assign n13827 = n13819 & n23530 ;
  assign n13828 = x101 | n13827 ;
  assign n13829 = x101 & n13827 ;
  assign n13830 = n13335 & n23322 ;
  assign n13831 = n138 & n13830 ;
  assign n23531 = ~n13341 ;
  assign n13832 = n23531 & n13831 ;
  assign n23532 = ~n13831 ;
  assign n13833 = n13341 & n23532 ;
  assign n13834 = n13832 | n13833 ;
  assign n23533 = ~n13829 ;
  assign n13835 = n23533 & n13834 ;
  assign n23534 = ~n13835 ;
  assign n13836 = n13828 & n23534 ;
  assign n13837 = x102 | n13836 ;
  assign n13838 = x102 & n13836 ;
  assign n13839 = n13344 & n23326 ;
  assign n13840 = n138 & n13839 ;
  assign n23535 = ~n13350 ;
  assign n13841 = n23535 & n13840 ;
  assign n23536 = ~n13840 ;
  assign n13842 = n13350 & n23536 ;
  assign n13843 = n13841 | n13842 ;
  assign n23537 = ~n13838 ;
  assign n13844 = n23537 & n13843 ;
  assign n23538 = ~n13844 ;
  assign n13845 = n13837 & n23538 ;
  assign n13846 = x103 | n13845 ;
  assign n13847 = x103 & n13845 ;
  assign n13848 = n13353 & n23330 ;
  assign n13849 = n138 & n13848 ;
  assign n13850 = n13359 & n13849 ;
  assign n13851 = n13359 | n13849 ;
  assign n23539 = ~n13850 ;
  assign n13852 = n23539 & n13851 ;
  assign n23540 = ~n13847 ;
  assign n13853 = n23540 & n13852 ;
  assign n23541 = ~n13853 ;
  assign n13854 = n13846 & n23541 ;
  assign n13855 = x104 | n13854 ;
  assign n13856 = x104 & n13854 ;
  assign n13857 = n13362 & n23334 ;
  assign n13858 = n138 & n13857 ;
  assign n23542 = ~n13368 ;
  assign n13859 = n23542 & n13858 ;
  assign n23543 = ~n13858 ;
  assign n13860 = n13368 & n23543 ;
  assign n13861 = n13859 | n13860 ;
  assign n23544 = ~n13856 ;
  assign n13862 = n23544 & n13861 ;
  assign n23545 = ~n13862 ;
  assign n13863 = n13855 & n23545 ;
  assign n13864 = x105 | n13863 ;
  assign n13865 = x105 & n13863 ;
  assign n13866 = n13371 & n23338 ;
  assign n13867 = n138 & n13866 ;
  assign n23546 = ~n13377 ;
  assign n13868 = n23546 & n13867 ;
  assign n23547 = ~n13867 ;
  assign n13869 = n13377 & n23547 ;
  assign n13870 = n13868 | n13869 ;
  assign n23548 = ~n13865 ;
  assign n13871 = n23548 & n13870 ;
  assign n23549 = ~n13871 ;
  assign n13872 = n13864 & n23549 ;
  assign n13873 = x106 | n13872 ;
  assign n13874 = x106 & n13872 ;
  assign n13875 = n13380 & n23342 ;
  assign n13876 = n138 & n13875 ;
  assign n23550 = ~n13386 ;
  assign n13877 = n23550 & n13876 ;
  assign n23551 = ~n13876 ;
  assign n13878 = n13386 & n23551 ;
  assign n13879 = n13877 | n13878 ;
  assign n23552 = ~n13874 ;
  assign n13880 = n23552 & n13879 ;
  assign n23553 = ~n13880 ;
  assign n13881 = n13873 & n23553 ;
  assign n13882 = x107 | n13881 ;
  assign n13883 = x107 & n13881 ;
  assign n13884 = n13389 & n23346 ;
  assign n13885 = n138 & n13884 ;
  assign n23554 = ~n13395 ;
  assign n13886 = n23554 & n13885 ;
  assign n23555 = ~n13885 ;
  assign n13887 = n13395 & n23555 ;
  assign n13888 = n13886 | n13887 ;
  assign n23556 = ~n13883 ;
  assign n13889 = n23556 & n13888 ;
  assign n23557 = ~n13889 ;
  assign n13890 = n13882 & n23557 ;
  assign n13891 = x108 | n13890 ;
  assign n13892 = x108 & n13890 ;
  assign n13893 = n13398 & n23350 ;
  assign n13894 = n138 & n13893 ;
  assign n13895 = n13404 & n13894 ;
  assign n13896 = n13404 | n13894 ;
  assign n23558 = ~n13895 ;
  assign n13897 = n23558 & n13896 ;
  assign n23559 = ~n13892 ;
  assign n13898 = n23559 & n13897 ;
  assign n23560 = ~n13898 ;
  assign n13899 = n13891 & n23560 ;
  assign n13900 = x109 | n13899 ;
  assign n13901 = x109 & n13899 ;
  assign n13902 = n13407 & n23354 ;
  assign n13903 = n138 & n13902 ;
  assign n13904 = n13413 & n13903 ;
  assign n13905 = n13413 | n13903 ;
  assign n23561 = ~n13904 ;
  assign n13906 = n23561 & n13905 ;
  assign n23562 = ~n13901 ;
  assign n13907 = n23562 & n13906 ;
  assign n23563 = ~n13907 ;
  assign n13908 = n13900 & n23563 ;
  assign n13909 = x110 | n13908 ;
  assign n13910 = x110 & n13908 ;
  assign n13911 = n13416 & n23358 ;
  assign n13912 = n138 & n13911 ;
  assign n13913 = n13422 & n13912 ;
  assign n13914 = n13422 | n13912 ;
  assign n23564 = ~n13913 ;
  assign n13915 = n23564 & n13914 ;
  assign n23565 = ~n13910 ;
  assign n13916 = n23565 & n13915 ;
  assign n23566 = ~n13916 ;
  assign n13917 = n13909 & n23566 ;
  assign n13918 = x111 | n13917 ;
  assign n13919 = x111 & n13917 ;
  assign n13920 = n13425 & n23362 ;
  assign n13921 = n138 & n13920 ;
  assign n23567 = ~n13431 ;
  assign n13922 = n23567 & n13921 ;
  assign n23568 = ~n13921 ;
  assign n13923 = n13431 & n23568 ;
  assign n13924 = n13922 | n13923 ;
  assign n23569 = ~n13919 ;
  assign n13925 = n23569 & n13924 ;
  assign n23570 = ~n13925 ;
  assign n13926 = n13918 & n23570 ;
  assign n13927 = x112 | n13926 ;
  assign n13928 = x112 & n13926 ;
  assign n13929 = n13434 & n23366 ;
  assign n13930 = n138 & n13929 ;
  assign n23571 = ~n13440 ;
  assign n13931 = n23571 & n13930 ;
  assign n23572 = ~n13930 ;
  assign n13932 = n13440 & n23572 ;
  assign n13933 = n13931 | n13932 ;
  assign n23573 = ~n13928 ;
  assign n13934 = n23573 & n13933 ;
  assign n23574 = ~n13934 ;
  assign n13935 = n13927 & n23574 ;
  assign n13936 = x113 | n13935 ;
  assign n13937 = x113 & n13935 ;
  assign n13938 = n13443 & n23370 ;
  assign n13939 = n138 & n13938 ;
  assign n23575 = ~n13449 ;
  assign n13940 = n23575 & n13939 ;
  assign n23576 = ~n13939 ;
  assign n13941 = n13449 & n23576 ;
  assign n13942 = n13940 | n13941 ;
  assign n23577 = ~n13937 ;
  assign n13943 = n23577 & n13942 ;
  assign n23578 = ~n13943 ;
  assign n13944 = n13936 & n23578 ;
  assign n13945 = x114 | n13944 ;
  assign n13946 = x114 & n13944 ;
  assign n13947 = n13452 & n23374 ;
  assign n13948 = n138 & n13947 ;
  assign n23579 = ~n13458 ;
  assign n13949 = n23579 & n13948 ;
  assign n23580 = ~n13948 ;
  assign n13950 = n13458 & n23580 ;
  assign n13951 = n13949 | n13950 ;
  assign n23581 = ~n13946 ;
  assign n13952 = n23581 & n13951 ;
  assign n23582 = ~n13952 ;
  assign n13953 = n13945 & n23582 ;
  assign n13954 = x115 | n13953 ;
  assign n13955 = x115 & n13953 ;
  assign n13956 = n13461 & n23378 ;
  assign n13957 = n138 & n13956 ;
  assign n23583 = ~n13467 ;
  assign n13958 = n23583 & n13957 ;
  assign n23584 = ~n13957 ;
  assign n13959 = n13467 & n23584 ;
  assign n13960 = n13958 | n13959 ;
  assign n23585 = ~n13955 ;
  assign n13961 = n23585 & n13960 ;
  assign n23586 = ~n13961 ;
  assign n13962 = n13954 & n23586 ;
  assign n13963 = x116 | n13962 ;
  assign n13964 = x116 & n13962 ;
  assign n13965 = n13470 & n23382 ;
  assign n13966 = n138 & n13965 ;
  assign n23587 = ~n13476 ;
  assign n13967 = n23587 & n13966 ;
  assign n23588 = ~n13966 ;
  assign n13968 = n13476 & n23588 ;
  assign n13969 = n13967 | n13968 ;
  assign n23589 = ~n13964 ;
  assign n13970 = n23589 & n13969 ;
  assign n23590 = ~n13970 ;
  assign n13971 = n13963 & n23590 ;
  assign n13972 = x117 | n13971 ;
  assign n13973 = x117 & n13971 ;
  assign n13974 = n13479 & n23386 ;
  assign n13975 = n138 & n13974 ;
  assign n23591 = ~n13485 ;
  assign n13976 = n23591 & n13975 ;
  assign n23592 = ~n13975 ;
  assign n13977 = n13485 & n23592 ;
  assign n13978 = n13976 | n13977 ;
  assign n23593 = ~n13973 ;
  assign n13979 = n23593 & n13978 ;
  assign n23594 = ~n13979 ;
  assign n13980 = n13972 & n23594 ;
  assign n13981 = x118 | n13980 ;
  assign n13982 = x118 & n13980 ;
  assign n23595 = ~n13982 ;
  assign n13983 = n13503 & n23595 ;
  assign n23596 = ~n13983 ;
  assign n13984 = n13981 & n23596 ;
  assign n13985 = x118 & n13491 ;
  assign n13986 = x118 | n13491 ;
  assign n23597 = ~n18303 ;
  assign n13987 = n23597 & n13986 ;
  assign n23598 = ~n13985 ;
  assign n13988 = n23598 & n13987 ;
  assign n23599 = ~n13988 ;
  assign n13989 = n13493 & n23599 ;
  assign n23600 = ~x119 ;
  assign n13991 = n23600 & n13989 ;
  assign n23601 = ~n13991 ;
  assign n13992 = n13984 & n23601 ;
  assign n23602 = ~n13989 ;
  assign n13990 = x119 & n23602 ;
  assign n13993 = n18298 | n13990 ;
  assign n13994 = n13992 | n13993 ;
  assign n13996 = n13981 & n23595 ;
  assign n137 = ~n13994 ;
  assign n13997 = n137 & n13996 ;
  assign n23604 = ~n13503 ;
  assign n13998 = n23604 & n13997 ;
  assign n23605 = ~n13997 ;
  assign n13999 = n13503 & n23605 ;
  assign n14000 = n13998 | n13999 ;
  assign n23606 = ~x7 ;
  assign n14001 = n23606 & x64 ;
  assign n14002 = x65 | n14001 ;
  assign n13995 = n13504 & n137 ;
  assign n14004 = x64 & n137 ;
  assign n23607 = ~n14004 ;
  assign n14005 = x8 & n23607 ;
  assign n14006 = n13995 | n14005 ;
  assign n14007 = x65 & n14001 ;
  assign n23608 = ~n14007 ;
  assign n14008 = n14006 & n23608 ;
  assign n23609 = ~n14008 ;
  assign n14009 = n14002 & n23609 ;
  assign n14010 = x66 & n14009 ;
  assign n14011 = n23399 & n13506 ;
  assign n14012 = n137 & n14011 ;
  assign n14013 = n13510 & n14012 ;
  assign n14014 = n13510 | n14012 ;
  assign n23610 = ~n14013 ;
  assign n14015 = n23610 & n14014 ;
  assign n14016 = x66 | n14009 ;
  assign n23611 = ~n14015 ;
  assign n14017 = n23611 & n14016 ;
  assign n14018 = n14010 | n14017 ;
  assign n14019 = x67 & n14018 ;
  assign n14020 = x67 | n14018 ;
  assign n14021 = n13513 & n23402 ;
  assign n14022 = n137 & n14021 ;
  assign n23612 = ~n13519 ;
  assign n14023 = n23612 & n14022 ;
  assign n23613 = ~n14022 ;
  assign n14024 = n13519 & n23613 ;
  assign n14025 = n14023 | n14024 ;
  assign n23614 = ~n14025 ;
  assign n14026 = n14020 & n23614 ;
  assign n14027 = n14019 | n14026 ;
  assign n14028 = x68 & n14027 ;
  assign n14029 = x68 | n14027 ;
  assign n14030 = n13522 & n23406 ;
  assign n14031 = n137 & n14030 ;
  assign n23615 = ~n13528 ;
  assign n14032 = n23615 & n14031 ;
  assign n23616 = ~n14031 ;
  assign n14033 = n13528 & n23616 ;
  assign n14034 = n14032 | n14033 ;
  assign n23617 = ~n14034 ;
  assign n14035 = n14029 & n23617 ;
  assign n14036 = n14028 | n14035 ;
  assign n14037 = x69 & n14036 ;
  assign n14038 = x69 | n14036 ;
  assign n14039 = n13531 & n23410 ;
  assign n14040 = n137 & n14039 ;
  assign n23618 = ~n13537 ;
  assign n14041 = n23618 & n14040 ;
  assign n23619 = ~n14040 ;
  assign n14042 = n13537 & n23619 ;
  assign n14043 = n14041 | n14042 ;
  assign n23620 = ~n14043 ;
  assign n14044 = n14038 & n23620 ;
  assign n14045 = n14037 | n14044 ;
  assign n14046 = x70 & n14045 ;
  assign n14047 = x70 | n14045 ;
  assign n14048 = n13540 & n23413 ;
  assign n14049 = n137 & n14048 ;
  assign n14050 = n13546 & n14049 ;
  assign n14051 = n13546 | n14049 ;
  assign n23621 = ~n14050 ;
  assign n14052 = n23621 & n14051 ;
  assign n23622 = ~n14052 ;
  assign n14053 = n14047 & n23622 ;
  assign n14054 = n14046 | n14053 ;
  assign n14055 = x71 & n14054 ;
  assign n14056 = x71 | n14054 ;
  assign n14057 = n13549 & n23417 ;
  assign n14058 = n137 & n14057 ;
  assign n23623 = ~n13555 ;
  assign n14059 = n23623 & n14058 ;
  assign n23624 = ~n14058 ;
  assign n14060 = n13555 & n23624 ;
  assign n14061 = n14059 | n14060 ;
  assign n23625 = ~n14061 ;
  assign n14062 = n14056 & n23625 ;
  assign n14063 = n14055 | n14062 ;
  assign n14064 = x72 & n14063 ;
  assign n14065 = x72 | n14063 ;
  assign n14066 = n13558 & n23420 ;
  assign n14067 = n137 & n14066 ;
  assign n23626 = ~n13564 ;
  assign n14068 = n23626 & n14067 ;
  assign n23627 = ~n14067 ;
  assign n14069 = n13564 & n23627 ;
  assign n14070 = n14068 | n14069 ;
  assign n23628 = ~n14070 ;
  assign n14071 = n14065 & n23628 ;
  assign n14072 = n14064 | n14071 ;
  assign n14073 = x73 & n14072 ;
  assign n14074 = x73 | n14072 ;
  assign n14075 = n13567 & n23423 ;
  assign n14076 = n137 & n14075 ;
  assign n14077 = n13573 & n14076 ;
  assign n14078 = n13573 | n14076 ;
  assign n23629 = ~n14077 ;
  assign n14079 = n23629 & n14078 ;
  assign n23630 = ~n14079 ;
  assign n14080 = n14074 & n23630 ;
  assign n14081 = n14073 | n14080 ;
  assign n14082 = x74 & n14081 ;
  assign n14083 = x74 | n14081 ;
  assign n14084 = n13576 & n23426 ;
  assign n14085 = n137 & n14084 ;
  assign n14086 = n13582 & n14085 ;
  assign n14087 = n13582 | n14085 ;
  assign n23631 = ~n14086 ;
  assign n14088 = n23631 & n14087 ;
  assign n23632 = ~n14088 ;
  assign n14089 = n14083 & n23632 ;
  assign n14090 = n14082 | n14089 ;
  assign n14091 = x75 & n14090 ;
  assign n14092 = x75 | n14090 ;
  assign n14093 = n13585 & n23430 ;
  assign n14094 = n137 & n14093 ;
  assign n23633 = ~n13591 ;
  assign n14095 = n23633 & n14094 ;
  assign n23634 = ~n14094 ;
  assign n14096 = n13591 & n23634 ;
  assign n14097 = n14095 | n14096 ;
  assign n23635 = ~n14097 ;
  assign n14098 = n14092 & n23635 ;
  assign n14099 = n14091 | n14098 ;
  assign n14100 = x76 & n14099 ;
  assign n14101 = x76 | n14099 ;
  assign n14102 = n13594 & n23434 ;
  assign n14103 = n137 & n14102 ;
  assign n23636 = ~n13600 ;
  assign n14104 = n23636 & n14103 ;
  assign n23637 = ~n14103 ;
  assign n14105 = n13600 & n23637 ;
  assign n14106 = n14104 | n14105 ;
  assign n23638 = ~n14106 ;
  assign n14107 = n14101 & n23638 ;
  assign n14108 = n14100 | n14107 ;
  assign n14109 = x77 & n14108 ;
  assign n14110 = x77 | n14108 ;
  assign n14111 = n13603 & n23438 ;
  assign n14112 = n137 & n14111 ;
  assign n14113 = n13609 & n14112 ;
  assign n14114 = n13609 | n14112 ;
  assign n23639 = ~n14113 ;
  assign n14115 = n23639 & n14114 ;
  assign n23640 = ~n14115 ;
  assign n14116 = n14110 & n23640 ;
  assign n14117 = n14109 | n14116 ;
  assign n14118 = x78 & n14117 ;
  assign n14119 = x78 | n14117 ;
  assign n14120 = n13612 & n23441 ;
  assign n14121 = n137 & n14120 ;
  assign n23641 = ~n13618 ;
  assign n14122 = n23641 & n14121 ;
  assign n23642 = ~n14121 ;
  assign n14123 = n13618 & n23642 ;
  assign n14124 = n14122 | n14123 ;
  assign n23643 = ~n14124 ;
  assign n14125 = n14119 & n23643 ;
  assign n14126 = n14118 | n14125 ;
  assign n14127 = x79 & n14126 ;
  assign n14128 = x79 | n14126 ;
  assign n14129 = n13621 & n23445 ;
  assign n14130 = n137 & n14129 ;
  assign n14131 = n13627 & n14130 ;
  assign n14132 = n13627 | n14130 ;
  assign n23644 = ~n14131 ;
  assign n14133 = n23644 & n14132 ;
  assign n23645 = ~n14133 ;
  assign n14134 = n14128 & n23645 ;
  assign n14135 = n14127 | n14134 ;
  assign n14136 = x80 & n14135 ;
  assign n14137 = x80 | n14135 ;
  assign n14138 = n13630 & n23449 ;
  assign n14139 = n137 & n14138 ;
  assign n23646 = ~n13636 ;
  assign n14140 = n23646 & n14139 ;
  assign n23647 = ~n14139 ;
  assign n14141 = n13636 & n23647 ;
  assign n14142 = n14140 | n14141 ;
  assign n23648 = ~n14142 ;
  assign n14143 = n14137 & n23648 ;
  assign n14144 = n14136 | n14143 ;
  assign n14145 = x81 & n14144 ;
  assign n14146 = x81 | n14144 ;
  assign n14147 = n13639 & n23453 ;
  assign n14148 = n137 & n14147 ;
  assign n23649 = ~n13645 ;
  assign n14149 = n23649 & n14148 ;
  assign n23650 = ~n14148 ;
  assign n14150 = n13645 & n23650 ;
  assign n14151 = n14149 | n14150 ;
  assign n23651 = ~n14151 ;
  assign n14152 = n14146 & n23651 ;
  assign n14153 = n14145 | n14152 ;
  assign n14154 = x82 & n14153 ;
  assign n14155 = x82 | n14153 ;
  assign n14156 = n13648 & n23456 ;
  assign n14157 = n137 & n14156 ;
  assign n14158 = n13654 & n14157 ;
  assign n14159 = n13654 | n14157 ;
  assign n23652 = ~n14158 ;
  assign n14160 = n23652 & n14159 ;
  assign n23653 = ~n14160 ;
  assign n14161 = n14155 & n23653 ;
  assign n14162 = n14154 | n14161 ;
  assign n14163 = x83 & n14162 ;
  assign n14164 = x83 | n14162 ;
  assign n14165 = n13657 & n23460 ;
  assign n14166 = n137 & n14165 ;
  assign n23654 = ~n13663 ;
  assign n14167 = n23654 & n14166 ;
  assign n23655 = ~n14166 ;
  assign n14168 = n13663 & n23655 ;
  assign n14169 = n14167 | n14168 ;
  assign n23656 = ~n14169 ;
  assign n14170 = n14164 & n23656 ;
  assign n14171 = n14163 | n14170 ;
  assign n14172 = x84 & n14171 ;
  assign n14173 = x84 | n14171 ;
  assign n14174 = n13666 & n23464 ;
  assign n14175 = n137 & n14174 ;
  assign n23657 = ~n13672 ;
  assign n14176 = n23657 & n14175 ;
  assign n23658 = ~n14175 ;
  assign n14177 = n13672 & n23658 ;
  assign n14178 = n14176 | n14177 ;
  assign n23659 = ~n14178 ;
  assign n14179 = n14173 & n23659 ;
  assign n14180 = n14172 | n14179 ;
  assign n14181 = x85 & n14180 ;
  assign n14182 = x85 | n14180 ;
  assign n14183 = n13675 & n23468 ;
  assign n14184 = n137 & n14183 ;
  assign n23660 = ~n13681 ;
  assign n14185 = n23660 & n14184 ;
  assign n23661 = ~n14184 ;
  assign n14186 = n13681 & n23661 ;
  assign n14187 = n14185 | n14186 ;
  assign n23662 = ~n14187 ;
  assign n14188 = n14182 & n23662 ;
  assign n14189 = n14181 | n14188 ;
  assign n14190 = x86 & n14189 ;
  assign n14191 = x86 | n14189 ;
  assign n14192 = n13684 & n23472 ;
  assign n14193 = n137 & n14192 ;
  assign n23663 = ~n13690 ;
  assign n14194 = n23663 & n14193 ;
  assign n23664 = ~n14193 ;
  assign n14195 = n13690 & n23664 ;
  assign n14196 = n14194 | n14195 ;
  assign n23665 = ~n14196 ;
  assign n14197 = n14191 & n23665 ;
  assign n14198 = n14190 | n14197 ;
  assign n14199 = x87 & n14198 ;
  assign n14200 = x87 | n14198 ;
  assign n14201 = n13693 & n23476 ;
  assign n14202 = n137 & n14201 ;
  assign n23666 = ~n13699 ;
  assign n14203 = n23666 & n14202 ;
  assign n23667 = ~n14202 ;
  assign n14204 = n13699 & n23667 ;
  assign n14205 = n14203 | n14204 ;
  assign n23668 = ~n14205 ;
  assign n14206 = n14200 & n23668 ;
  assign n14207 = n14199 | n14206 ;
  assign n14208 = x88 & n14207 ;
  assign n14209 = x88 | n14207 ;
  assign n14210 = n13702 & n23480 ;
  assign n14211 = n137 & n14210 ;
  assign n23669 = ~n13708 ;
  assign n14212 = n23669 & n14211 ;
  assign n23670 = ~n14211 ;
  assign n14213 = n13708 & n23670 ;
  assign n14214 = n14212 | n14213 ;
  assign n23671 = ~n14214 ;
  assign n14215 = n14209 & n23671 ;
  assign n14216 = n14208 | n14215 ;
  assign n14217 = x89 & n14216 ;
  assign n14218 = x89 | n14216 ;
  assign n14219 = n13711 & n23483 ;
  assign n14220 = n137 & n14219 ;
  assign n14221 = n13717 & n14220 ;
  assign n14222 = n13717 | n14220 ;
  assign n23672 = ~n14221 ;
  assign n14223 = n23672 & n14222 ;
  assign n23673 = ~n14223 ;
  assign n14224 = n14218 & n23673 ;
  assign n14225 = n14217 | n14224 ;
  assign n14226 = x90 & n14225 ;
  assign n14227 = x90 | n14225 ;
  assign n14228 = n13720 & n23487 ;
  assign n14229 = n137 & n14228 ;
  assign n23674 = ~n13726 ;
  assign n14230 = n23674 & n14229 ;
  assign n23675 = ~n14229 ;
  assign n14231 = n13726 & n23675 ;
  assign n14232 = n14230 | n14231 ;
  assign n23676 = ~n14232 ;
  assign n14233 = n14227 & n23676 ;
  assign n14234 = n14226 | n14233 ;
  assign n14235 = x91 & n14234 ;
  assign n14236 = x91 | n14234 ;
  assign n14237 = n13729 & n23491 ;
  assign n14238 = n137 & n14237 ;
  assign n23677 = ~n13735 ;
  assign n14239 = n23677 & n14238 ;
  assign n23678 = ~n14238 ;
  assign n14240 = n13735 & n23678 ;
  assign n14241 = n14239 | n14240 ;
  assign n23679 = ~n14241 ;
  assign n14242 = n14236 & n23679 ;
  assign n14243 = n14235 | n14242 ;
  assign n14244 = x92 & n14243 ;
  assign n14245 = x92 | n14243 ;
  assign n14246 = n13738 & n23495 ;
  assign n14247 = n137 & n14246 ;
  assign n23680 = ~n13744 ;
  assign n14248 = n23680 & n14247 ;
  assign n23681 = ~n14247 ;
  assign n14249 = n13744 & n23681 ;
  assign n14250 = n14248 | n14249 ;
  assign n23682 = ~n14250 ;
  assign n14251 = n14245 & n23682 ;
  assign n14252 = n14244 | n14251 ;
  assign n14253 = x93 & n14252 ;
  assign n14254 = x93 | n14252 ;
  assign n14255 = n13747 & n23499 ;
  assign n14256 = n137 & n14255 ;
  assign n14257 = n13753 & n14256 ;
  assign n14258 = n13753 | n14256 ;
  assign n23683 = ~n14257 ;
  assign n14259 = n23683 & n14258 ;
  assign n23684 = ~n14259 ;
  assign n14260 = n14254 & n23684 ;
  assign n14261 = n14253 | n14260 ;
  assign n14262 = x94 & n14261 ;
  assign n14263 = x94 | n14261 ;
  assign n14264 = n13756 & n23503 ;
  assign n14265 = n137 & n14264 ;
  assign n23685 = ~n13762 ;
  assign n14266 = n23685 & n14265 ;
  assign n23686 = ~n14265 ;
  assign n14267 = n13762 & n23686 ;
  assign n14268 = n14266 | n14267 ;
  assign n23687 = ~n14268 ;
  assign n14269 = n14263 & n23687 ;
  assign n14270 = n14262 | n14269 ;
  assign n14271 = x95 & n14270 ;
  assign n14272 = x95 | n14270 ;
  assign n14273 = n13765 & n23506 ;
  assign n14274 = n137 & n14273 ;
  assign n23688 = ~n13771 ;
  assign n14275 = n23688 & n14274 ;
  assign n23689 = ~n14274 ;
  assign n14276 = n13771 & n23689 ;
  assign n14277 = n14275 | n14276 ;
  assign n23690 = ~n14277 ;
  assign n14278 = n14272 & n23690 ;
  assign n14279 = n14271 | n14278 ;
  assign n14280 = x96 & n14279 ;
  assign n14281 = x96 | n14279 ;
  assign n14282 = n13774 & n23510 ;
  assign n14283 = n137 & n14282 ;
  assign n23691 = ~n13780 ;
  assign n14284 = n23691 & n14283 ;
  assign n23692 = ~n14283 ;
  assign n14285 = n13780 & n23692 ;
  assign n14286 = n14284 | n14285 ;
  assign n23693 = ~n14286 ;
  assign n14287 = n14281 & n23693 ;
  assign n14288 = n14280 | n14287 ;
  assign n14289 = x97 & n14288 ;
  assign n14290 = x97 | n14288 ;
  assign n14291 = n13783 & n23514 ;
  assign n14292 = n137 & n14291 ;
  assign n23694 = ~n13789 ;
  assign n14293 = n23694 & n14292 ;
  assign n23695 = ~n14292 ;
  assign n14294 = n13789 & n23695 ;
  assign n14295 = n14293 | n14294 ;
  assign n23696 = ~n14295 ;
  assign n14296 = n14290 & n23696 ;
  assign n14297 = n14289 | n14296 ;
  assign n14298 = x98 & n14297 ;
  assign n14299 = x98 | n14297 ;
  assign n14300 = n13792 & n23517 ;
  assign n14301 = n137 & n14300 ;
  assign n14302 = n13798 & n14301 ;
  assign n14303 = n13798 | n14301 ;
  assign n23697 = ~n14302 ;
  assign n14304 = n23697 & n14303 ;
  assign n23698 = ~n14304 ;
  assign n14305 = n14299 & n23698 ;
  assign n14306 = n14298 | n14305 ;
  assign n14307 = x99 & n14306 ;
  assign n14308 = x99 | n14306 ;
  assign n14309 = n13801 & n23521 ;
  assign n14310 = n137 & n14309 ;
  assign n23699 = ~n13807 ;
  assign n14311 = n23699 & n14310 ;
  assign n23700 = ~n14310 ;
  assign n14312 = n13807 & n23700 ;
  assign n14313 = n14311 | n14312 ;
  assign n23701 = ~n14313 ;
  assign n14314 = n14308 & n23701 ;
  assign n14315 = n14307 | n14314 ;
  assign n14316 = x100 & n14315 ;
  assign n14317 = x100 | n14315 ;
  assign n14318 = n13810 & n23525 ;
  assign n14319 = n137 & n14318 ;
  assign n23702 = ~n13816 ;
  assign n14320 = n23702 & n14319 ;
  assign n23703 = ~n14319 ;
  assign n14321 = n13816 & n23703 ;
  assign n14322 = n14320 | n14321 ;
  assign n23704 = ~n14322 ;
  assign n14323 = n14317 & n23704 ;
  assign n14324 = n14316 | n14323 ;
  assign n14325 = x101 & n14324 ;
  assign n14326 = x101 | n14324 ;
  assign n14327 = n13819 & n23529 ;
  assign n14328 = n137 & n14327 ;
  assign n23705 = ~n13825 ;
  assign n14329 = n23705 & n14328 ;
  assign n23706 = ~n14328 ;
  assign n14330 = n13825 & n23706 ;
  assign n14331 = n14329 | n14330 ;
  assign n23707 = ~n14331 ;
  assign n14332 = n14326 & n23707 ;
  assign n14333 = n14325 | n14332 ;
  assign n14334 = x102 & n14333 ;
  assign n14335 = x102 | n14333 ;
  assign n14336 = n13828 & n23533 ;
  assign n14337 = n137 & n14336 ;
  assign n23708 = ~n13834 ;
  assign n14338 = n23708 & n14337 ;
  assign n23709 = ~n14337 ;
  assign n14339 = n13834 & n23709 ;
  assign n14340 = n14338 | n14339 ;
  assign n23710 = ~n14340 ;
  assign n14341 = n14335 & n23710 ;
  assign n14342 = n14334 | n14341 ;
  assign n14343 = x103 & n14342 ;
  assign n14344 = x103 | n14342 ;
  assign n14345 = n13837 & n23537 ;
  assign n14346 = n137 & n14345 ;
  assign n23711 = ~n13843 ;
  assign n14347 = n23711 & n14346 ;
  assign n23712 = ~n14346 ;
  assign n14348 = n13843 & n23712 ;
  assign n14349 = n14347 | n14348 ;
  assign n23713 = ~n14349 ;
  assign n14350 = n14344 & n23713 ;
  assign n14351 = n14343 | n14350 ;
  assign n14352 = x104 & n14351 ;
  assign n14353 = x104 | n14351 ;
  assign n14354 = n13846 & n23540 ;
  assign n14355 = n137 & n14354 ;
  assign n23714 = ~n13852 ;
  assign n14356 = n23714 & n14355 ;
  assign n23715 = ~n14355 ;
  assign n14357 = n13852 & n23715 ;
  assign n14358 = n14356 | n14357 ;
  assign n23716 = ~n14358 ;
  assign n14359 = n14353 & n23716 ;
  assign n14360 = n14352 | n14359 ;
  assign n14361 = x105 & n14360 ;
  assign n14362 = x105 | n14360 ;
  assign n14363 = n13855 & n23544 ;
  assign n14364 = n137 & n14363 ;
  assign n23717 = ~n13861 ;
  assign n14365 = n23717 & n14364 ;
  assign n23718 = ~n14364 ;
  assign n14366 = n13861 & n23718 ;
  assign n14367 = n14365 | n14366 ;
  assign n23719 = ~n14367 ;
  assign n14368 = n14362 & n23719 ;
  assign n14369 = n14361 | n14368 ;
  assign n14370 = x106 & n14369 ;
  assign n14371 = x106 | n14369 ;
  assign n14372 = n13864 & n23548 ;
  assign n14373 = n137 & n14372 ;
  assign n23720 = ~n13870 ;
  assign n14374 = n23720 & n14373 ;
  assign n23721 = ~n14373 ;
  assign n14375 = n13870 & n23721 ;
  assign n14376 = n14374 | n14375 ;
  assign n23722 = ~n14376 ;
  assign n14377 = n14371 & n23722 ;
  assign n14378 = n14370 | n14377 ;
  assign n14379 = x107 & n14378 ;
  assign n14380 = x107 | n14378 ;
  assign n14381 = n13873 & n23552 ;
  assign n14382 = n137 & n14381 ;
  assign n23723 = ~n13879 ;
  assign n14383 = n23723 & n14382 ;
  assign n23724 = ~n14382 ;
  assign n14384 = n13879 & n23724 ;
  assign n14385 = n14383 | n14384 ;
  assign n23725 = ~n14385 ;
  assign n14386 = n14380 & n23725 ;
  assign n14387 = n14379 | n14386 ;
  assign n14388 = x108 & n14387 ;
  assign n14389 = x108 | n14387 ;
  assign n14390 = n13882 & n23556 ;
  assign n14391 = n137 & n14390 ;
  assign n23726 = ~n13888 ;
  assign n14392 = n23726 & n14391 ;
  assign n23727 = ~n14391 ;
  assign n14393 = n13888 & n23727 ;
  assign n14394 = n14392 | n14393 ;
  assign n23728 = ~n14394 ;
  assign n14395 = n14389 & n23728 ;
  assign n14396 = n14388 | n14395 ;
  assign n14397 = x109 & n14396 ;
  assign n14398 = x109 | n14396 ;
  assign n14399 = n13891 & n23559 ;
  assign n14400 = n137 & n14399 ;
  assign n14401 = n13897 & n14400 ;
  assign n14402 = n13897 | n14400 ;
  assign n23729 = ~n14401 ;
  assign n14403 = n23729 & n14402 ;
  assign n23730 = ~n14403 ;
  assign n14404 = n14398 & n23730 ;
  assign n14405 = n14397 | n14404 ;
  assign n14406 = x110 & n14405 ;
  assign n14407 = x110 | n14405 ;
  assign n14408 = n13900 & n23562 ;
  assign n14409 = n137 & n14408 ;
  assign n14410 = n13906 & n14409 ;
  assign n14411 = n13906 | n14409 ;
  assign n23731 = ~n14410 ;
  assign n14412 = n23731 & n14411 ;
  assign n23732 = ~n14412 ;
  assign n14413 = n14407 & n23732 ;
  assign n14414 = n14406 | n14413 ;
  assign n14415 = x111 & n14414 ;
  assign n14416 = x111 | n14414 ;
  assign n14417 = n13909 & n23565 ;
  assign n14418 = n137 & n14417 ;
  assign n23733 = ~n13915 ;
  assign n14419 = n23733 & n14418 ;
  assign n23734 = ~n14418 ;
  assign n14420 = n13915 & n23734 ;
  assign n14421 = n14419 | n14420 ;
  assign n23735 = ~n14421 ;
  assign n14422 = n14416 & n23735 ;
  assign n14423 = n14415 | n14422 ;
  assign n14424 = x112 & n14423 ;
  assign n14425 = x112 | n14423 ;
  assign n14426 = n13918 & n23569 ;
  assign n14427 = n137 & n14426 ;
  assign n23736 = ~n13924 ;
  assign n14428 = n23736 & n14427 ;
  assign n23737 = ~n14427 ;
  assign n14429 = n13924 & n23737 ;
  assign n14430 = n14428 | n14429 ;
  assign n23738 = ~n14430 ;
  assign n14431 = n14425 & n23738 ;
  assign n14432 = n14424 | n14431 ;
  assign n14433 = x113 & n14432 ;
  assign n14434 = x113 | n14432 ;
  assign n14435 = n13927 & n23573 ;
  assign n14436 = n137 & n14435 ;
  assign n23739 = ~n13933 ;
  assign n14437 = n23739 & n14436 ;
  assign n23740 = ~n14436 ;
  assign n14438 = n13933 & n23740 ;
  assign n14439 = n14437 | n14438 ;
  assign n23741 = ~n14439 ;
  assign n14440 = n14434 & n23741 ;
  assign n14441 = n14433 | n14440 ;
  assign n14442 = x114 & n14441 ;
  assign n14443 = x114 | n14441 ;
  assign n14444 = n13936 & n23577 ;
  assign n14445 = n137 & n14444 ;
  assign n23742 = ~n13942 ;
  assign n14446 = n23742 & n14445 ;
  assign n23743 = ~n14445 ;
  assign n14447 = n13942 & n23743 ;
  assign n14448 = n14446 | n14447 ;
  assign n23744 = ~n14448 ;
  assign n14449 = n14443 & n23744 ;
  assign n14450 = n14442 | n14449 ;
  assign n14451 = x115 & n14450 ;
  assign n14452 = x115 | n14450 ;
  assign n14453 = n13945 & n23581 ;
  assign n14454 = n137 & n14453 ;
  assign n23745 = ~n13951 ;
  assign n14455 = n23745 & n14454 ;
  assign n23746 = ~n14454 ;
  assign n14456 = n13951 & n23746 ;
  assign n14457 = n14455 | n14456 ;
  assign n23747 = ~n14457 ;
  assign n14458 = n14452 & n23747 ;
  assign n14459 = n14451 | n14458 ;
  assign n14460 = x116 & n14459 ;
  assign n14461 = x116 | n14459 ;
  assign n14462 = n13954 & n23585 ;
  assign n14463 = n137 & n14462 ;
  assign n23748 = ~n13960 ;
  assign n14464 = n23748 & n14463 ;
  assign n23749 = ~n14463 ;
  assign n14465 = n13960 & n23749 ;
  assign n14466 = n14464 | n14465 ;
  assign n23750 = ~n14466 ;
  assign n14467 = n14461 & n23750 ;
  assign n14468 = n14460 | n14467 ;
  assign n14469 = x117 & n14468 ;
  assign n14470 = x117 | n14468 ;
  assign n14471 = n13963 & n23589 ;
  assign n14472 = n137 & n14471 ;
  assign n23751 = ~n13969 ;
  assign n14473 = n23751 & n14472 ;
  assign n23752 = ~n14472 ;
  assign n14474 = n13969 & n23752 ;
  assign n14475 = n14473 | n14474 ;
  assign n23753 = ~n14475 ;
  assign n14476 = n14470 & n23753 ;
  assign n14477 = n14469 | n14476 ;
  assign n14478 = x118 & n14477 ;
  assign n14479 = x118 | n14477 ;
  assign n14480 = n13972 & n23593 ;
  assign n14481 = n137 & n14480 ;
  assign n23754 = ~n13978 ;
  assign n14482 = n23754 & n14481 ;
  assign n23755 = ~n14481 ;
  assign n14483 = n13978 & n23755 ;
  assign n14484 = n14482 | n14483 ;
  assign n23756 = ~n14484 ;
  assign n14485 = n14479 & n23756 ;
  assign n14486 = n14478 | n14485 ;
  assign n14488 = x119 & n14486 ;
  assign n23757 = ~n14488 ;
  assign n14489 = n14000 & n23757 ;
  assign n14487 = x119 | n14486 ;
  assign n14490 = x119 & n13984 ;
  assign n14003 = x119 | n13984 ;
  assign n23758 = ~n18298 ;
  assign n14491 = n23758 & n14003 ;
  assign n23759 = ~n14490 ;
  assign n14492 = n23759 & n14491 ;
  assign n23760 = ~n14492 ;
  assign n14493 = n13989 & n23760 ;
  assign n23761 = ~x120 ;
  assign n14494 = n23761 & n14493 ;
  assign n23762 = ~n14494 ;
  assign n14495 = n14487 & n23762 ;
  assign n23763 = ~n14489 ;
  assign n14496 = n23763 & n14495 ;
  assign n14497 = n18293 | n14496 ;
  assign n23764 = ~n14493 ;
  assign n14498 = x120 & n23764 ;
  assign n14499 = n14497 | n14498 ;
  assign n136 = ~n14499 ;
  assign n14500 = x64 & n136 ;
  assign n14501 = x7 & n14500 ;
  assign n14502 = x7 | n14500 ;
  assign n23766 = ~n14501 ;
  assign n14503 = n23766 & n14502 ;
  assign n23767 = ~n5500 ;
  assign n14504 = n23767 & n14503 ;
  assign n23768 = ~n14504 ;
  assign n14505 = n5501 & n23768 ;
  assign n14506 = x66 | n14505 ;
  assign n14507 = x66 & n14505 ;
  assign n14508 = n14002 & n136 ;
  assign n14509 = n23608 & n14508 ;
  assign n14510 = n14006 | n14509 ;
  assign n14511 = n14008 & n14508 ;
  assign n23769 = ~n14511 ;
  assign n14512 = n14510 & n23769 ;
  assign n23770 = ~n14507 ;
  assign n14513 = n23770 & n14512 ;
  assign n23771 = ~n14513 ;
  assign n14514 = n14506 & n23771 ;
  assign n14515 = x67 | n14514 ;
  assign n14516 = x67 & n14514 ;
  assign n23772 = ~n14010 ;
  assign n14517 = n23772 & n14016 ;
  assign n14518 = n136 & n14517 ;
  assign n14519 = n14015 & n14518 ;
  assign n14520 = n14015 | n14518 ;
  assign n23773 = ~n14519 ;
  assign n14521 = n23773 & n14520 ;
  assign n23774 = ~n14516 ;
  assign n14522 = n23774 & n14521 ;
  assign n23775 = ~n14522 ;
  assign n14523 = n14515 & n23775 ;
  assign n14524 = x68 | n14523 ;
  assign n14525 = x68 & n14523 ;
  assign n23776 = ~n14019 ;
  assign n14526 = n23776 & n14020 ;
  assign n14527 = n136 & n14526 ;
  assign n14528 = n14025 & n14527 ;
  assign n14529 = n14025 | n14527 ;
  assign n23777 = ~n14528 ;
  assign n14530 = n23777 & n14529 ;
  assign n23778 = ~n14525 ;
  assign n14531 = n23778 & n14530 ;
  assign n23779 = ~n14531 ;
  assign n14532 = n14524 & n23779 ;
  assign n14533 = x69 | n14532 ;
  assign n14534 = x69 & n14532 ;
  assign n23780 = ~n14028 ;
  assign n14535 = n23780 & n14029 ;
  assign n14536 = n136 & n14535 ;
  assign n14537 = n23617 & n14536 ;
  assign n23781 = ~n14536 ;
  assign n14538 = n14034 & n23781 ;
  assign n14539 = n14537 | n14538 ;
  assign n23782 = ~n14534 ;
  assign n14540 = n23782 & n14539 ;
  assign n23783 = ~n14540 ;
  assign n14541 = n14533 & n23783 ;
  assign n14542 = x70 | n14541 ;
  assign n14543 = x70 & n14541 ;
  assign n23784 = ~n14037 ;
  assign n14544 = n23784 & n14038 ;
  assign n14545 = n136 & n14544 ;
  assign n14546 = n14043 & n14545 ;
  assign n14547 = n14043 | n14545 ;
  assign n23785 = ~n14546 ;
  assign n14548 = n23785 & n14547 ;
  assign n23786 = ~n14543 ;
  assign n14549 = n23786 & n14548 ;
  assign n23787 = ~n14549 ;
  assign n14550 = n14542 & n23787 ;
  assign n14551 = x71 | n14550 ;
  assign n14552 = x71 & n14550 ;
  assign n23788 = ~n14046 ;
  assign n14553 = n23788 & n14047 ;
  assign n14554 = n136 & n14553 ;
  assign n14555 = n14052 & n14554 ;
  assign n14556 = n14052 | n14554 ;
  assign n23789 = ~n14555 ;
  assign n14557 = n23789 & n14556 ;
  assign n23790 = ~n14552 ;
  assign n14558 = n23790 & n14557 ;
  assign n23791 = ~n14558 ;
  assign n14559 = n14551 & n23791 ;
  assign n14560 = x72 | n14559 ;
  assign n14561 = x72 & n14559 ;
  assign n23792 = ~n14055 ;
  assign n14562 = n23792 & n14056 ;
  assign n14563 = n136 & n14562 ;
  assign n14564 = n14061 & n14563 ;
  assign n14565 = n14061 | n14563 ;
  assign n23793 = ~n14564 ;
  assign n14566 = n23793 & n14565 ;
  assign n23794 = ~n14561 ;
  assign n14567 = n23794 & n14566 ;
  assign n23795 = ~n14567 ;
  assign n14568 = n14560 & n23795 ;
  assign n14569 = x73 | n14568 ;
  assign n14570 = x73 & n14568 ;
  assign n23796 = ~n14064 ;
  assign n14571 = n23796 & n14065 ;
  assign n14572 = n136 & n14571 ;
  assign n14573 = n23628 & n14572 ;
  assign n23797 = ~n14572 ;
  assign n14574 = n14070 & n23797 ;
  assign n14575 = n14573 | n14574 ;
  assign n23798 = ~n14570 ;
  assign n14576 = n23798 & n14575 ;
  assign n23799 = ~n14576 ;
  assign n14577 = n14569 & n23799 ;
  assign n14578 = x74 | n14577 ;
  assign n14579 = x74 & n14577 ;
  assign n23800 = ~n14073 ;
  assign n14580 = n23800 & n14074 ;
  assign n14581 = n136 & n14580 ;
  assign n14582 = n14079 & n14581 ;
  assign n14583 = n14079 | n14581 ;
  assign n23801 = ~n14582 ;
  assign n14584 = n23801 & n14583 ;
  assign n23802 = ~n14579 ;
  assign n14585 = n23802 & n14584 ;
  assign n23803 = ~n14585 ;
  assign n14586 = n14578 & n23803 ;
  assign n14587 = x75 | n14586 ;
  assign n14588 = x75 & n14586 ;
  assign n23804 = ~n14082 ;
  assign n14589 = n23804 & n14083 ;
  assign n14590 = n136 & n14589 ;
  assign n14591 = n14088 & n14590 ;
  assign n14592 = n14088 | n14590 ;
  assign n23805 = ~n14591 ;
  assign n14593 = n23805 & n14592 ;
  assign n23806 = ~n14588 ;
  assign n14594 = n23806 & n14593 ;
  assign n23807 = ~n14594 ;
  assign n14595 = n14587 & n23807 ;
  assign n14596 = x76 | n14595 ;
  assign n14597 = x76 & n14595 ;
  assign n23808 = ~n14091 ;
  assign n14598 = n23808 & n14092 ;
  assign n14599 = n136 & n14598 ;
  assign n14600 = n14097 & n14599 ;
  assign n14601 = n14097 | n14599 ;
  assign n23809 = ~n14600 ;
  assign n14602 = n23809 & n14601 ;
  assign n23810 = ~n14597 ;
  assign n14603 = n23810 & n14602 ;
  assign n23811 = ~n14603 ;
  assign n14604 = n14596 & n23811 ;
  assign n14605 = x77 | n14604 ;
  assign n14606 = x77 & n14604 ;
  assign n23812 = ~n14100 ;
  assign n14607 = n23812 & n14101 ;
  assign n14608 = n136 & n14607 ;
  assign n14609 = n14106 & n14608 ;
  assign n14610 = n14106 | n14608 ;
  assign n23813 = ~n14609 ;
  assign n14611 = n23813 & n14610 ;
  assign n23814 = ~n14606 ;
  assign n14612 = n23814 & n14611 ;
  assign n23815 = ~n14612 ;
  assign n14613 = n14605 & n23815 ;
  assign n14614 = x78 | n14613 ;
  assign n14615 = x78 & n14613 ;
  assign n23816 = ~n14109 ;
  assign n14616 = n23816 & n14110 ;
  assign n14617 = n136 & n14616 ;
  assign n14618 = n14115 & n14617 ;
  assign n14619 = n14115 | n14617 ;
  assign n23817 = ~n14618 ;
  assign n14620 = n23817 & n14619 ;
  assign n23818 = ~n14615 ;
  assign n14621 = n23818 & n14620 ;
  assign n23819 = ~n14621 ;
  assign n14622 = n14614 & n23819 ;
  assign n14623 = x79 | n14622 ;
  assign n14624 = x79 & n14622 ;
  assign n23820 = ~n14118 ;
  assign n14625 = n23820 & n14119 ;
  assign n14626 = n136 & n14625 ;
  assign n14627 = n23643 & n14626 ;
  assign n23821 = ~n14626 ;
  assign n14628 = n14124 & n23821 ;
  assign n14629 = n14627 | n14628 ;
  assign n23822 = ~n14624 ;
  assign n14630 = n23822 & n14629 ;
  assign n23823 = ~n14630 ;
  assign n14631 = n14623 & n23823 ;
  assign n14632 = x80 | n14631 ;
  assign n14633 = x80 & n14631 ;
  assign n23824 = ~n14127 ;
  assign n14634 = n23824 & n14128 ;
  assign n14635 = n136 & n14634 ;
  assign n14636 = n14133 & n14635 ;
  assign n14637 = n14133 | n14635 ;
  assign n23825 = ~n14636 ;
  assign n14638 = n23825 & n14637 ;
  assign n23826 = ~n14633 ;
  assign n14639 = n23826 & n14638 ;
  assign n23827 = ~n14639 ;
  assign n14640 = n14632 & n23827 ;
  assign n14641 = x81 | n14640 ;
  assign n14642 = x81 & n14640 ;
  assign n23828 = ~n14136 ;
  assign n14643 = n23828 & n14137 ;
  assign n14644 = n136 & n14643 ;
  assign n14645 = n23648 & n14644 ;
  assign n23829 = ~n14644 ;
  assign n14646 = n14142 & n23829 ;
  assign n14647 = n14645 | n14646 ;
  assign n23830 = ~n14642 ;
  assign n14648 = n23830 & n14647 ;
  assign n23831 = ~n14648 ;
  assign n14649 = n14641 & n23831 ;
  assign n14650 = x82 | n14649 ;
  assign n14651 = x82 & n14649 ;
  assign n23832 = ~n14145 ;
  assign n14652 = n23832 & n14146 ;
  assign n14653 = n136 & n14652 ;
  assign n14654 = n23651 & n14653 ;
  assign n23833 = ~n14653 ;
  assign n14655 = n14151 & n23833 ;
  assign n14656 = n14654 | n14655 ;
  assign n23834 = ~n14651 ;
  assign n14657 = n23834 & n14656 ;
  assign n23835 = ~n14657 ;
  assign n14658 = n14650 & n23835 ;
  assign n14659 = x83 | n14658 ;
  assign n14660 = x83 & n14658 ;
  assign n23836 = ~n14154 ;
  assign n14661 = n23836 & n14155 ;
  assign n14662 = n136 & n14661 ;
  assign n14663 = n14160 & n14662 ;
  assign n14664 = n14160 | n14662 ;
  assign n23837 = ~n14663 ;
  assign n14665 = n23837 & n14664 ;
  assign n23838 = ~n14660 ;
  assign n14666 = n23838 & n14665 ;
  assign n23839 = ~n14666 ;
  assign n14667 = n14659 & n23839 ;
  assign n14668 = x84 | n14667 ;
  assign n14669 = x84 & n14667 ;
  assign n23840 = ~n14163 ;
  assign n14670 = n23840 & n14164 ;
  assign n14671 = n136 & n14670 ;
  assign n14672 = n14169 & n14671 ;
  assign n14673 = n14169 | n14671 ;
  assign n23841 = ~n14672 ;
  assign n14674 = n23841 & n14673 ;
  assign n23842 = ~n14669 ;
  assign n14675 = n23842 & n14674 ;
  assign n23843 = ~n14675 ;
  assign n14676 = n14668 & n23843 ;
  assign n14677 = x85 | n14676 ;
  assign n14678 = x85 & n14676 ;
  assign n23844 = ~n14172 ;
  assign n14679 = n23844 & n14173 ;
  assign n14680 = n136 & n14679 ;
  assign n14681 = n14178 & n14680 ;
  assign n14682 = n14178 | n14680 ;
  assign n23845 = ~n14681 ;
  assign n14683 = n23845 & n14682 ;
  assign n23846 = ~n14678 ;
  assign n14684 = n23846 & n14683 ;
  assign n23847 = ~n14684 ;
  assign n14685 = n14677 & n23847 ;
  assign n14686 = x86 | n14685 ;
  assign n14687 = x86 & n14685 ;
  assign n23848 = ~n14181 ;
  assign n14688 = n23848 & n14182 ;
  assign n14689 = n136 & n14688 ;
  assign n14690 = n14187 & n14689 ;
  assign n14691 = n14187 | n14689 ;
  assign n23849 = ~n14690 ;
  assign n14692 = n23849 & n14691 ;
  assign n23850 = ~n14687 ;
  assign n14693 = n23850 & n14692 ;
  assign n23851 = ~n14693 ;
  assign n14694 = n14686 & n23851 ;
  assign n14695 = x87 | n14694 ;
  assign n14696 = x87 & n14694 ;
  assign n23852 = ~n14190 ;
  assign n14697 = n23852 & n14191 ;
  assign n14698 = n136 & n14697 ;
  assign n14699 = n14196 & n14698 ;
  assign n14700 = n14196 | n14698 ;
  assign n23853 = ~n14699 ;
  assign n14701 = n23853 & n14700 ;
  assign n23854 = ~n14696 ;
  assign n14702 = n23854 & n14701 ;
  assign n23855 = ~n14702 ;
  assign n14703 = n14695 & n23855 ;
  assign n14704 = x88 | n14703 ;
  assign n14705 = x88 & n14703 ;
  assign n23856 = ~n14199 ;
  assign n14706 = n23856 & n14200 ;
  assign n14707 = n136 & n14706 ;
  assign n14708 = n14205 & n14707 ;
  assign n14709 = n14205 | n14707 ;
  assign n23857 = ~n14708 ;
  assign n14710 = n23857 & n14709 ;
  assign n23858 = ~n14705 ;
  assign n14711 = n23858 & n14710 ;
  assign n23859 = ~n14711 ;
  assign n14712 = n14704 & n23859 ;
  assign n14713 = x89 | n14712 ;
  assign n14714 = x89 & n14712 ;
  assign n23860 = ~n14208 ;
  assign n14715 = n23860 & n14209 ;
  assign n14716 = n136 & n14715 ;
  assign n14717 = n23671 & n14716 ;
  assign n23861 = ~n14716 ;
  assign n14718 = n14214 & n23861 ;
  assign n14719 = n14717 | n14718 ;
  assign n23862 = ~n14714 ;
  assign n14720 = n23862 & n14719 ;
  assign n23863 = ~n14720 ;
  assign n14721 = n14713 & n23863 ;
  assign n14722 = x90 | n14721 ;
  assign n14723 = x90 & n14721 ;
  assign n23864 = ~n14217 ;
  assign n14724 = n23864 & n14218 ;
  assign n14725 = n136 & n14724 ;
  assign n14726 = n14223 & n14725 ;
  assign n14727 = n14223 | n14725 ;
  assign n23865 = ~n14726 ;
  assign n14728 = n23865 & n14727 ;
  assign n23866 = ~n14723 ;
  assign n14729 = n23866 & n14728 ;
  assign n23867 = ~n14729 ;
  assign n14730 = n14722 & n23867 ;
  assign n14731 = x91 | n14730 ;
  assign n14732 = x91 & n14730 ;
  assign n23868 = ~n14226 ;
  assign n14733 = n23868 & n14227 ;
  assign n14734 = n136 & n14733 ;
  assign n14735 = n14232 & n14734 ;
  assign n14736 = n14232 | n14734 ;
  assign n23869 = ~n14735 ;
  assign n14737 = n23869 & n14736 ;
  assign n23870 = ~n14732 ;
  assign n14738 = n23870 & n14737 ;
  assign n23871 = ~n14738 ;
  assign n14739 = n14731 & n23871 ;
  assign n14740 = x92 | n14739 ;
  assign n14741 = x92 & n14739 ;
  assign n23872 = ~n14235 ;
  assign n14742 = n23872 & n14236 ;
  assign n14743 = n136 & n14742 ;
  assign n14744 = n14241 & n14743 ;
  assign n14745 = n14241 | n14743 ;
  assign n23873 = ~n14744 ;
  assign n14746 = n23873 & n14745 ;
  assign n23874 = ~n14741 ;
  assign n14747 = n23874 & n14746 ;
  assign n23875 = ~n14747 ;
  assign n14748 = n14740 & n23875 ;
  assign n14749 = x93 | n14748 ;
  assign n14750 = x93 & n14748 ;
  assign n23876 = ~n14244 ;
  assign n14751 = n23876 & n14245 ;
  assign n14752 = n136 & n14751 ;
  assign n14753 = n14250 & n14752 ;
  assign n14754 = n14250 | n14752 ;
  assign n23877 = ~n14753 ;
  assign n14755 = n23877 & n14754 ;
  assign n23878 = ~n14750 ;
  assign n14756 = n23878 & n14755 ;
  assign n23879 = ~n14756 ;
  assign n14757 = n14749 & n23879 ;
  assign n14758 = x94 | n14757 ;
  assign n14759 = x94 & n14757 ;
  assign n23880 = ~n14253 ;
  assign n14760 = n23880 & n14254 ;
  assign n14761 = n136 & n14760 ;
  assign n14762 = n14259 & n14761 ;
  assign n14763 = n14259 | n14761 ;
  assign n23881 = ~n14762 ;
  assign n14764 = n23881 & n14763 ;
  assign n23882 = ~n14759 ;
  assign n14765 = n23882 & n14764 ;
  assign n23883 = ~n14765 ;
  assign n14766 = n14758 & n23883 ;
  assign n14767 = x95 | n14766 ;
  assign n14768 = x95 & n14766 ;
  assign n23884 = ~n14262 ;
  assign n14769 = n23884 & n14263 ;
  assign n14770 = n136 & n14769 ;
  assign n14771 = n14268 & n14770 ;
  assign n14772 = n14268 | n14770 ;
  assign n23885 = ~n14771 ;
  assign n14773 = n23885 & n14772 ;
  assign n23886 = ~n14768 ;
  assign n14774 = n23886 & n14773 ;
  assign n23887 = ~n14774 ;
  assign n14775 = n14767 & n23887 ;
  assign n14776 = x96 | n14775 ;
  assign n14777 = x96 & n14775 ;
  assign n23888 = ~n14271 ;
  assign n14778 = n23888 & n14272 ;
  assign n14779 = n136 & n14778 ;
  assign n14780 = n23690 & n14779 ;
  assign n23889 = ~n14779 ;
  assign n14781 = n14277 & n23889 ;
  assign n14782 = n14780 | n14781 ;
  assign n23890 = ~n14777 ;
  assign n14783 = n23890 & n14782 ;
  assign n23891 = ~n14783 ;
  assign n14784 = n14776 & n23891 ;
  assign n14785 = x97 | n14784 ;
  assign n14786 = x97 & n14784 ;
  assign n23892 = ~n14280 ;
  assign n14787 = n23892 & n14281 ;
  assign n14788 = n136 & n14787 ;
  assign n14789 = n14286 & n14788 ;
  assign n14790 = n14286 | n14788 ;
  assign n23893 = ~n14789 ;
  assign n14791 = n23893 & n14790 ;
  assign n23894 = ~n14786 ;
  assign n14792 = n23894 & n14791 ;
  assign n23895 = ~n14792 ;
  assign n14793 = n14785 & n23895 ;
  assign n14794 = x98 | n14793 ;
  assign n14795 = x98 & n14793 ;
  assign n23896 = ~n14289 ;
  assign n14796 = n23896 & n14290 ;
  assign n14797 = n136 & n14796 ;
  assign n14798 = n23696 & n14797 ;
  assign n23897 = ~n14797 ;
  assign n14799 = n14295 & n23897 ;
  assign n14800 = n14798 | n14799 ;
  assign n23898 = ~n14795 ;
  assign n14801 = n23898 & n14800 ;
  assign n23899 = ~n14801 ;
  assign n14802 = n14794 & n23899 ;
  assign n14803 = x99 | n14802 ;
  assign n14804 = x99 & n14802 ;
  assign n23900 = ~n14298 ;
  assign n14805 = n23900 & n14299 ;
  assign n14806 = n136 & n14805 ;
  assign n14807 = n14304 & n14806 ;
  assign n14808 = n14304 | n14806 ;
  assign n23901 = ~n14807 ;
  assign n14809 = n23901 & n14808 ;
  assign n23902 = ~n14804 ;
  assign n14810 = n23902 & n14809 ;
  assign n23903 = ~n14810 ;
  assign n14811 = n14803 & n23903 ;
  assign n14812 = x100 | n14811 ;
  assign n14813 = x100 & n14811 ;
  assign n23904 = ~n14307 ;
  assign n14814 = n23904 & n14308 ;
  assign n14815 = n136 & n14814 ;
  assign n14816 = n23701 & n14815 ;
  assign n23905 = ~n14815 ;
  assign n14817 = n14313 & n23905 ;
  assign n14818 = n14816 | n14817 ;
  assign n23906 = ~n14813 ;
  assign n14819 = n23906 & n14818 ;
  assign n23907 = ~n14819 ;
  assign n14820 = n14812 & n23907 ;
  assign n14821 = x101 | n14820 ;
  assign n14822 = x101 & n14820 ;
  assign n23908 = ~n14316 ;
  assign n14823 = n23908 & n14317 ;
  assign n14824 = n136 & n14823 ;
  assign n14825 = n14322 & n14824 ;
  assign n14826 = n14322 | n14824 ;
  assign n23909 = ~n14825 ;
  assign n14827 = n23909 & n14826 ;
  assign n23910 = ~n14822 ;
  assign n14828 = n23910 & n14827 ;
  assign n23911 = ~n14828 ;
  assign n14829 = n14821 & n23911 ;
  assign n14830 = x102 | n14829 ;
  assign n14831 = x102 & n14829 ;
  assign n23912 = ~n14325 ;
  assign n14832 = n23912 & n14326 ;
  assign n14833 = n136 & n14832 ;
  assign n14834 = n23707 & n14833 ;
  assign n23913 = ~n14833 ;
  assign n14835 = n14331 & n23913 ;
  assign n14836 = n14834 | n14835 ;
  assign n23914 = ~n14831 ;
  assign n14837 = n23914 & n14836 ;
  assign n23915 = ~n14837 ;
  assign n14838 = n14830 & n23915 ;
  assign n14839 = x103 | n14838 ;
  assign n14840 = x103 & n14838 ;
  assign n23916 = ~n14334 ;
  assign n14841 = n23916 & n14335 ;
  assign n14842 = n136 & n14841 ;
  assign n14843 = n23710 & n14842 ;
  assign n23917 = ~n14842 ;
  assign n14844 = n14340 & n23917 ;
  assign n14845 = n14843 | n14844 ;
  assign n23918 = ~n14840 ;
  assign n14846 = n23918 & n14845 ;
  assign n23919 = ~n14846 ;
  assign n14847 = n14839 & n23919 ;
  assign n14848 = x104 | n14847 ;
  assign n14849 = x104 & n14847 ;
  assign n23920 = ~n14343 ;
  assign n14850 = n23920 & n14344 ;
  assign n14851 = n136 & n14850 ;
  assign n14852 = n14349 & n14851 ;
  assign n14853 = n14349 | n14851 ;
  assign n23921 = ~n14852 ;
  assign n14854 = n23921 & n14853 ;
  assign n23922 = ~n14849 ;
  assign n14855 = n23922 & n14854 ;
  assign n23923 = ~n14855 ;
  assign n14856 = n14848 & n23923 ;
  assign n14857 = x105 | n14856 ;
  assign n14858 = x105 & n14856 ;
  assign n23924 = ~n14352 ;
  assign n14859 = n23924 & n14353 ;
  assign n14860 = n136 & n14859 ;
  assign n14861 = n23716 & n14860 ;
  assign n23925 = ~n14860 ;
  assign n14862 = n14358 & n23925 ;
  assign n14863 = n14861 | n14862 ;
  assign n23926 = ~n14858 ;
  assign n14864 = n23926 & n14863 ;
  assign n23927 = ~n14864 ;
  assign n14865 = n14857 & n23927 ;
  assign n14866 = x106 | n14865 ;
  assign n14867 = x106 & n14865 ;
  assign n23928 = ~n14361 ;
  assign n14868 = n23928 & n14362 ;
  assign n14869 = n136 & n14868 ;
  assign n14870 = n23719 & n14869 ;
  assign n23929 = ~n14869 ;
  assign n14871 = n14367 & n23929 ;
  assign n14872 = n14870 | n14871 ;
  assign n23930 = ~n14867 ;
  assign n14873 = n23930 & n14872 ;
  assign n23931 = ~n14873 ;
  assign n14874 = n14866 & n23931 ;
  assign n14875 = x107 | n14874 ;
  assign n14876 = x107 & n14874 ;
  assign n23932 = ~n14370 ;
  assign n14877 = n23932 & n14371 ;
  assign n14878 = n136 & n14877 ;
  assign n14879 = n23722 & n14878 ;
  assign n23933 = ~n14878 ;
  assign n14880 = n14376 & n23933 ;
  assign n14881 = n14879 | n14880 ;
  assign n23934 = ~n14876 ;
  assign n14882 = n23934 & n14881 ;
  assign n23935 = ~n14882 ;
  assign n14883 = n14875 & n23935 ;
  assign n14884 = x108 | n14883 ;
  assign n14885 = x108 & n14883 ;
  assign n23936 = ~n14379 ;
  assign n14886 = n23936 & n14380 ;
  assign n14887 = n136 & n14886 ;
  assign n14888 = n14385 & n14887 ;
  assign n14889 = n14385 | n14887 ;
  assign n23937 = ~n14888 ;
  assign n14890 = n23937 & n14889 ;
  assign n23938 = ~n14885 ;
  assign n14891 = n23938 & n14890 ;
  assign n23939 = ~n14891 ;
  assign n14892 = n14884 & n23939 ;
  assign n14893 = x109 | n14892 ;
  assign n14894 = x109 & n14892 ;
  assign n23940 = ~n14388 ;
  assign n14895 = n23940 & n14389 ;
  assign n14896 = n136 & n14895 ;
  assign n14897 = n14394 & n14896 ;
  assign n14898 = n14394 | n14896 ;
  assign n23941 = ~n14897 ;
  assign n14899 = n23941 & n14898 ;
  assign n23942 = ~n14894 ;
  assign n14900 = n23942 & n14899 ;
  assign n23943 = ~n14900 ;
  assign n14901 = n14893 & n23943 ;
  assign n14902 = x110 | n14901 ;
  assign n14903 = x110 & n14901 ;
  assign n23944 = ~n14397 ;
  assign n14904 = n23944 & n14398 ;
  assign n14905 = n136 & n14904 ;
  assign n14906 = n14403 & n14905 ;
  assign n14907 = n14403 | n14905 ;
  assign n23945 = ~n14906 ;
  assign n14908 = n23945 & n14907 ;
  assign n23946 = ~n14903 ;
  assign n14909 = n23946 & n14908 ;
  assign n23947 = ~n14909 ;
  assign n14910 = n14902 & n23947 ;
  assign n14911 = x111 | n14910 ;
  assign n14912 = x111 & n14910 ;
  assign n23948 = ~n14406 ;
  assign n14913 = n23948 & n14407 ;
  assign n14914 = n136 & n14913 ;
  assign n14915 = n14412 & n14914 ;
  assign n14916 = n14412 | n14914 ;
  assign n23949 = ~n14915 ;
  assign n14917 = n23949 & n14916 ;
  assign n23950 = ~n14912 ;
  assign n14918 = n23950 & n14917 ;
  assign n23951 = ~n14918 ;
  assign n14919 = n14911 & n23951 ;
  assign n14920 = x112 | n14919 ;
  assign n14921 = x112 & n14919 ;
  assign n23952 = ~n14415 ;
  assign n14922 = n23952 & n14416 ;
  assign n14923 = n136 & n14922 ;
  assign n14924 = n23735 & n14923 ;
  assign n23953 = ~n14923 ;
  assign n14925 = n14421 & n23953 ;
  assign n14926 = n14924 | n14925 ;
  assign n23954 = ~n14921 ;
  assign n14927 = n23954 & n14926 ;
  assign n23955 = ~n14927 ;
  assign n14928 = n14920 & n23955 ;
  assign n14929 = x113 | n14928 ;
  assign n14930 = x113 & n14928 ;
  assign n23956 = ~n14424 ;
  assign n14931 = n23956 & n14425 ;
  assign n14932 = n136 & n14931 ;
  assign n14933 = n23738 & n14932 ;
  assign n23957 = ~n14932 ;
  assign n14934 = n14430 & n23957 ;
  assign n14935 = n14933 | n14934 ;
  assign n23958 = ~n14930 ;
  assign n14936 = n23958 & n14935 ;
  assign n23959 = ~n14936 ;
  assign n14937 = n14929 & n23959 ;
  assign n14938 = x114 | n14937 ;
  assign n14939 = x114 & n14937 ;
  assign n23960 = ~n14433 ;
  assign n14940 = n23960 & n14434 ;
  assign n14941 = n136 & n14940 ;
  assign n14942 = n23741 & n14941 ;
  assign n23961 = ~n14941 ;
  assign n14943 = n14439 & n23961 ;
  assign n14944 = n14942 | n14943 ;
  assign n23962 = ~n14939 ;
  assign n14945 = n23962 & n14944 ;
  assign n23963 = ~n14945 ;
  assign n14946 = n14938 & n23963 ;
  assign n14947 = x115 | n14946 ;
  assign n14948 = x115 & n14946 ;
  assign n23964 = ~n14442 ;
  assign n14949 = n23964 & n14443 ;
  assign n14950 = n136 & n14949 ;
  assign n14951 = n23744 & n14950 ;
  assign n23965 = ~n14950 ;
  assign n14952 = n14448 & n23965 ;
  assign n14953 = n14951 | n14952 ;
  assign n23966 = ~n14948 ;
  assign n14954 = n23966 & n14953 ;
  assign n23967 = ~n14954 ;
  assign n14955 = n14947 & n23967 ;
  assign n14956 = x116 | n14955 ;
  assign n14957 = x116 & n14955 ;
  assign n23968 = ~n14451 ;
  assign n14958 = n23968 & n14452 ;
  assign n14959 = n136 & n14958 ;
  assign n14960 = n23747 & n14959 ;
  assign n23969 = ~n14959 ;
  assign n14961 = n14457 & n23969 ;
  assign n14962 = n14960 | n14961 ;
  assign n23970 = ~n14957 ;
  assign n14963 = n23970 & n14962 ;
  assign n23971 = ~n14963 ;
  assign n14964 = n14956 & n23971 ;
  assign n14965 = x117 | n14964 ;
  assign n14966 = x117 & n14964 ;
  assign n23972 = ~n14460 ;
  assign n14967 = n23972 & n14461 ;
  assign n14968 = n136 & n14967 ;
  assign n14969 = n14466 & n14968 ;
  assign n14970 = n14466 | n14968 ;
  assign n23973 = ~n14969 ;
  assign n14971 = n23973 & n14970 ;
  assign n23974 = ~n14966 ;
  assign n14972 = n23974 & n14971 ;
  assign n23975 = ~n14972 ;
  assign n14973 = n14965 & n23975 ;
  assign n14974 = x118 | n14973 ;
  assign n14975 = x118 & n14973 ;
  assign n23976 = ~n14469 ;
  assign n14976 = n23976 & n14470 ;
  assign n14977 = n136 & n14976 ;
  assign n14978 = n14475 & n14977 ;
  assign n14979 = n14475 | n14977 ;
  assign n23977 = ~n14978 ;
  assign n14980 = n23977 & n14979 ;
  assign n23978 = ~n14975 ;
  assign n14981 = n23978 & n14980 ;
  assign n23979 = ~n14981 ;
  assign n14982 = n14974 & n23979 ;
  assign n14983 = x119 | n14982 ;
  assign n14984 = x119 & n14982 ;
  assign n23980 = ~n14478 ;
  assign n14985 = n23980 & n14479 ;
  assign n14986 = n136 & n14985 ;
  assign n14987 = n23756 & n14986 ;
  assign n23981 = ~n14986 ;
  assign n14988 = n14484 & n23981 ;
  assign n14989 = n14987 | n14988 ;
  assign n23982 = ~n14984 ;
  assign n14990 = n23982 & n14989 ;
  assign n23983 = ~n14990 ;
  assign n14991 = n14983 & n23983 ;
  assign n14992 = x120 | n14991 ;
  assign n14993 = n14487 & n136 ;
  assign n14994 = n23757 & n14993 ;
  assign n14995 = n14000 | n14994 ;
  assign n14996 = n14489 & n14993 ;
  assign n23984 = ~n14996 ;
  assign n14997 = n14995 & n23984 ;
  assign n14998 = x120 & n14991 ;
  assign n23985 = ~n14998 ;
  assign n14999 = n14997 & n23985 ;
  assign n23986 = ~n14999 ;
  assign n15000 = n14992 & n23986 ;
  assign n15001 = x121 & n15000 ;
  assign n15002 = x121 | n15000 ;
  assign n23987 = ~n15001 ;
  assign n15003 = n23987 & n15002 ;
  assign n15004 = n14493 & n14497 ;
  assign n15005 = n21884 | n15004 ;
  assign n23988 = ~n18288 ;
  assign n15008 = n23988 & n15005 ;
  assign n23989 = ~n15003 ;
  assign n15009 = n23989 & n15008 ;
  assign n23990 = ~n15005 ;
  assign n15006 = n15002 & n23990 ;
  assign n15010 = n18288 | n15001 ;
  assign n15011 = n15006 | n15010 ;
  assign n15012 = n14992 & n23985 ;
  assign n135 = ~n15011 ;
  assign n15013 = n135 & n15012 ;
  assign n15014 = n14997 & n15013 ;
  assign n15015 = n14997 | n15013 ;
  assign n23992 = ~n15014 ;
  assign n15016 = n23992 & n15015 ;
  assign n23993 = ~x5 ;
  assign n15017 = n23993 & x64 ;
  assign n15019 = x65 | n15017 ;
  assign n15018 = x65 & n15017 ;
  assign n15020 = x64 & n135 ;
  assign n15021 = x6 & n15020 ;
  assign n15022 = x6 | n15020 ;
  assign n23994 = ~n15021 ;
  assign n15023 = n23994 & n15022 ;
  assign n23995 = ~n15018 ;
  assign n15024 = n23995 & n15023 ;
  assign n23996 = ~n15024 ;
  assign n15025 = n15019 & n23996 ;
  assign n15026 = x66 | n15025 ;
  assign n15027 = x66 & n15025 ;
  assign n15028 = n23767 & n5501 ;
  assign n15029 = n135 & n15028 ;
  assign n15030 = n14503 & n15029 ;
  assign n15031 = n14503 | n15029 ;
  assign n23997 = ~n15030 ;
  assign n15032 = n23997 & n15031 ;
  assign n23998 = ~n15027 ;
  assign n15033 = n23998 & n15032 ;
  assign n23999 = ~n15033 ;
  assign n15034 = n15026 & n23999 ;
  assign n15035 = x67 | n15034 ;
  assign n15036 = x67 & n15034 ;
  assign n15037 = n14506 & n23770 ;
  assign n15038 = n135 & n15037 ;
  assign n24000 = ~n14512 ;
  assign n15039 = n24000 & n15038 ;
  assign n24001 = ~n15038 ;
  assign n15040 = n14512 & n24001 ;
  assign n15041 = n15039 | n15040 ;
  assign n24002 = ~n15036 ;
  assign n15042 = n24002 & n15041 ;
  assign n24003 = ~n15042 ;
  assign n15043 = n15035 & n24003 ;
  assign n15044 = x68 | n15043 ;
  assign n15045 = x68 & n15043 ;
  assign n15046 = n14515 & n23774 ;
  assign n15047 = n135 & n15046 ;
  assign n24004 = ~n14521 ;
  assign n15048 = n24004 & n15047 ;
  assign n24005 = ~n15047 ;
  assign n15049 = n14521 & n24005 ;
  assign n15050 = n15048 | n15049 ;
  assign n24006 = ~n15045 ;
  assign n15051 = n24006 & n15050 ;
  assign n24007 = ~n15051 ;
  assign n15052 = n15044 & n24007 ;
  assign n15053 = x69 | n15052 ;
  assign n15054 = x69 & n15052 ;
  assign n15055 = n14524 & n23778 ;
  assign n15056 = n135 & n15055 ;
  assign n24008 = ~n14530 ;
  assign n15057 = n24008 & n15056 ;
  assign n24009 = ~n15056 ;
  assign n15058 = n14530 & n24009 ;
  assign n15059 = n15057 | n15058 ;
  assign n24010 = ~n15054 ;
  assign n15060 = n24010 & n15059 ;
  assign n24011 = ~n15060 ;
  assign n15061 = n15053 & n24011 ;
  assign n15062 = x70 | n15061 ;
  assign n15063 = x70 & n15061 ;
  assign n15064 = n14533 & n23782 ;
  assign n15065 = n135 & n15064 ;
  assign n24012 = ~n14539 ;
  assign n15066 = n24012 & n15065 ;
  assign n24013 = ~n15065 ;
  assign n15067 = n14539 & n24013 ;
  assign n15068 = n15066 | n15067 ;
  assign n24014 = ~n15063 ;
  assign n15069 = n24014 & n15068 ;
  assign n24015 = ~n15069 ;
  assign n15070 = n15062 & n24015 ;
  assign n15071 = x71 | n15070 ;
  assign n15072 = x71 & n15070 ;
  assign n15073 = n14542 & n23786 ;
  assign n15074 = n135 & n15073 ;
  assign n15075 = n14548 & n15074 ;
  assign n15076 = n14548 | n15074 ;
  assign n24016 = ~n15075 ;
  assign n15077 = n24016 & n15076 ;
  assign n24017 = ~n15072 ;
  assign n15078 = n24017 & n15077 ;
  assign n24018 = ~n15078 ;
  assign n15079 = n15071 & n24018 ;
  assign n15080 = x72 | n15079 ;
  assign n15081 = x72 & n15079 ;
  assign n15082 = n14551 & n23790 ;
  assign n15083 = n135 & n15082 ;
  assign n24019 = ~n14557 ;
  assign n15084 = n24019 & n15083 ;
  assign n24020 = ~n15083 ;
  assign n15085 = n14557 & n24020 ;
  assign n15086 = n15084 | n15085 ;
  assign n24021 = ~n15081 ;
  assign n15087 = n24021 & n15086 ;
  assign n24022 = ~n15087 ;
  assign n15088 = n15080 & n24022 ;
  assign n15089 = x73 | n15088 ;
  assign n15090 = x73 & n15088 ;
  assign n15091 = n14560 & n23794 ;
  assign n15092 = n135 & n15091 ;
  assign n15093 = n14566 & n15092 ;
  assign n15094 = n14566 | n15092 ;
  assign n24023 = ~n15093 ;
  assign n15095 = n24023 & n15094 ;
  assign n24024 = ~n15090 ;
  assign n15096 = n24024 & n15095 ;
  assign n24025 = ~n15096 ;
  assign n15097 = n15089 & n24025 ;
  assign n15098 = x74 | n15097 ;
  assign n15099 = x74 & n15097 ;
  assign n15100 = n14569 & n23798 ;
  assign n15101 = n135 & n15100 ;
  assign n24026 = ~n14575 ;
  assign n15102 = n24026 & n15101 ;
  assign n24027 = ~n15101 ;
  assign n15103 = n14575 & n24027 ;
  assign n15104 = n15102 | n15103 ;
  assign n24028 = ~n15099 ;
  assign n15105 = n24028 & n15104 ;
  assign n24029 = ~n15105 ;
  assign n15106 = n15098 & n24029 ;
  assign n15107 = x75 | n15106 ;
  assign n15108 = x75 & n15106 ;
  assign n15109 = n14578 & n23802 ;
  assign n15110 = n135 & n15109 ;
  assign n24030 = ~n14584 ;
  assign n15111 = n24030 & n15110 ;
  assign n24031 = ~n15110 ;
  assign n15112 = n14584 & n24031 ;
  assign n15113 = n15111 | n15112 ;
  assign n24032 = ~n15108 ;
  assign n15114 = n24032 & n15113 ;
  assign n24033 = ~n15114 ;
  assign n15115 = n15107 & n24033 ;
  assign n15116 = x76 | n15115 ;
  assign n15117 = x76 & n15115 ;
  assign n15118 = n14587 & n23806 ;
  assign n15119 = n135 & n15118 ;
  assign n24034 = ~n14593 ;
  assign n15120 = n24034 & n15119 ;
  assign n24035 = ~n15119 ;
  assign n15121 = n14593 & n24035 ;
  assign n15122 = n15120 | n15121 ;
  assign n24036 = ~n15117 ;
  assign n15123 = n24036 & n15122 ;
  assign n24037 = ~n15123 ;
  assign n15124 = n15116 & n24037 ;
  assign n15125 = x77 | n15124 ;
  assign n15126 = x77 & n15124 ;
  assign n15127 = n14596 & n23810 ;
  assign n15128 = n135 & n15127 ;
  assign n15129 = n14602 & n15128 ;
  assign n15130 = n14602 | n15128 ;
  assign n24038 = ~n15129 ;
  assign n15131 = n24038 & n15130 ;
  assign n24039 = ~n15126 ;
  assign n15132 = n24039 & n15131 ;
  assign n24040 = ~n15132 ;
  assign n15133 = n15125 & n24040 ;
  assign n15134 = x78 | n15133 ;
  assign n15135 = x78 & n15133 ;
  assign n15136 = n14605 & n23814 ;
  assign n15137 = n135 & n15136 ;
  assign n15138 = n14611 & n15137 ;
  assign n15139 = n14611 | n15137 ;
  assign n24041 = ~n15138 ;
  assign n15140 = n24041 & n15139 ;
  assign n24042 = ~n15135 ;
  assign n15141 = n24042 & n15140 ;
  assign n24043 = ~n15141 ;
  assign n15142 = n15134 & n24043 ;
  assign n15143 = x79 | n15142 ;
  assign n15144 = x79 & n15142 ;
  assign n15145 = n14614 & n23818 ;
  assign n15146 = n135 & n15145 ;
  assign n24044 = ~n14620 ;
  assign n15147 = n24044 & n15146 ;
  assign n24045 = ~n15146 ;
  assign n15148 = n14620 & n24045 ;
  assign n15149 = n15147 | n15148 ;
  assign n24046 = ~n15144 ;
  assign n15150 = n24046 & n15149 ;
  assign n24047 = ~n15150 ;
  assign n15151 = n15143 & n24047 ;
  assign n15152 = x80 | n15151 ;
  assign n15153 = x80 & n15151 ;
  assign n15154 = n14623 & n23822 ;
  assign n15155 = n135 & n15154 ;
  assign n24048 = ~n14629 ;
  assign n15156 = n24048 & n15155 ;
  assign n24049 = ~n15155 ;
  assign n15157 = n14629 & n24049 ;
  assign n15158 = n15156 | n15157 ;
  assign n24050 = ~n15153 ;
  assign n15159 = n24050 & n15158 ;
  assign n24051 = ~n15159 ;
  assign n15160 = n15152 & n24051 ;
  assign n15161 = x81 | n15160 ;
  assign n15162 = x81 & n15160 ;
  assign n15163 = n14632 & n23826 ;
  assign n15164 = n135 & n15163 ;
  assign n24052 = ~n14638 ;
  assign n15165 = n24052 & n15164 ;
  assign n24053 = ~n15164 ;
  assign n15166 = n14638 & n24053 ;
  assign n15167 = n15165 | n15166 ;
  assign n24054 = ~n15162 ;
  assign n15168 = n24054 & n15167 ;
  assign n24055 = ~n15168 ;
  assign n15169 = n15161 & n24055 ;
  assign n15170 = x82 | n15169 ;
  assign n15171 = x82 & n15169 ;
  assign n15172 = n14641 & n23830 ;
  assign n15173 = n135 & n15172 ;
  assign n24056 = ~n14647 ;
  assign n15174 = n24056 & n15173 ;
  assign n24057 = ~n15173 ;
  assign n15175 = n14647 & n24057 ;
  assign n15176 = n15174 | n15175 ;
  assign n24058 = ~n15171 ;
  assign n15177 = n24058 & n15176 ;
  assign n24059 = ~n15177 ;
  assign n15178 = n15170 & n24059 ;
  assign n15179 = x83 | n15178 ;
  assign n15180 = x83 & n15178 ;
  assign n15181 = n14650 & n23834 ;
  assign n15182 = n135 & n15181 ;
  assign n24060 = ~n14656 ;
  assign n15183 = n24060 & n15182 ;
  assign n24061 = ~n15182 ;
  assign n15184 = n14656 & n24061 ;
  assign n15185 = n15183 | n15184 ;
  assign n24062 = ~n15180 ;
  assign n15186 = n24062 & n15185 ;
  assign n24063 = ~n15186 ;
  assign n15187 = n15179 & n24063 ;
  assign n15188 = x84 | n15187 ;
  assign n15189 = x84 & n15187 ;
  assign n15190 = n14659 & n23838 ;
  assign n15191 = n135 & n15190 ;
  assign n24064 = ~n14665 ;
  assign n15192 = n24064 & n15191 ;
  assign n24065 = ~n15191 ;
  assign n15193 = n14665 & n24065 ;
  assign n15194 = n15192 | n15193 ;
  assign n24066 = ~n15189 ;
  assign n15195 = n24066 & n15194 ;
  assign n24067 = ~n15195 ;
  assign n15196 = n15188 & n24067 ;
  assign n15197 = x85 | n15196 ;
  assign n15198 = x85 & n15196 ;
  assign n15199 = n14668 & n23842 ;
  assign n15200 = n135 & n15199 ;
  assign n15201 = n14674 & n15200 ;
  assign n15202 = n14674 | n15200 ;
  assign n24068 = ~n15201 ;
  assign n15203 = n24068 & n15202 ;
  assign n24069 = ~n15198 ;
  assign n15204 = n24069 & n15203 ;
  assign n24070 = ~n15204 ;
  assign n15205 = n15197 & n24070 ;
  assign n15206 = x86 | n15205 ;
  assign n15207 = x86 & n15205 ;
  assign n15208 = n14677 & n23846 ;
  assign n15209 = n135 & n15208 ;
  assign n15210 = n14683 & n15209 ;
  assign n15211 = n14683 | n15209 ;
  assign n24071 = ~n15210 ;
  assign n15212 = n24071 & n15211 ;
  assign n24072 = ~n15207 ;
  assign n15213 = n24072 & n15212 ;
  assign n24073 = ~n15213 ;
  assign n15214 = n15206 & n24073 ;
  assign n15215 = x87 | n15214 ;
  assign n15216 = x87 & n15214 ;
  assign n15217 = n14686 & n23850 ;
  assign n15218 = n135 & n15217 ;
  assign n15219 = n14692 & n15218 ;
  assign n15220 = n14692 | n15218 ;
  assign n24074 = ~n15219 ;
  assign n15221 = n24074 & n15220 ;
  assign n24075 = ~n15216 ;
  assign n15222 = n24075 & n15221 ;
  assign n24076 = ~n15222 ;
  assign n15223 = n15215 & n24076 ;
  assign n15224 = x88 | n15223 ;
  assign n15225 = x88 & n15223 ;
  assign n15226 = n14695 & n23854 ;
  assign n15227 = n135 & n15226 ;
  assign n15228 = n14701 & n15227 ;
  assign n15229 = n14701 | n15227 ;
  assign n24077 = ~n15228 ;
  assign n15230 = n24077 & n15229 ;
  assign n24078 = ~n15225 ;
  assign n15231 = n24078 & n15230 ;
  assign n24079 = ~n15231 ;
  assign n15232 = n15224 & n24079 ;
  assign n15233 = x89 | n15232 ;
  assign n15234 = x89 & n15232 ;
  assign n15235 = n14704 & n23858 ;
  assign n15236 = n135 & n15235 ;
  assign n15237 = n14710 & n15236 ;
  assign n15238 = n14710 | n15236 ;
  assign n24080 = ~n15237 ;
  assign n15239 = n24080 & n15238 ;
  assign n24081 = ~n15234 ;
  assign n15240 = n24081 & n15239 ;
  assign n24082 = ~n15240 ;
  assign n15241 = n15233 & n24082 ;
  assign n15242 = x90 | n15241 ;
  assign n15243 = x90 & n15241 ;
  assign n15244 = n14713 & n23862 ;
  assign n15245 = n135 & n15244 ;
  assign n24083 = ~n14719 ;
  assign n15246 = n24083 & n15245 ;
  assign n24084 = ~n15245 ;
  assign n15247 = n14719 & n24084 ;
  assign n15248 = n15246 | n15247 ;
  assign n24085 = ~n15243 ;
  assign n15249 = n24085 & n15248 ;
  assign n24086 = ~n15249 ;
  assign n15250 = n15242 & n24086 ;
  assign n15251 = x91 | n15250 ;
  assign n15252 = x91 & n15250 ;
  assign n15253 = n14722 & n23866 ;
  assign n15254 = n135 & n15253 ;
  assign n24087 = ~n14728 ;
  assign n15255 = n24087 & n15254 ;
  assign n24088 = ~n15254 ;
  assign n15256 = n14728 & n24088 ;
  assign n15257 = n15255 | n15256 ;
  assign n24089 = ~n15252 ;
  assign n15258 = n24089 & n15257 ;
  assign n24090 = ~n15258 ;
  assign n15259 = n15251 & n24090 ;
  assign n15260 = x92 | n15259 ;
  assign n15261 = x92 & n15259 ;
  assign n15262 = n14731 & n23870 ;
  assign n15263 = n135 & n15262 ;
  assign n15264 = n14737 & n15263 ;
  assign n15265 = n14737 | n15263 ;
  assign n24091 = ~n15264 ;
  assign n15266 = n24091 & n15265 ;
  assign n24092 = ~n15261 ;
  assign n15267 = n24092 & n15266 ;
  assign n24093 = ~n15267 ;
  assign n15268 = n15260 & n24093 ;
  assign n15269 = x93 | n15268 ;
  assign n15270 = x93 & n15268 ;
  assign n15271 = n14740 & n23874 ;
  assign n15272 = n135 & n15271 ;
  assign n15273 = n14746 & n15272 ;
  assign n15274 = n14746 | n15272 ;
  assign n24094 = ~n15273 ;
  assign n15275 = n24094 & n15274 ;
  assign n24095 = ~n15270 ;
  assign n15276 = n24095 & n15275 ;
  assign n24096 = ~n15276 ;
  assign n15277 = n15269 & n24096 ;
  assign n15278 = x94 | n15277 ;
  assign n15279 = x94 & n15277 ;
  assign n15280 = n14749 & n23878 ;
  assign n15281 = n135 & n15280 ;
  assign n15282 = n14755 & n15281 ;
  assign n15283 = n14755 | n15281 ;
  assign n24097 = ~n15282 ;
  assign n15284 = n24097 & n15283 ;
  assign n24098 = ~n15279 ;
  assign n15285 = n24098 & n15284 ;
  assign n24099 = ~n15285 ;
  assign n15286 = n15278 & n24099 ;
  assign n15287 = x95 | n15286 ;
  assign n15288 = x95 & n15286 ;
  assign n15289 = n14758 & n23882 ;
  assign n15290 = n135 & n15289 ;
  assign n24100 = ~n14764 ;
  assign n15291 = n24100 & n15290 ;
  assign n24101 = ~n15290 ;
  assign n15292 = n14764 & n24101 ;
  assign n15293 = n15291 | n15292 ;
  assign n24102 = ~n15288 ;
  assign n15294 = n24102 & n15293 ;
  assign n24103 = ~n15294 ;
  assign n15295 = n15287 & n24103 ;
  assign n15296 = x96 | n15295 ;
  assign n15297 = x96 & n15295 ;
  assign n15298 = n14767 & n23886 ;
  assign n15299 = n135 & n15298 ;
  assign n15300 = n14773 & n15299 ;
  assign n15301 = n14773 | n15299 ;
  assign n24104 = ~n15300 ;
  assign n15302 = n24104 & n15301 ;
  assign n24105 = ~n15297 ;
  assign n15303 = n24105 & n15302 ;
  assign n24106 = ~n15303 ;
  assign n15304 = n15296 & n24106 ;
  assign n15305 = x97 | n15304 ;
  assign n15306 = x97 & n15304 ;
  assign n15307 = n14776 & n23890 ;
  assign n15308 = n135 & n15307 ;
  assign n24107 = ~n14782 ;
  assign n15309 = n24107 & n15308 ;
  assign n24108 = ~n15308 ;
  assign n15310 = n14782 & n24108 ;
  assign n15311 = n15309 | n15310 ;
  assign n24109 = ~n15306 ;
  assign n15312 = n24109 & n15311 ;
  assign n24110 = ~n15312 ;
  assign n15313 = n15305 & n24110 ;
  assign n15314 = x98 | n15313 ;
  assign n15315 = x98 & n15313 ;
  assign n15316 = n14785 & n23894 ;
  assign n15317 = n135 & n15316 ;
  assign n15318 = n14791 & n15317 ;
  assign n15319 = n14791 | n15317 ;
  assign n24111 = ~n15318 ;
  assign n15320 = n24111 & n15319 ;
  assign n24112 = ~n15315 ;
  assign n15321 = n24112 & n15320 ;
  assign n24113 = ~n15321 ;
  assign n15322 = n15314 & n24113 ;
  assign n15323 = x99 | n15322 ;
  assign n15324 = x99 & n15322 ;
  assign n15325 = n14794 & n23898 ;
  assign n15326 = n135 & n15325 ;
  assign n24114 = ~n14800 ;
  assign n15327 = n24114 & n15326 ;
  assign n24115 = ~n15326 ;
  assign n15328 = n14800 & n24115 ;
  assign n15329 = n15327 | n15328 ;
  assign n24116 = ~n15324 ;
  assign n15330 = n24116 & n15329 ;
  assign n24117 = ~n15330 ;
  assign n15331 = n15323 & n24117 ;
  assign n15332 = x100 | n15331 ;
  assign n15333 = x100 & n15331 ;
  assign n15334 = n14803 & n23902 ;
  assign n15335 = n135 & n15334 ;
  assign n24118 = ~n14809 ;
  assign n15336 = n24118 & n15335 ;
  assign n24119 = ~n15335 ;
  assign n15337 = n14809 & n24119 ;
  assign n15338 = n15336 | n15337 ;
  assign n24120 = ~n15333 ;
  assign n15339 = n24120 & n15338 ;
  assign n24121 = ~n15339 ;
  assign n15340 = n15332 & n24121 ;
  assign n15341 = x101 | n15340 ;
  assign n15342 = x101 & n15340 ;
  assign n15343 = n14812 & n23906 ;
  assign n15344 = n135 & n15343 ;
  assign n24122 = ~n14818 ;
  assign n15345 = n24122 & n15344 ;
  assign n24123 = ~n15344 ;
  assign n15346 = n14818 & n24123 ;
  assign n15347 = n15345 | n15346 ;
  assign n24124 = ~n15342 ;
  assign n15348 = n24124 & n15347 ;
  assign n24125 = ~n15348 ;
  assign n15349 = n15341 & n24125 ;
  assign n15350 = x102 | n15349 ;
  assign n15351 = x102 & n15349 ;
  assign n15352 = n14821 & n23910 ;
  assign n15353 = n135 & n15352 ;
  assign n15354 = n14827 & n15353 ;
  assign n15355 = n14827 | n15353 ;
  assign n24126 = ~n15354 ;
  assign n15356 = n24126 & n15355 ;
  assign n24127 = ~n15351 ;
  assign n15357 = n24127 & n15356 ;
  assign n24128 = ~n15357 ;
  assign n15358 = n15350 & n24128 ;
  assign n15359 = x103 | n15358 ;
  assign n15360 = x103 & n15358 ;
  assign n15361 = n14830 & n23914 ;
  assign n15362 = n135 & n15361 ;
  assign n24129 = ~n14836 ;
  assign n15363 = n24129 & n15362 ;
  assign n24130 = ~n15362 ;
  assign n15364 = n14836 & n24130 ;
  assign n15365 = n15363 | n15364 ;
  assign n24131 = ~n15360 ;
  assign n15366 = n24131 & n15365 ;
  assign n24132 = ~n15366 ;
  assign n15367 = n15359 & n24132 ;
  assign n15368 = x104 | n15367 ;
  assign n15369 = x104 & n15367 ;
  assign n15370 = n14839 & n23918 ;
  assign n15371 = n135 & n15370 ;
  assign n24133 = ~n14845 ;
  assign n15372 = n24133 & n15371 ;
  assign n24134 = ~n15371 ;
  assign n15373 = n14845 & n24134 ;
  assign n15374 = n15372 | n15373 ;
  assign n24135 = ~n15369 ;
  assign n15375 = n24135 & n15374 ;
  assign n24136 = ~n15375 ;
  assign n15376 = n15368 & n24136 ;
  assign n15377 = x105 | n15376 ;
  assign n15378 = x105 & n15376 ;
  assign n15379 = n14848 & n23922 ;
  assign n15380 = n135 & n15379 ;
  assign n15381 = n14854 & n15380 ;
  assign n15382 = n14854 | n15380 ;
  assign n24137 = ~n15381 ;
  assign n15383 = n24137 & n15382 ;
  assign n24138 = ~n15378 ;
  assign n15384 = n24138 & n15383 ;
  assign n24139 = ~n15384 ;
  assign n15385 = n15377 & n24139 ;
  assign n15386 = x106 | n15385 ;
  assign n15387 = x106 & n15385 ;
  assign n15388 = n14857 & n23926 ;
  assign n15389 = n135 & n15388 ;
  assign n24140 = ~n14863 ;
  assign n15390 = n24140 & n15389 ;
  assign n24141 = ~n15389 ;
  assign n15391 = n14863 & n24141 ;
  assign n15392 = n15390 | n15391 ;
  assign n24142 = ~n15387 ;
  assign n15393 = n24142 & n15392 ;
  assign n24143 = ~n15393 ;
  assign n15394 = n15386 & n24143 ;
  assign n15395 = x107 | n15394 ;
  assign n15396 = x107 & n15394 ;
  assign n15397 = n14866 & n23930 ;
  assign n15398 = n135 & n15397 ;
  assign n24144 = ~n14872 ;
  assign n15399 = n24144 & n15398 ;
  assign n24145 = ~n15398 ;
  assign n15400 = n14872 & n24145 ;
  assign n15401 = n15399 | n15400 ;
  assign n24146 = ~n15396 ;
  assign n15402 = n24146 & n15401 ;
  assign n24147 = ~n15402 ;
  assign n15403 = n15395 & n24147 ;
  assign n15404 = x108 | n15403 ;
  assign n15405 = x108 & n15403 ;
  assign n15406 = n14875 & n23934 ;
  assign n15407 = n135 & n15406 ;
  assign n24148 = ~n14881 ;
  assign n15408 = n24148 & n15407 ;
  assign n24149 = ~n15407 ;
  assign n15409 = n14881 & n24149 ;
  assign n15410 = n15408 | n15409 ;
  assign n24150 = ~n15405 ;
  assign n15411 = n24150 & n15410 ;
  assign n24151 = ~n15411 ;
  assign n15412 = n15404 & n24151 ;
  assign n15413 = x109 | n15412 ;
  assign n15414 = x109 & n15412 ;
  assign n15415 = n14884 & n23938 ;
  assign n15416 = n135 & n15415 ;
  assign n15417 = n14890 & n15416 ;
  assign n15418 = n14890 | n15416 ;
  assign n24152 = ~n15417 ;
  assign n15419 = n24152 & n15418 ;
  assign n24153 = ~n15414 ;
  assign n15420 = n24153 & n15419 ;
  assign n24154 = ~n15420 ;
  assign n15421 = n15413 & n24154 ;
  assign n15422 = x110 | n15421 ;
  assign n15423 = x110 & n15421 ;
  assign n15424 = n14893 & n23942 ;
  assign n15425 = n135 & n15424 ;
  assign n15426 = n14899 & n15425 ;
  assign n15427 = n14899 | n15425 ;
  assign n24155 = ~n15426 ;
  assign n15428 = n24155 & n15427 ;
  assign n24156 = ~n15423 ;
  assign n15429 = n24156 & n15428 ;
  assign n24157 = ~n15429 ;
  assign n15430 = n15422 & n24157 ;
  assign n15431 = x111 | n15430 ;
  assign n15432 = x111 & n15430 ;
  assign n15433 = n14902 & n23946 ;
  assign n15434 = n135 & n15433 ;
  assign n24158 = ~n14908 ;
  assign n15435 = n24158 & n15434 ;
  assign n24159 = ~n15434 ;
  assign n15436 = n14908 & n24159 ;
  assign n15437 = n15435 | n15436 ;
  assign n24160 = ~n15432 ;
  assign n15438 = n24160 & n15437 ;
  assign n24161 = ~n15438 ;
  assign n15439 = n15431 & n24161 ;
  assign n15440 = x112 | n15439 ;
  assign n15441 = x112 & n15439 ;
  assign n15442 = n14911 & n23950 ;
  assign n15443 = n135 & n15442 ;
  assign n24162 = ~n14917 ;
  assign n15444 = n24162 & n15443 ;
  assign n24163 = ~n15443 ;
  assign n15445 = n14917 & n24163 ;
  assign n15446 = n15444 | n15445 ;
  assign n24164 = ~n15441 ;
  assign n15447 = n24164 & n15446 ;
  assign n24165 = ~n15447 ;
  assign n15448 = n15440 & n24165 ;
  assign n15449 = x113 | n15448 ;
  assign n15450 = x113 & n15448 ;
  assign n15451 = n14920 & n23954 ;
  assign n15452 = n135 & n15451 ;
  assign n24166 = ~n14926 ;
  assign n15453 = n24166 & n15452 ;
  assign n24167 = ~n15452 ;
  assign n15454 = n14926 & n24167 ;
  assign n15455 = n15453 | n15454 ;
  assign n24168 = ~n15450 ;
  assign n15456 = n24168 & n15455 ;
  assign n24169 = ~n15456 ;
  assign n15457 = n15449 & n24169 ;
  assign n15458 = x114 | n15457 ;
  assign n15459 = x114 & n15457 ;
  assign n15460 = n14929 & n23958 ;
  assign n15461 = n135 & n15460 ;
  assign n24170 = ~n14935 ;
  assign n15462 = n24170 & n15461 ;
  assign n24171 = ~n15461 ;
  assign n15463 = n14935 & n24171 ;
  assign n15464 = n15462 | n15463 ;
  assign n24172 = ~n15459 ;
  assign n15465 = n24172 & n15464 ;
  assign n24173 = ~n15465 ;
  assign n15466 = n15458 & n24173 ;
  assign n15467 = x115 | n15466 ;
  assign n15468 = x115 & n15466 ;
  assign n15469 = n14938 & n23962 ;
  assign n15470 = n135 & n15469 ;
  assign n24174 = ~n14944 ;
  assign n15471 = n24174 & n15470 ;
  assign n24175 = ~n15470 ;
  assign n15472 = n14944 & n24175 ;
  assign n15473 = n15471 | n15472 ;
  assign n24176 = ~n15468 ;
  assign n15474 = n24176 & n15473 ;
  assign n24177 = ~n15474 ;
  assign n15475 = n15467 & n24177 ;
  assign n15476 = x116 | n15475 ;
  assign n15477 = x116 & n15475 ;
  assign n15478 = n14947 & n23966 ;
  assign n15479 = n135 & n15478 ;
  assign n24178 = ~n14953 ;
  assign n15480 = n24178 & n15479 ;
  assign n24179 = ~n15479 ;
  assign n15481 = n14953 & n24179 ;
  assign n15482 = n15480 | n15481 ;
  assign n24180 = ~n15477 ;
  assign n15483 = n24180 & n15482 ;
  assign n24181 = ~n15483 ;
  assign n15484 = n15476 & n24181 ;
  assign n15485 = x117 | n15484 ;
  assign n15486 = x117 & n15484 ;
  assign n15487 = n14956 & n23970 ;
  assign n15488 = n135 & n15487 ;
  assign n24182 = ~n14962 ;
  assign n15489 = n24182 & n15488 ;
  assign n24183 = ~n15488 ;
  assign n15490 = n14962 & n24183 ;
  assign n15491 = n15489 | n15490 ;
  assign n24184 = ~n15486 ;
  assign n15492 = n24184 & n15491 ;
  assign n24185 = ~n15492 ;
  assign n15493 = n15485 & n24185 ;
  assign n15494 = x118 | n15493 ;
  assign n15495 = x118 & n15493 ;
  assign n15496 = n14965 & n23974 ;
  assign n15497 = n135 & n15496 ;
  assign n15498 = n14971 & n15497 ;
  assign n15499 = n14971 | n15497 ;
  assign n24186 = ~n15498 ;
  assign n15500 = n24186 & n15499 ;
  assign n24187 = ~n15495 ;
  assign n15501 = n24187 & n15500 ;
  assign n24188 = ~n15501 ;
  assign n15502 = n15494 & n24188 ;
  assign n15503 = x119 | n15502 ;
  assign n15504 = x119 & n15502 ;
  assign n15505 = n14974 & n23978 ;
  assign n15506 = n135 & n15505 ;
  assign n15507 = n14980 & n15506 ;
  assign n15508 = n14980 | n15506 ;
  assign n24189 = ~n15507 ;
  assign n15509 = n24189 & n15508 ;
  assign n24190 = ~n15504 ;
  assign n15510 = n24190 & n15509 ;
  assign n24191 = ~n15510 ;
  assign n15511 = n15503 & n24191 ;
  assign n15512 = x120 | n15511 ;
  assign n15513 = x120 & n15511 ;
  assign n15514 = n14983 & n23982 ;
  assign n15515 = n135 & n15514 ;
  assign n24192 = ~n14989 ;
  assign n15516 = n24192 & n15515 ;
  assign n24193 = ~n15515 ;
  assign n15517 = n14989 & n24193 ;
  assign n15518 = n15516 | n15517 ;
  assign n24194 = ~n15513 ;
  assign n15519 = n24194 & n15518 ;
  assign n24195 = ~n15519 ;
  assign n15520 = n15512 & n24195 ;
  assign n15522 = x121 | n15520 ;
  assign n24196 = ~n15016 ;
  assign n15523 = n24196 & n15522 ;
  assign n15521 = x121 & n15520 ;
  assign n15007 = x122 & n23990 ;
  assign n15524 = n18283 | n15007 ;
  assign n15525 = n15009 | n15524 ;
  assign n15526 = n15521 | n15525 ;
  assign n15527 = n15523 | n15526 ;
  assign n24197 = ~n15009 ;
  assign n15528 = n24197 & n15527 ;
  assign n134 = ~n15528 ;
  assign n15529 = x64 & n134 ;
  assign n24199 = ~n15529 ;
  assign n15530 = x5 & n24199 ;
  assign n15531 = n15017 & n134 ;
  assign n15532 = n15530 | n15531 ;
  assign n15533 = x65 & n5497 ;
  assign n24200 = ~n15533 ;
  assign n15534 = n15532 & n24200 ;
  assign n24201 = ~n15534 ;
  assign n15535 = n5498 & n24201 ;
  assign n15536 = x66 & n15535 ;
  assign n15537 = n23995 & n15019 ;
  assign n15538 = n134 & n15537 ;
  assign n15539 = n15023 & n15538 ;
  assign n15540 = n15023 | n15538 ;
  assign n24202 = ~n15539 ;
  assign n15541 = n24202 & n15540 ;
  assign n15542 = x66 | n15535 ;
  assign n24203 = ~n15541 ;
  assign n15543 = n24203 & n15542 ;
  assign n15544 = n15536 | n15543 ;
  assign n15545 = x67 & n15544 ;
  assign n15546 = x67 | n15544 ;
  assign n15547 = n15026 & n23998 ;
  assign n15548 = n134 & n15547 ;
  assign n24204 = ~n15032 ;
  assign n15549 = n24204 & n15548 ;
  assign n24205 = ~n15548 ;
  assign n15550 = n15032 & n24205 ;
  assign n15551 = n15549 | n15550 ;
  assign n24206 = ~n15551 ;
  assign n15552 = n15546 & n24206 ;
  assign n15553 = n15545 | n15552 ;
  assign n15554 = x68 & n15553 ;
  assign n15555 = x68 | n15553 ;
  assign n15556 = n15035 & n24002 ;
  assign n15557 = n134 & n15556 ;
  assign n24207 = ~n15041 ;
  assign n15558 = n24207 & n15557 ;
  assign n24208 = ~n15557 ;
  assign n15559 = n15041 & n24208 ;
  assign n15560 = n15558 | n15559 ;
  assign n24209 = ~n15560 ;
  assign n15561 = n15555 & n24209 ;
  assign n15562 = n15554 | n15561 ;
  assign n15563 = x69 & n15562 ;
  assign n15564 = x69 | n15562 ;
  assign n15565 = n15044 & n24006 ;
  assign n15566 = n134 & n15565 ;
  assign n24210 = ~n15050 ;
  assign n15567 = n24210 & n15566 ;
  assign n24211 = ~n15566 ;
  assign n15568 = n15050 & n24211 ;
  assign n15569 = n15567 | n15568 ;
  assign n24212 = ~n15569 ;
  assign n15570 = n15564 & n24212 ;
  assign n15571 = n15563 | n15570 ;
  assign n15572 = x70 & n15571 ;
  assign n15573 = x70 | n15571 ;
  assign n15574 = n15053 & n24010 ;
  assign n15575 = n134 & n15574 ;
  assign n24213 = ~n15059 ;
  assign n15576 = n24213 & n15575 ;
  assign n24214 = ~n15575 ;
  assign n15577 = n15059 & n24214 ;
  assign n15578 = n15576 | n15577 ;
  assign n24215 = ~n15578 ;
  assign n15579 = n15573 & n24215 ;
  assign n15580 = n15572 | n15579 ;
  assign n15581 = x71 & n15580 ;
  assign n15582 = x71 | n15580 ;
  assign n15583 = n15062 & n24014 ;
  assign n15584 = n134 & n15583 ;
  assign n24216 = ~n15068 ;
  assign n15585 = n24216 & n15584 ;
  assign n24217 = ~n15584 ;
  assign n15586 = n15068 & n24217 ;
  assign n15587 = n15585 | n15586 ;
  assign n24218 = ~n15587 ;
  assign n15588 = n15582 & n24218 ;
  assign n15589 = n15581 | n15588 ;
  assign n15590 = x72 & n15589 ;
  assign n15591 = x72 | n15589 ;
  assign n15592 = n15071 & n24017 ;
  assign n15593 = n134 & n15592 ;
  assign n24219 = ~n15077 ;
  assign n15594 = n24219 & n15593 ;
  assign n24220 = ~n15593 ;
  assign n15595 = n15077 & n24220 ;
  assign n15596 = n15594 | n15595 ;
  assign n24221 = ~n15596 ;
  assign n15597 = n15591 & n24221 ;
  assign n15598 = n15590 | n15597 ;
  assign n15599 = x73 & n15598 ;
  assign n15600 = x73 | n15598 ;
  assign n15601 = n15080 & n24021 ;
  assign n15602 = n134 & n15601 ;
  assign n24222 = ~n15086 ;
  assign n15603 = n24222 & n15602 ;
  assign n24223 = ~n15602 ;
  assign n15604 = n15086 & n24223 ;
  assign n15605 = n15603 | n15604 ;
  assign n24224 = ~n15605 ;
  assign n15606 = n15600 & n24224 ;
  assign n15607 = n15599 | n15606 ;
  assign n15608 = x74 & n15607 ;
  assign n15609 = x74 | n15607 ;
  assign n15610 = n15089 & n24024 ;
  assign n15611 = n134 & n15610 ;
  assign n15612 = n15095 & n15611 ;
  assign n15613 = n15095 | n15611 ;
  assign n24225 = ~n15612 ;
  assign n15614 = n24225 & n15613 ;
  assign n24226 = ~n15614 ;
  assign n15615 = n15609 & n24226 ;
  assign n15616 = n15608 | n15615 ;
  assign n15617 = x75 & n15616 ;
  assign n15618 = x75 | n15616 ;
  assign n15619 = n15098 & n24028 ;
  assign n15620 = n134 & n15619 ;
  assign n24227 = ~n15104 ;
  assign n15621 = n24227 & n15620 ;
  assign n24228 = ~n15620 ;
  assign n15622 = n15104 & n24228 ;
  assign n15623 = n15621 | n15622 ;
  assign n24229 = ~n15623 ;
  assign n15624 = n15618 & n24229 ;
  assign n15625 = n15617 | n15624 ;
  assign n15626 = x76 & n15625 ;
  assign n15627 = x76 | n15625 ;
  assign n15628 = n15107 & n24032 ;
  assign n15629 = n134 & n15628 ;
  assign n24230 = ~n15113 ;
  assign n15630 = n24230 & n15629 ;
  assign n24231 = ~n15629 ;
  assign n15631 = n15113 & n24231 ;
  assign n15632 = n15630 | n15631 ;
  assign n24232 = ~n15632 ;
  assign n15633 = n15627 & n24232 ;
  assign n15634 = n15626 | n15633 ;
  assign n15635 = x77 & n15634 ;
  assign n15636 = x77 | n15634 ;
  assign n15637 = n15116 & n24036 ;
  assign n15638 = n134 & n15637 ;
  assign n24233 = ~n15122 ;
  assign n15639 = n24233 & n15638 ;
  assign n24234 = ~n15638 ;
  assign n15640 = n15122 & n24234 ;
  assign n15641 = n15639 | n15640 ;
  assign n24235 = ~n15641 ;
  assign n15642 = n15636 & n24235 ;
  assign n15643 = n15635 | n15642 ;
  assign n15644 = x78 & n15643 ;
  assign n15645 = x78 | n15643 ;
  assign n15646 = n15125 & n24039 ;
  assign n15647 = n134 & n15646 ;
  assign n15648 = n15131 & n15647 ;
  assign n15649 = n15131 | n15647 ;
  assign n24236 = ~n15648 ;
  assign n15650 = n24236 & n15649 ;
  assign n24237 = ~n15650 ;
  assign n15651 = n15645 & n24237 ;
  assign n15652 = n15644 | n15651 ;
  assign n15653 = x79 & n15652 ;
  assign n15654 = x79 | n15652 ;
  assign n15655 = n15134 & n24042 ;
  assign n15656 = n134 & n15655 ;
  assign n24238 = ~n15140 ;
  assign n15657 = n24238 & n15656 ;
  assign n24239 = ~n15656 ;
  assign n15658 = n15140 & n24239 ;
  assign n15659 = n15657 | n15658 ;
  assign n24240 = ~n15659 ;
  assign n15660 = n15654 & n24240 ;
  assign n15661 = n15653 | n15660 ;
  assign n15662 = x80 & n15661 ;
  assign n15663 = x80 | n15661 ;
  assign n15664 = n15143 & n24046 ;
  assign n15665 = n134 & n15664 ;
  assign n24241 = ~n15149 ;
  assign n15666 = n24241 & n15665 ;
  assign n24242 = ~n15665 ;
  assign n15667 = n15149 & n24242 ;
  assign n15668 = n15666 | n15667 ;
  assign n24243 = ~n15668 ;
  assign n15669 = n15663 & n24243 ;
  assign n15670 = n15662 | n15669 ;
  assign n15671 = x81 & n15670 ;
  assign n15672 = x81 | n15670 ;
  assign n15673 = n15152 & n24050 ;
  assign n15674 = n134 & n15673 ;
  assign n24244 = ~n15158 ;
  assign n15675 = n24244 & n15674 ;
  assign n24245 = ~n15674 ;
  assign n15676 = n15158 & n24245 ;
  assign n15677 = n15675 | n15676 ;
  assign n24246 = ~n15677 ;
  assign n15678 = n15672 & n24246 ;
  assign n15679 = n15671 | n15678 ;
  assign n15680 = x82 & n15679 ;
  assign n15681 = x82 | n15679 ;
  assign n15682 = n15161 & n24054 ;
  assign n15683 = n134 & n15682 ;
  assign n24247 = ~n15167 ;
  assign n15684 = n24247 & n15683 ;
  assign n24248 = ~n15683 ;
  assign n15685 = n15167 & n24248 ;
  assign n15686 = n15684 | n15685 ;
  assign n24249 = ~n15686 ;
  assign n15687 = n15681 & n24249 ;
  assign n15688 = n15680 | n15687 ;
  assign n15689 = x83 & n15688 ;
  assign n15690 = x83 | n15688 ;
  assign n15691 = n15170 & n24058 ;
  assign n15692 = n134 & n15691 ;
  assign n15693 = n15176 & n15692 ;
  assign n15694 = n15176 | n15692 ;
  assign n24250 = ~n15693 ;
  assign n15695 = n24250 & n15694 ;
  assign n24251 = ~n15695 ;
  assign n15696 = n15690 & n24251 ;
  assign n15697 = n15689 | n15696 ;
  assign n15698 = x84 & n15697 ;
  assign n15699 = x84 | n15697 ;
  assign n15700 = n15179 & n24062 ;
  assign n15701 = n134 & n15700 ;
  assign n24252 = ~n15185 ;
  assign n15702 = n24252 & n15701 ;
  assign n24253 = ~n15701 ;
  assign n15703 = n15185 & n24253 ;
  assign n15704 = n15702 | n15703 ;
  assign n24254 = ~n15704 ;
  assign n15705 = n15699 & n24254 ;
  assign n15706 = n15698 | n15705 ;
  assign n15707 = x85 & n15706 ;
  assign n15708 = x85 | n15706 ;
  assign n15709 = n15188 & n24066 ;
  assign n15710 = n134 & n15709 ;
  assign n24255 = ~n15194 ;
  assign n15711 = n24255 & n15710 ;
  assign n24256 = ~n15710 ;
  assign n15712 = n15194 & n24256 ;
  assign n15713 = n15711 | n15712 ;
  assign n24257 = ~n15713 ;
  assign n15714 = n15708 & n24257 ;
  assign n15715 = n15707 | n15714 ;
  assign n15716 = x86 & n15715 ;
  assign n15717 = x86 | n15715 ;
  assign n15718 = n15197 & n24069 ;
  assign n15719 = n134 & n15718 ;
  assign n24258 = ~n15203 ;
  assign n15720 = n24258 & n15719 ;
  assign n24259 = ~n15719 ;
  assign n15721 = n15203 & n24259 ;
  assign n15722 = n15720 | n15721 ;
  assign n24260 = ~n15722 ;
  assign n15723 = n15717 & n24260 ;
  assign n15724 = n15716 | n15723 ;
  assign n15725 = x87 & n15724 ;
  assign n15726 = x87 | n15724 ;
  assign n15727 = n15206 & n24072 ;
  assign n15728 = n134 & n15727 ;
  assign n24261 = ~n15212 ;
  assign n15729 = n24261 & n15728 ;
  assign n24262 = ~n15728 ;
  assign n15730 = n15212 & n24262 ;
  assign n15731 = n15729 | n15730 ;
  assign n24263 = ~n15731 ;
  assign n15732 = n15726 & n24263 ;
  assign n15733 = n15725 | n15732 ;
  assign n15734 = x88 & n15733 ;
  assign n15735 = x88 | n15733 ;
  assign n15736 = n15215 & n24075 ;
  assign n15737 = n134 & n15736 ;
  assign n15738 = n15221 & n15737 ;
  assign n15739 = n15221 | n15737 ;
  assign n24264 = ~n15738 ;
  assign n15740 = n24264 & n15739 ;
  assign n24265 = ~n15740 ;
  assign n15741 = n15735 & n24265 ;
  assign n15742 = n15734 | n15741 ;
  assign n15743 = x89 & n15742 ;
  assign n15744 = x89 | n15742 ;
  assign n15745 = n15224 & n24078 ;
  assign n15746 = n134 & n15745 ;
  assign n15747 = n15230 & n15746 ;
  assign n15748 = n15230 | n15746 ;
  assign n24266 = ~n15747 ;
  assign n15749 = n24266 & n15748 ;
  assign n24267 = ~n15749 ;
  assign n15750 = n15744 & n24267 ;
  assign n15751 = n15743 | n15750 ;
  assign n15752 = x90 & n15751 ;
  assign n15753 = x90 | n15751 ;
  assign n15754 = n15233 & n24081 ;
  assign n15755 = n134 & n15754 ;
  assign n24268 = ~n15239 ;
  assign n15756 = n24268 & n15755 ;
  assign n24269 = ~n15755 ;
  assign n15757 = n15239 & n24269 ;
  assign n15758 = n15756 | n15757 ;
  assign n24270 = ~n15758 ;
  assign n15759 = n15753 & n24270 ;
  assign n15760 = n15752 | n15759 ;
  assign n15761 = x91 & n15760 ;
  assign n15762 = x91 | n15760 ;
  assign n15763 = n15242 & n24085 ;
  assign n15764 = n134 & n15763 ;
  assign n15765 = n15248 & n15764 ;
  assign n15766 = n15248 | n15764 ;
  assign n24271 = ~n15765 ;
  assign n15767 = n24271 & n15766 ;
  assign n24272 = ~n15767 ;
  assign n15768 = n15762 & n24272 ;
  assign n15769 = n15761 | n15768 ;
  assign n15770 = x92 & n15769 ;
  assign n15771 = x92 | n15769 ;
  assign n15772 = n15251 & n24089 ;
  assign n15773 = n134 & n15772 ;
  assign n24273 = ~n15257 ;
  assign n15774 = n24273 & n15773 ;
  assign n24274 = ~n15773 ;
  assign n15775 = n15257 & n24274 ;
  assign n15776 = n15774 | n15775 ;
  assign n24275 = ~n15776 ;
  assign n15777 = n15771 & n24275 ;
  assign n15778 = n15770 | n15777 ;
  assign n15779 = x93 & n15778 ;
  assign n15780 = x93 | n15778 ;
  assign n15781 = n15260 & n24092 ;
  assign n15782 = n134 & n15781 ;
  assign n15783 = n15266 & n15782 ;
  assign n15784 = n15266 | n15782 ;
  assign n24276 = ~n15783 ;
  assign n15785 = n24276 & n15784 ;
  assign n24277 = ~n15785 ;
  assign n15786 = n15780 & n24277 ;
  assign n15787 = n15779 | n15786 ;
  assign n15788 = x94 & n15787 ;
  assign n15789 = x94 | n15787 ;
  assign n15790 = n15269 & n24095 ;
  assign n15791 = n134 & n15790 ;
  assign n15792 = n15275 & n15791 ;
  assign n15793 = n15275 | n15791 ;
  assign n24278 = ~n15792 ;
  assign n15794 = n24278 & n15793 ;
  assign n24279 = ~n15794 ;
  assign n15795 = n15789 & n24279 ;
  assign n15796 = n15788 | n15795 ;
  assign n15797 = x95 & n15796 ;
  assign n15798 = x95 | n15796 ;
  assign n15799 = n15278 & n24098 ;
  assign n15800 = n134 & n15799 ;
  assign n15801 = n15284 & n15800 ;
  assign n15802 = n15284 | n15800 ;
  assign n24280 = ~n15801 ;
  assign n15803 = n24280 & n15802 ;
  assign n24281 = ~n15803 ;
  assign n15804 = n15798 & n24281 ;
  assign n15805 = n15797 | n15804 ;
  assign n15806 = x96 & n15805 ;
  assign n15807 = x96 | n15805 ;
  assign n15808 = n15287 & n24102 ;
  assign n15809 = n134 & n15808 ;
  assign n24282 = ~n15293 ;
  assign n15810 = n24282 & n15809 ;
  assign n24283 = ~n15809 ;
  assign n15811 = n15293 & n24283 ;
  assign n15812 = n15810 | n15811 ;
  assign n24284 = ~n15812 ;
  assign n15813 = n15807 & n24284 ;
  assign n15814 = n15806 | n15813 ;
  assign n15815 = x97 & n15814 ;
  assign n15816 = x97 | n15814 ;
  assign n15817 = n15296 & n24105 ;
  assign n15818 = n134 & n15817 ;
  assign n24285 = ~n15302 ;
  assign n15819 = n24285 & n15818 ;
  assign n24286 = ~n15818 ;
  assign n15820 = n15302 & n24286 ;
  assign n15821 = n15819 | n15820 ;
  assign n24287 = ~n15821 ;
  assign n15822 = n15816 & n24287 ;
  assign n15823 = n15815 | n15822 ;
  assign n15824 = x98 & n15823 ;
  assign n15825 = x98 | n15823 ;
  assign n15826 = n15305 & n24109 ;
  assign n15827 = n134 & n15826 ;
  assign n24288 = ~n15311 ;
  assign n15828 = n24288 & n15827 ;
  assign n24289 = ~n15827 ;
  assign n15829 = n15311 & n24289 ;
  assign n15830 = n15828 | n15829 ;
  assign n24290 = ~n15830 ;
  assign n15831 = n15825 & n24290 ;
  assign n15832 = n15824 | n15831 ;
  assign n15833 = x99 & n15832 ;
  assign n15834 = x99 | n15832 ;
  assign n15835 = n15314 & n24112 ;
  assign n15836 = n134 & n15835 ;
  assign n24291 = ~n15320 ;
  assign n15837 = n24291 & n15836 ;
  assign n24292 = ~n15836 ;
  assign n15838 = n15320 & n24292 ;
  assign n15839 = n15837 | n15838 ;
  assign n24293 = ~n15839 ;
  assign n15840 = n15834 & n24293 ;
  assign n15841 = n15833 | n15840 ;
  assign n15842 = x100 & n15841 ;
  assign n15843 = x100 | n15841 ;
  assign n15844 = n15323 & n24116 ;
  assign n15845 = n134 & n15844 ;
  assign n15846 = n15329 & n15845 ;
  assign n15847 = n15329 | n15845 ;
  assign n24294 = ~n15846 ;
  assign n15848 = n24294 & n15847 ;
  assign n24295 = ~n15848 ;
  assign n15849 = n15843 & n24295 ;
  assign n15850 = n15842 | n15849 ;
  assign n15851 = x101 & n15850 ;
  assign n15852 = x101 | n15850 ;
  assign n15853 = n15332 & n24120 ;
  assign n15854 = n134 & n15853 ;
  assign n24296 = ~n15338 ;
  assign n15855 = n24296 & n15854 ;
  assign n24297 = ~n15854 ;
  assign n15856 = n15338 & n24297 ;
  assign n15857 = n15855 | n15856 ;
  assign n24298 = ~n15857 ;
  assign n15858 = n15852 & n24298 ;
  assign n15859 = n15851 | n15858 ;
  assign n15860 = x102 & n15859 ;
  assign n15861 = x102 | n15859 ;
  assign n15862 = n15341 & n24124 ;
  assign n15863 = n134 & n15862 ;
  assign n24299 = ~n15347 ;
  assign n15864 = n24299 & n15863 ;
  assign n24300 = ~n15863 ;
  assign n15865 = n15347 & n24300 ;
  assign n15866 = n15864 | n15865 ;
  assign n24301 = ~n15866 ;
  assign n15867 = n15861 & n24301 ;
  assign n15868 = n15860 | n15867 ;
  assign n15869 = x103 & n15868 ;
  assign n15870 = x103 | n15868 ;
  assign n15871 = n15350 & n24127 ;
  assign n15872 = n134 & n15871 ;
  assign n24302 = ~n15356 ;
  assign n15873 = n24302 & n15872 ;
  assign n24303 = ~n15872 ;
  assign n15874 = n15356 & n24303 ;
  assign n15875 = n15873 | n15874 ;
  assign n24304 = ~n15875 ;
  assign n15876 = n15870 & n24304 ;
  assign n15877 = n15869 | n15876 ;
  assign n15878 = x104 & n15877 ;
  assign n15879 = x104 | n15877 ;
  assign n15880 = n15359 & n24131 ;
  assign n15881 = n134 & n15880 ;
  assign n24305 = ~n15365 ;
  assign n15882 = n24305 & n15881 ;
  assign n24306 = ~n15881 ;
  assign n15883 = n15365 & n24306 ;
  assign n15884 = n15882 | n15883 ;
  assign n24307 = ~n15884 ;
  assign n15885 = n15879 & n24307 ;
  assign n15886 = n15878 | n15885 ;
  assign n15887 = x105 & n15886 ;
  assign n15888 = x105 | n15886 ;
  assign n15889 = n15368 & n24135 ;
  assign n15890 = n134 & n15889 ;
  assign n24308 = ~n15374 ;
  assign n15891 = n24308 & n15890 ;
  assign n24309 = ~n15890 ;
  assign n15892 = n15374 & n24309 ;
  assign n15893 = n15891 | n15892 ;
  assign n24310 = ~n15893 ;
  assign n15894 = n15888 & n24310 ;
  assign n15895 = n15887 | n15894 ;
  assign n15896 = x106 & n15895 ;
  assign n15897 = x106 | n15895 ;
  assign n15898 = n15377 & n24138 ;
  assign n15899 = n134 & n15898 ;
  assign n24311 = ~n15383 ;
  assign n15900 = n24311 & n15899 ;
  assign n24312 = ~n15899 ;
  assign n15901 = n15383 & n24312 ;
  assign n15902 = n15900 | n15901 ;
  assign n24313 = ~n15902 ;
  assign n15903 = n15897 & n24313 ;
  assign n15904 = n15896 | n15903 ;
  assign n15905 = x107 & n15904 ;
  assign n15906 = x107 | n15904 ;
  assign n15907 = n15386 & n24142 ;
  assign n15908 = n134 & n15907 ;
  assign n24314 = ~n15392 ;
  assign n15909 = n24314 & n15908 ;
  assign n24315 = ~n15908 ;
  assign n15910 = n15392 & n24315 ;
  assign n15911 = n15909 | n15910 ;
  assign n24316 = ~n15911 ;
  assign n15912 = n15906 & n24316 ;
  assign n15913 = n15905 | n15912 ;
  assign n15914 = x108 & n15913 ;
  assign n15915 = x108 | n15913 ;
  assign n15916 = n15395 & n24146 ;
  assign n15917 = n134 & n15916 ;
  assign n24317 = ~n15401 ;
  assign n15918 = n24317 & n15917 ;
  assign n24318 = ~n15917 ;
  assign n15919 = n15401 & n24318 ;
  assign n15920 = n15918 | n15919 ;
  assign n24319 = ~n15920 ;
  assign n15921 = n15915 & n24319 ;
  assign n15922 = n15914 | n15921 ;
  assign n15923 = x109 & n15922 ;
  assign n15924 = x109 | n15922 ;
  assign n15925 = n15404 & n24150 ;
  assign n15926 = n134 & n15925 ;
  assign n15927 = n15410 & n15926 ;
  assign n15928 = n15410 | n15926 ;
  assign n24320 = ~n15927 ;
  assign n15929 = n24320 & n15928 ;
  assign n24321 = ~n15929 ;
  assign n15930 = n15924 & n24321 ;
  assign n15931 = n15923 | n15930 ;
  assign n15932 = x110 & n15931 ;
  assign n15933 = x110 | n15931 ;
  assign n15934 = n15413 & n24153 ;
  assign n15935 = n134 & n15934 ;
  assign n15936 = n15419 & n15935 ;
  assign n15937 = n15419 | n15935 ;
  assign n24322 = ~n15936 ;
  assign n15938 = n24322 & n15937 ;
  assign n24323 = ~n15938 ;
  assign n15939 = n15933 & n24323 ;
  assign n15940 = n15932 | n15939 ;
  assign n15941 = x111 & n15940 ;
  assign n15942 = x111 | n15940 ;
  assign n15943 = n15422 & n24156 ;
  assign n15944 = n134 & n15943 ;
  assign n15945 = n15428 & n15944 ;
  assign n15946 = n15428 | n15944 ;
  assign n24324 = ~n15945 ;
  assign n15947 = n24324 & n15946 ;
  assign n24325 = ~n15947 ;
  assign n15948 = n15942 & n24325 ;
  assign n15949 = n15941 | n15948 ;
  assign n15950 = x112 & n15949 ;
  assign n15951 = x112 | n15949 ;
  assign n15952 = n15431 & n24160 ;
  assign n15953 = n134 & n15952 ;
  assign n24326 = ~n15437 ;
  assign n15954 = n24326 & n15953 ;
  assign n24327 = ~n15953 ;
  assign n15955 = n15437 & n24327 ;
  assign n15956 = n15954 | n15955 ;
  assign n24328 = ~n15956 ;
  assign n15957 = n15951 & n24328 ;
  assign n15958 = n15950 | n15957 ;
  assign n15959 = x113 & n15958 ;
  assign n15960 = x113 | n15958 ;
  assign n15961 = n15440 & n24164 ;
  assign n15962 = n134 & n15961 ;
  assign n24329 = ~n15446 ;
  assign n15963 = n24329 & n15962 ;
  assign n24330 = ~n15962 ;
  assign n15964 = n15446 & n24330 ;
  assign n15965 = n15963 | n15964 ;
  assign n24331 = ~n15965 ;
  assign n15966 = n15960 & n24331 ;
  assign n15967 = n15959 | n15966 ;
  assign n15968 = x114 & n15967 ;
  assign n15969 = x114 | n15967 ;
  assign n15970 = n15449 & n24168 ;
  assign n15971 = n134 & n15970 ;
  assign n24332 = ~n15455 ;
  assign n15972 = n24332 & n15971 ;
  assign n24333 = ~n15971 ;
  assign n15973 = n15455 & n24333 ;
  assign n15974 = n15972 | n15973 ;
  assign n24334 = ~n15974 ;
  assign n15975 = n15969 & n24334 ;
  assign n15976 = n15968 | n15975 ;
  assign n15977 = x115 & n15976 ;
  assign n15978 = x115 | n15976 ;
  assign n15979 = n15458 & n24172 ;
  assign n15980 = n134 & n15979 ;
  assign n24335 = ~n15464 ;
  assign n15981 = n24335 & n15980 ;
  assign n24336 = ~n15980 ;
  assign n15982 = n15464 & n24336 ;
  assign n15983 = n15981 | n15982 ;
  assign n24337 = ~n15983 ;
  assign n15984 = n15978 & n24337 ;
  assign n15985 = n15977 | n15984 ;
  assign n15986 = x116 & n15985 ;
  assign n15987 = x116 | n15985 ;
  assign n15988 = n15467 & n24176 ;
  assign n15989 = n134 & n15988 ;
  assign n24338 = ~n15473 ;
  assign n15990 = n24338 & n15989 ;
  assign n24339 = ~n15989 ;
  assign n15991 = n15473 & n24339 ;
  assign n15992 = n15990 | n15991 ;
  assign n24340 = ~n15992 ;
  assign n15993 = n15987 & n24340 ;
  assign n15994 = n15986 | n15993 ;
  assign n15995 = x117 & n15994 ;
  assign n15996 = x117 | n15994 ;
  assign n15997 = n15476 & n24180 ;
  assign n15998 = n134 & n15997 ;
  assign n24341 = ~n15482 ;
  assign n15999 = n24341 & n15998 ;
  assign n24342 = ~n15998 ;
  assign n16000 = n15482 & n24342 ;
  assign n16001 = n15999 | n16000 ;
  assign n24343 = ~n16001 ;
  assign n16002 = n15996 & n24343 ;
  assign n16003 = n15995 | n16002 ;
  assign n16004 = x118 & n16003 ;
  assign n16005 = x118 | n16003 ;
  assign n16006 = n15485 & n24184 ;
  assign n16007 = n134 & n16006 ;
  assign n16008 = n15491 & n16007 ;
  assign n16009 = n15491 | n16007 ;
  assign n24344 = ~n16008 ;
  assign n16010 = n24344 & n16009 ;
  assign n24345 = ~n16010 ;
  assign n16011 = n16005 & n24345 ;
  assign n16012 = n16004 | n16011 ;
  assign n16013 = x119 & n16012 ;
  assign n16014 = x119 | n16012 ;
  assign n16015 = n15494 & n24187 ;
  assign n16016 = n134 & n16015 ;
  assign n16017 = n15500 & n16016 ;
  assign n16018 = n15500 | n16016 ;
  assign n24346 = ~n16017 ;
  assign n16019 = n24346 & n16018 ;
  assign n24347 = ~n16019 ;
  assign n16020 = n16014 & n24347 ;
  assign n16021 = n16013 | n16020 ;
  assign n16022 = x120 & n16021 ;
  assign n16023 = x120 | n16021 ;
  assign n16024 = n15503 & n24190 ;
  assign n16025 = n134 & n16024 ;
  assign n24348 = ~n15509 ;
  assign n16026 = n24348 & n16025 ;
  assign n24349 = ~n16025 ;
  assign n16027 = n15509 & n24349 ;
  assign n16028 = n16026 | n16027 ;
  assign n24350 = ~n16028 ;
  assign n16029 = n16023 & n24350 ;
  assign n16030 = n16022 | n16029 ;
  assign n16031 = x121 & n16030 ;
  assign n16032 = x121 | n16030 ;
  assign n16033 = n15512 & n24194 ;
  assign n16034 = n134 & n16033 ;
  assign n24351 = ~n15518 ;
  assign n16035 = n24351 & n16034 ;
  assign n24352 = ~n16034 ;
  assign n16036 = n15518 & n24352 ;
  assign n16037 = n16035 | n16036 ;
  assign n24353 = ~n16037 ;
  assign n16038 = n16032 & n24353 ;
  assign n16039 = n16031 | n16038 ;
  assign n16040 = x122 & n16039 ;
  assign n16041 = x122 | n16039 ;
  assign n24354 = ~n15521 ;
  assign n16042 = n24354 & n15522 ;
  assign n16043 = n134 & n16042 ;
  assign n16044 = n24196 & n16043 ;
  assign n24355 = ~n16043 ;
  assign n16045 = n15016 & n24355 ;
  assign n16046 = n16044 | n16045 ;
  assign n24356 = ~n16046 ;
  assign n16047 = n16041 & n24356 ;
  assign n16048 = n16040 | n16047 ;
  assign n16049 = x123 | n16048 ;
  assign n16050 = x123 & n16048 ;
  assign n16051 = n18278 | n16050 ;
  assign n24357 = ~n16051 ;
  assign n16052 = n16049 & n24357 ;
  assign n16053 = n18288 & n15005 ;
  assign n16054 = n15527 & n16053 ;
  assign n16055 = n21884 | n16054 ;
  assign n24358 = ~n16052 ;
  assign n16057 = n24358 & n16055 ;
  assign n16058 = n18273 & n16057 ;
  assign n24359 = ~x2 ;
  assign n5494 = n24359 & x64 ;
  assign n5495 = x65 | n5494 ;
  assign n5496 = x65 & n5494 ;
  assign n24360 = ~n16055 ;
  assign n16056 = n16049 & n24360 ;
  assign n16063 = n16051 | n16056 ;
  assign n24361 = ~n16040 ;
  assign n16584 = n24361 & n16041 ;
  assign n133 = ~n16063 ;
  assign n16585 = n133 & n16584 ;
  assign n16586 = n24356 & n16585 ;
  assign n24363 = ~n16585 ;
  assign n16587 = n16046 & n24363 ;
  assign n16588 = n16586 | n16587 ;
  assign n24364 = ~x3 ;
  assign n16060 = n24364 & x64 ;
  assign n16062 = x65 | n16060 ;
  assign n16061 = x65 & n16060 ;
  assign n16064 = x64 & n133 ;
  assign n16065 = x4 & n16064 ;
  assign n16066 = x4 | n16064 ;
  assign n24365 = ~n16065 ;
  assign n16067 = n24365 & n16066 ;
  assign n24366 = ~n16061 ;
  assign n16068 = n24366 & n16067 ;
  assign n24367 = ~n16068 ;
  assign n16069 = n16062 & n24367 ;
  assign n16070 = x66 | n16069 ;
  assign n16071 = x66 & n16069 ;
  assign n16072 = n5498 & n133 ;
  assign n16073 = n24200 & n16072 ;
  assign n16074 = n15532 | n16073 ;
  assign n16075 = n15534 & n16072 ;
  assign n24368 = ~n16075 ;
  assign n16076 = n16074 & n24368 ;
  assign n24369 = ~n16071 ;
  assign n16077 = n24369 & n16076 ;
  assign n24370 = ~n16077 ;
  assign n16078 = n16070 & n24370 ;
  assign n16079 = x67 | n16078 ;
  assign n16080 = x67 & n16078 ;
  assign n24371 = ~n15536 ;
  assign n16081 = n24371 & n15542 ;
  assign n16082 = n133 & n16081 ;
  assign n16083 = n15541 & n16082 ;
  assign n16084 = n15541 | n16082 ;
  assign n24372 = ~n16083 ;
  assign n16085 = n24372 & n16084 ;
  assign n24373 = ~n16080 ;
  assign n16086 = n24373 & n16085 ;
  assign n24374 = ~n16086 ;
  assign n16087 = n16079 & n24374 ;
  assign n16088 = x68 | n16087 ;
  assign n16089 = x68 & n16087 ;
  assign n24375 = ~n15545 ;
  assign n16090 = n24375 & n15546 ;
  assign n16091 = n133 & n16090 ;
  assign n16092 = n15551 & n16091 ;
  assign n16093 = n15551 | n16091 ;
  assign n24376 = ~n16092 ;
  assign n16094 = n24376 & n16093 ;
  assign n24377 = ~n16089 ;
  assign n16095 = n24377 & n16094 ;
  assign n24378 = ~n16095 ;
  assign n16096 = n16088 & n24378 ;
  assign n16097 = x69 | n16096 ;
  assign n16098 = x69 & n16096 ;
  assign n24379 = ~n15554 ;
  assign n16099 = n24379 & n15555 ;
  assign n16100 = n133 & n16099 ;
  assign n16101 = n24209 & n16100 ;
  assign n24380 = ~n16100 ;
  assign n16102 = n15560 & n24380 ;
  assign n16103 = n16101 | n16102 ;
  assign n24381 = ~n16098 ;
  assign n16104 = n24381 & n16103 ;
  assign n24382 = ~n16104 ;
  assign n16105 = n16097 & n24382 ;
  assign n16106 = x70 | n16105 ;
  assign n16107 = x70 & n16105 ;
  assign n24383 = ~n15563 ;
  assign n16108 = n24383 & n15564 ;
  assign n16109 = n133 & n16108 ;
  assign n16110 = n15569 & n16109 ;
  assign n16111 = n15569 | n16109 ;
  assign n24384 = ~n16110 ;
  assign n16112 = n24384 & n16111 ;
  assign n24385 = ~n16107 ;
  assign n16113 = n24385 & n16112 ;
  assign n24386 = ~n16113 ;
  assign n16114 = n16106 & n24386 ;
  assign n16115 = x71 | n16114 ;
  assign n16116 = x71 & n16114 ;
  assign n24387 = ~n15572 ;
  assign n16117 = n24387 & n15573 ;
  assign n16118 = n133 & n16117 ;
  assign n16119 = n15578 & n16118 ;
  assign n16120 = n15578 | n16118 ;
  assign n24388 = ~n16119 ;
  assign n16121 = n24388 & n16120 ;
  assign n24389 = ~n16116 ;
  assign n16122 = n24389 & n16121 ;
  assign n24390 = ~n16122 ;
  assign n16123 = n16115 & n24390 ;
  assign n16124 = x72 | n16123 ;
  assign n16125 = x72 & n16123 ;
  assign n24391 = ~n15581 ;
  assign n16126 = n24391 & n15582 ;
  assign n16127 = n133 & n16126 ;
  assign n16128 = n15587 & n16127 ;
  assign n16129 = n15587 | n16127 ;
  assign n24392 = ~n16128 ;
  assign n16130 = n24392 & n16129 ;
  assign n24393 = ~n16125 ;
  assign n16131 = n24393 & n16130 ;
  assign n24394 = ~n16131 ;
  assign n16132 = n16124 & n24394 ;
  assign n16133 = x73 | n16132 ;
  assign n16134 = x73 & n16132 ;
  assign n24395 = ~n15590 ;
  assign n16135 = n24395 & n15591 ;
  assign n16136 = n133 & n16135 ;
  assign n16137 = n24221 & n16136 ;
  assign n24396 = ~n16136 ;
  assign n16138 = n15596 & n24396 ;
  assign n16139 = n16137 | n16138 ;
  assign n24397 = ~n16134 ;
  assign n16140 = n24397 & n16139 ;
  assign n24398 = ~n16140 ;
  assign n16141 = n16133 & n24398 ;
  assign n16142 = x74 | n16141 ;
  assign n16143 = x74 & n16141 ;
  assign n24399 = ~n15599 ;
  assign n16144 = n24399 & n15600 ;
  assign n16145 = n133 & n16144 ;
  assign n16146 = n24224 & n16145 ;
  assign n24400 = ~n16145 ;
  assign n16147 = n15605 & n24400 ;
  assign n16148 = n16146 | n16147 ;
  assign n24401 = ~n16143 ;
  assign n16149 = n24401 & n16148 ;
  assign n24402 = ~n16149 ;
  assign n16150 = n16142 & n24402 ;
  assign n16151 = x75 | n16150 ;
  assign n16152 = x75 & n16150 ;
  assign n24403 = ~n15608 ;
  assign n16153 = n24403 & n15609 ;
  assign n16154 = n133 & n16153 ;
  assign n16155 = n15614 & n16154 ;
  assign n16156 = n15614 | n16154 ;
  assign n24404 = ~n16155 ;
  assign n16157 = n24404 & n16156 ;
  assign n24405 = ~n16152 ;
  assign n16158 = n24405 & n16157 ;
  assign n24406 = ~n16158 ;
  assign n16159 = n16151 & n24406 ;
  assign n16160 = x76 | n16159 ;
  assign n16161 = x76 & n16159 ;
  assign n24407 = ~n15617 ;
  assign n16162 = n24407 & n15618 ;
  assign n16163 = n133 & n16162 ;
  assign n16164 = n15623 & n16163 ;
  assign n16165 = n15623 | n16163 ;
  assign n24408 = ~n16164 ;
  assign n16166 = n24408 & n16165 ;
  assign n24409 = ~n16161 ;
  assign n16167 = n24409 & n16166 ;
  assign n24410 = ~n16167 ;
  assign n16168 = n16160 & n24410 ;
  assign n16169 = x77 | n16168 ;
  assign n16170 = x77 & n16168 ;
  assign n24411 = ~n15626 ;
  assign n16171 = n24411 & n15627 ;
  assign n16172 = n133 & n16171 ;
  assign n16173 = n15632 & n16172 ;
  assign n16174 = n15632 | n16172 ;
  assign n24412 = ~n16173 ;
  assign n16175 = n24412 & n16174 ;
  assign n24413 = ~n16170 ;
  assign n16176 = n24413 & n16175 ;
  assign n24414 = ~n16176 ;
  assign n16177 = n16169 & n24414 ;
  assign n16178 = x78 | n16177 ;
  assign n16179 = x78 & n16177 ;
  assign n24415 = ~n15635 ;
  assign n16180 = n24415 & n15636 ;
  assign n16181 = n133 & n16180 ;
  assign n16182 = n15641 & n16181 ;
  assign n16183 = n15641 | n16181 ;
  assign n24416 = ~n16182 ;
  assign n16184 = n24416 & n16183 ;
  assign n24417 = ~n16179 ;
  assign n16185 = n24417 & n16184 ;
  assign n24418 = ~n16185 ;
  assign n16186 = n16178 & n24418 ;
  assign n16187 = x79 | n16186 ;
  assign n16188 = x79 & n16186 ;
  assign n24419 = ~n15644 ;
  assign n16189 = n24419 & n15645 ;
  assign n16190 = n133 & n16189 ;
  assign n16191 = n15650 & n16190 ;
  assign n16192 = n15650 | n16190 ;
  assign n24420 = ~n16191 ;
  assign n16193 = n24420 & n16192 ;
  assign n24421 = ~n16188 ;
  assign n16194 = n24421 & n16193 ;
  assign n24422 = ~n16194 ;
  assign n16195 = n16187 & n24422 ;
  assign n16196 = x80 | n16195 ;
  assign n16197 = x80 & n16195 ;
  assign n24423 = ~n15653 ;
  assign n16198 = n24423 & n15654 ;
  assign n16199 = n133 & n16198 ;
  assign n16200 = n24240 & n16199 ;
  assign n24424 = ~n16199 ;
  assign n16201 = n15659 & n24424 ;
  assign n16202 = n16200 | n16201 ;
  assign n24425 = ~n16197 ;
  assign n16203 = n24425 & n16202 ;
  assign n24426 = ~n16203 ;
  assign n16204 = n16196 & n24426 ;
  assign n16205 = x81 | n16204 ;
  assign n16206 = x81 & n16204 ;
  assign n24427 = ~n15662 ;
  assign n16207 = n24427 & n15663 ;
  assign n16208 = n133 & n16207 ;
  assign n16209 = n24243 & n16208 ;
  assign n24428 = ~n16208 ;
  assign n16210 = n15668 & n24428 ;
  assign n16211 = n16209 | n16210 ;
  assign n24429 = ~n16206 ;
  assign n16212 = n24429 & n16211 ;
  assign n24430 = ~n16212 ;
  assign n16213 = n16205 & n24430 ;
  assign n16214 = x82 | n16213 ;
  assign n16215 = x82 & n16213 ;
  assign n24431 = ~n15671 ;
  assign n16216 = n24431 & n15672 ;
  assign n16217 = n133 & n16216 ;
  assign n16218 = n15677 & n16217 ;
  assign n16219 = n15677 | n16217 ;
  assign n24432 = ~n16218 ;
  assign n16220 = n24432 & n16219 ;
  assign n24433 = ~n16215 ;
  assign n16221 = n24433 & n16220 ;
  assign n24434 = ~n16221 ;
  assign n16222 = n16214 & n24434 ;
  assign n16223 = x83 | n16222 ;
  assign n16224 = x83 & n16222 ;
  assign n24435 = ~n15680 ;
  assign n16225 = n24435 & n15681 ;
  assign n16226 = n133 & n16225 ;
  assign n16227 = n24249 & n16226 ;
  assign n24436 = ~n16226 ;
  assign n16228 = n15686 & n24436 ;
  assign n16229 = n16227 | n16228 ;
  assign n24437 = ~n16224 ;
  assign n16230 = n24437 & n16229 ;
  assign n24438 = ~n16230 ;
  assign n16231 = n16223 & n24438 ;
  assign n16232 = x84 | n16231 ;
  assign n16233 = x84 & n16231 ;
  assign n24439 = ~n15689 ;
  assign n16234 = n24439 & n15690 ;
  assign n16235 = n133 & n16234 ;
  assign n16236 = n15695 & n16235 ;
  assign n16237 = n15695 | n16235 ;
  assign n24440 = ~n16236 ;
  assign n16238 = n24440 & n16237 ;
  assign n24441 = ~n16233 ;
  assign n16239 = n24441 & n16238 ;
  assign n24442 = ~n16239 ;
  assign n16240 = n16232 & n24442 ;
  assign n16241 = x85 | n16240 ;
  assign n16242 = x85 & n16240 ;
  assign n24443 = ~n15698 ;
  assign n16243 = n24443 & n15699 ;
  assign n16244 = n133 & n16243 ;
  assign n16245 = n15704 & n16244 ;
  assign n16246 = n15704 | n16244 ;
  assign n24444 = ~n16245 ;
  assign n16247 = n24444 & n16246 ;
  assign n24445 = ~n16242 ;
  assign n16248 = n24445 & n16247 ;
  assign n24446 = ~n16248 ;
  assign n16249 = n16241 & n24446 ;
  assign n16250 = x86 | n16249 ;
  assign n16251 = x86 & n16249 ;
  assign n24447 = ~n15707 ;
  assign n16252 = n24447 & n15708 ;
  assign n16253 = n133 & n16252 ;
  assign n16254 = n15713 & n16253 ;
  assign n16255 = n15713 | n16253 ;
  assign n24448 = ~n16254 ;
  assign n16256 = n24448 & n16255 ;
  assign n24449 = ~n16251 ;
  assign n16257 = n24449 & n16256 ;
  assign n24450 = ~n16257 ;
  assign n16258 = n16250 & n24450 ;
  assign n16259 = x87 | n16258 ;
  assign n16260 = x87 & n16258 ;
  assign n24451 = ~n15716 ;
  assign n16261 = n24451 & n15717 ;
  assign n16262 = n133 & n16261 ;
  assign n16263 = n24260 & n16262 ;
  assign n24452 = ~n16262 ;
  assign n16264 = n15722 & n24452 ;
  assign n16265 = n16263 | n16264 ;
  assign n24453 = ~n16260 ;
  assign n16266 = n24453 & n16265 ;
  assign n24454 = ~n16266 ;
  assign n16267 = n16259 & n24454 ;
  assign n16268 = x88 | n16267 ;
  assign n16269 = x88 & n16267 ;
  assign n24455 = ~n15725 ;
  assign n16270 = n24455 & n15726 ;
  assign n16271 = n133 & n16270 ;
  assign n16272 = n24263 & n16271 ;
  assign n24456 = ~n16271 ;
  assign n16273 = n15731 & n24456 ;
  assign n16274 = n16272 | n16273 ;
  assign n24457 = ~n16269 ;
  assign n16275 = n24457 & n16274 ;
  assign n24458 = ~n16275 ;
  assign n16276 = n16268 & n24458 ;
  assign n16277 = x89 | n16276 ;
  assign n16278 = x89 & n16276 ;
  assign n24459 = ~n15734 ;
  assign n16279 = n24459 & n15735 ;
  assign n16280 = n133 & n16279 ;
  assign n16281 = n15740 & n16280 ;
  assign n16282 = n15740 | n16280 ;
  assign n24460 = ~n16281 ;
  assign n16283 = n24460 & n16282 ;
  assign n24461 = ~n16278 ;
  assign n16284 = n24461 & n16283 ;
  assign n24462 = ~n16284 ;
  assign n16285 = n16277 & n24462 ;
  assign n16286 = x90 | n16285 ;
  assign n16287 = x90 & n16285 ;
  assign n24463 = ~n15743 ;
  assign n16288 = n24463 & n15744 ;
  assign n16289 = n133 & n16288 ;
  assign n16290 = n15749 & n16289 ;
  assign n16291 = n15749 | n16289 ;
  assign n24464 = ~n16290 ;
  assign n16292 = n24464 & n16291 ;
  assign n24465 = ~n16287 ;
  assign n16293 = n24465 & n16292 ;
  assign n24466 = ~n16293 ;
  assign n16294 = n16286 & n24466 ;
  assign n16295 = x91 | n16294 ;
  assign n16296 = x91 & n16294 ;
  assign n24467 = ~n15752 ;
  assign n16297 = n24467 & n15753 ;
  assign n16298 = n133 & n16297 ;
  assign n16299 = n24270 & n16298 ;
  assign n24468 = ~n16298 ;
  assign n16300 = n15758 & n24468 ;
  assign n16301 = n16299 | n16300 ;
  assign n24469 = ~n16296 ;
  assign n16302 = n24469 & n16301 ;
  assign n24470 = ~n16302 ;
  assign n16303 = n16295 & n24470 ;
  assign n16304 = x92 | n16303 ;
  assign n16305 = x92 & n16303 ;
  assign n24471 = ~n15761 ;
  assign n16306 = n24471 & n15762 ;
  assign n16307 = n133 & n16306 ;
  assign n16308 = n15767 & n16307 ;
  assign n16309 = n15767 | n16307 ;
  assign n24472 = ~n16308 ;
  assign n16310 = n24472 & n16309 ;
  assign n24473 = ~n16305 ;
  assign n16311 = n24473 & n16310 ;
  assign n24474 = ~n16311 ;
  assign n16312 = n16304 & n24474 ;
  assign n16313 = x93 | n16312 ;
  assign n16314 = x93 & n16312 ;
  assign n24475 = ~n15770 ;
  assign n16315 = n24475 & n15771 ;
  assign n16316 = n133 & n16315 ;
  assign n16317 = n15776 & n16316 ;
  assign n16318 = n15776 | n16316 ;
  assign n24476 = ~n16317 ;
  assign n16319 = n24476 & n16318 ;
  assign n24477 = ~n16314 ;
  assign n16320 = n24477 & n16319 ;
  assign n24478 = ~n16320 ;
  assign n16321 = n16313 & n24478 ;
  assign n16322 = x94 | n16321 ;
  assign n16323 = x94 & n16321 ;
  assign n24479 = ~n15779 ;
  assign n16324 = n24479 & n15780 ;
  assign n16325 = n133 & n16324 ;
  assign n16326 = n15785 & n16325 ;
  assign n16327 = n15785 | n16325 ;
  assign n24480 = ~n16326 ;
  assign n16328 = n24480 & n16327 ;
  assign n24481 = ~n16323 ;
  assign n16329 = n24481 & n16328 ;
  assign n24482 = ~n16329 ;
  assign n16330 = n16322 & n24482 ;
  assign n16331 = x95 | n16330 ;
  assign n16332 = x95 & n16330 ;
  assign n24483 = ~n15788 ;
  assign n16333 = n24483 & n15789 ;
  assign n16334 = n133 & n16333 ;
  assign n16335 = n15794 & n16334 ;
  assign n16336 = n15794 | n16334 ;
  assign n24484 = ~n16335 ;
  assign n16337 = n24484 & n16336 ;
  assign n24485 = ~n16332 ;
  assign n16338 = n24485 & n16337 ;
  assign n24486 = ~n16338 ;
  assign n16339 = n16331 & n24486 ;
  assign n16340 = x96 | n16339 ;
  assign n16341 = x96 & n16339 ;
  assign n24487 = ~n15797 ;
  assign n16342 = n24487 & n15798 ;
  assign n16343 = n133 & n16342 ;
  assign n16344 = n15803 & n16343 ;
  assign n16345 = n15803 | n16343 ;
  assign n24488 = ~n16344 ;
  assign n16346 = n24488 & n16345 ;
  assign n24489 = ~n16341 ;
  assign n16347 = n24489 & n16346 ;
  assign n24490 = ~n16347 ;
  assign n16348 = n16340 & n24490 ;
  assign n16349 = x97 | n16348 ;
  assign n16350 = x97 & n16348 ;
  assign n24491 = ~n15806 ;
  assign n16351 = n24491 & n15807 ;
  assign n16352 = n133 & n16351 ;
  assign n16353 = n24284 & n16352 ;
  assign n24492 = ~n16352 ;
  assign n16354 = n15812 & n24492 ;
  assign n16355 = n16353 | n16354 ;
  assign n24493 = ~n16350 ;
  assign n16356 = n24493 & n16355 ;
  assign n24494 = ~n16356 ;
  assign n16357 = n16349 & n24494 ;
  assign n16358 = x98 | n16357 ;
  assign n16359 = x98 & n16357 ;
  assign n24495 = ~n15815 ;
  assign n16360 = n24495 & n15816 ;
  assign n16361 = n133 & n16360 ;
  assign n16362 = n24287 & n16361 ;
  assign n24496 = ~n16361 ;
  assign n16363 = n15821 & n24496 ;
  assign n16364 = n16362 | n16363 ;
  assign n24497 = ~n16359 ;
  assign n16365 = n24497 & n16364 ;
  assign n24498 = ~n16365 ;
  assign n16366 = n16358 & n24498 ;
  assign n16367 = x99 | n16366 ;
  assign n16368 = x99 & n16366 ;
  assign n24499 = ~n15824 ;
  assign n16369 = n24499 & n15825 ;
  assign n16370 = n133 & n16369 ;
  assign n16371 = n15830 & n16370 ;
  assign n16372 = n15830 | n16370 ;
  assign n24500 = ~n16371 ;
  assign n16373 = n24500 & n16372 ;
  assign n24501 = ~n16368 ;
  assign n16374 = n24501 & n16373 ;
  assign n24502 = ~n16374 ;
  assign n16375 = n16367 & n24502 ;
  assign n16376 = x100 | n16375 ;
  assign n16377 = x100 & n16375 ;
  assign n24503 = ~n15833 ;
  assign n16378 = n24503 & n15834 ;
  assign n16379 = n133 & n16378 ;
  assign n16380 = n24293 & n16379 ;
  assign n24504 = ~n16379 ;
  assign n16381 = n15839 & n24504 ;
  assign n16382 = n16380 | n16381 ;
  assign n24505 = ~n16377 ;
  assign n16383 = n24505 & n16382 ;
  assign n24506 = ~n16383 ;
  assign n16384 = n16376 & n24506 ;
  assign n16385 = x101 | n16384 ;
  assign n16386 = x101 & n16384 ;
  assign n24507 = ~n15842 ;
  assign n16387 = n24507 & n15843 ;
  assign n16388 = n133 & n16387 ;
  assign n16389 = n15848 & n16388 ;
  assign n16390 = n15848 | n16388 ;
  assign n24508 = ~n16389 ;
  assign n16391 = n24508 & n16390 ;
  assign n24509 = ~n16386 ;
  assign n16392 = n24509 & n16391 ;
  assign n24510 = ~n16392 ;
  assign n16393 = n16385 & n24510 ;
  assign n16394 = x102 | n16393 ;
  assign n16395 = x102 & n16393 ;
  assign n24511 = ~n15851 ;
  assign n16396 = n24511 & n15852 ;
  assign n16397 = n133 & n16396 ;
  assign n16398 = n15857 & n16397 ;
  assign n16399 = n15857 | n16397 ;
  assign n24512 = ~n16398 ;
  assign n16400 = n24512 & n16399 ;
  assign n24513 = ~n16395 ;
  assign n16401 = n24513 & n16400 ;
  assign n24514 = ~n16401 ;
  assign n16402 = n16394 & n24514 ;
  assign n16403 = x103 | n16402 ;
  assign n16404 = x103 & n16402 ;
  assign n24515 = ~n15860 ;
  assign n16405 = n24515 & n15861 ;
  assign n16406 = n133 & n16405 ;
  assign n16407 = n15866 & n16406 ;
  assign n16408 = n15866 | n16406 ;
  assign n24516 = ~n16407 ;
  assign n16409 = n24516 & n16408 ;
  assign n24517 = ~n16404 ;
  assign n16410 = n24517 & n16409 ;
  assign n24518 = ~n16410 ;
  assign n16411 = n16403 & n24518 ;
  assign n16412 = x104 | n16411 ;
  assign n16413 = x104 & n16411 ;
  assign n24519 = ~n15869 ;
  assign n16414 = n24519 & n15870 ;
  assign n16415 = n133 & n16414 ;
  assign n16416 = n24304 & n16415 ;
  assign n24520 = ~n16415 ;
  assign n16417 = n15875 & n24520 ;
  assign n16418 = n16416 | n16417 ;
  assign n24521 = ~n16413 ;
  assign n16419 = n24521 & n16418 ;
  assign n24522 = ~n16419 ;
  assign n16420 = n16412 & n24522 ;
  assign n16421 = x105 | n16420 ;
  assign n16422 = x105 & n16420 ;
  assign n24523 = ~n15878 ;
  assign n16423 = n24523 & n15879 ;
  assign n16424 = n133 & n16423 ;
  assign n16425 = n24307 & n16424 ;
  assign n24524 = ~n16424 ;
  assign n16426 = n15884 & n24524 ;
  assign n16427 = n16425 | n16426 ;
  assign n24525 = ~n16422 ;
  assign n16428 = n24525 & n16427 ;
  assign n24526 = ~n16428 ;
  assign n16429 = n16421 & n24526 ;
  assign n16430 = x106 | n16429 ;
  assign n16431 = x106 & n16429 ;
  assign n24527 = ~n15887 ;
  assign n16432 = n24527 & n15888 ;
  assign n16433 = n133 & n16432 ;
  assign n16434 = n24310 & n16433 ;
  assign n24528 = ~n16433 ;
  assign n16435 = n15893 & n24528 ;
  assign n16436 = n16434 | n16435 ;
  assign n24529 = ~n16431 ;
  assign n16437 = n24529 & n16436 ;
  assign n24530 = ~n16437 ;
  assign n16438 = n16430 & n24530 ;
  assign n16439 = x107 | n16438 ;
  assign n16440 = x107 & n16438 ;
  assign n24531 = ~n15896 ;
  assign n16441 = n24531 & n15897 ;
  assign n16442 = n133 & n16441 ;
  assign n16443 = n24313 & n16442 ;
  assign n24532 = ~n16442 ;
  assign n16444 = n15902 & n24532 ;
  assign n16445 = n16443 | n16444 ;
  assign n24533 = ~n16440 ;
  assign n16446 = n24533 & n16445 ;
  assign n24534 = ~n16446 ;
  assign n16447 = n16439 & n24534 ;
  assign n16448 = x108 | n16447 ;
  assign n16449 = x108 & n16447 ;
  assign n24535 = ~n15905 ;
  assign n16450 = n24535 & n15906 ;
  assign n16451 = n133 & n16450 ;
  assign n16452 = n24316 & n16451 ;
  assign n24536 = ~n16451 ;
  assign n16453 = n15911 & n24536 ;
  assign n16454 = n16452 | n16453 ;
  assign n24537 = ~n16449 ;
  assign n16455 = n24537 & n16454 ;
  assign n24538 = ~n16455 ;
  assign n16456 = n16448 & n24538 ;
  assign n16457 = x109 | n16456 ;
  assign n16458 = x109 & n16456 ;
  assign n24539 = ~n15914 ;
  assign n16459 = n24539 & n15915 ;
  assign n16460 = n133 & n16459 ;
  assign n16461 = n15920 & n16460 ;
  assign n16462 = n15920 | n16460 ;
  assign n24540 = ~n16461 ;
  assign n16463 = n24540 & n16462 ;
  assign n24541 = ~n16458 ;
  assign n16464 = n24541 & n16463 ;
  assign n24542 = ~n16464 ;
  assign n16465 = n16457 & n24542 ;
  assign n16466 = x110 | n16465 ;
  assign n16467 = x110 & n16465 ;
  assign n24543 = ~n15923 ;
  assign n16468 = n24543 & n15924 ;
  assign n16469 = n133 & n16468 ;
  assign n16470 = n15929 & n16469 ;
  assign n16471 = n15929 | n16469 ;
  assign n24544 = ~n16470 ;
  assign n16472 = n24544 & n16471 ;
  assign n24545 = ~n16467 ;
  assign n16473 = n24545 & n16472 ;
  assign n24546 = ~n16473 ;
  assign n16474 = n16466 & n24546 ;
  assign n16475 = x111 | n16474 ;
  assign n16476 = x111 & n16474 ;
  assign n24547 = ~n15932 ;
  assign n16477 = n24547 & n15933 ;
  assign n16478 = n133 & n16477 ;
  assign n16479 = n15938 & n16478 ;
  assign n16480 = n15938 | n16478 ;
  assign n24548 = ~n16479 ;
  assign n16481 = n24548 & n16480 ;
  assign n24549 = ~n16476 ;
  assign n16482 = n24549 & n16481 ;
  assign n24550 = ~n16482 ;
  assign n16483 = n16475 & n24550 ;
  assign n16484 = x112 | n16483 ;
  assign n16485 = x112 & n16483 ;
  assign n24551 = ~n15941 ;
  assign n16486 = n24551 & n15942 ;
  assign n16487 = n133 & n16486 ;
  assign n16488 = n15947 & n16487 ;
  assign n16489 = n15947 | n16487 ;
  assign n24552 = ~n16488 ;
  assign n16490 = n24552 & n16489 ;
  assign n24553 = ~n16485 ;
  assign n16491 = n24553 & n16490 ;
  assign n24554 = ~n16491 ;
  assign n16492 = n16484 & n24554 ;
  assign n16493 = x113 | n16492 ;
  assign n16494 = x113 & n16492 ;
  assign n24555 = ~n15950 ;
  assign n16495 = n24555 & n15951 ;
  assign n16496 = n133 & n16495 ;
  assign n16497 = n15956 & n16496 ;
  assign n16498 = n15956 | n16496 ;
  assign n24556 = ~n16497 ;
  assign n16499 = n24556 & n16498 ;
  assign n24557 = ~n16494 ;
  assign n16500 = n24557 & n16499 ;
  assign n24558 = ~n16500 ;
  assign n16501 = n16493 & n24558 ;
  assign n16502 = x114 | n16501 ;
  assign n16503 = x114 & n16501 ;
  assign n24559 = ~n15959 ;
  assign n16504 = n24559 & n15960 ;
  assign n16505 = n133 & n16504 ;
  assign n16506 = n15965 & n16505 ;
  assign n16507 = n15965 | n16505 ;
  assign n24560 = ~n16506 ;
  assign n16508 = n24560 & n16507 ;
  assign n24561 = ~n16503 ;
  assign n16509 = n24561 & n16508 ;
  assign n24562 = ~n16509 ;
  assign n16510 = n16502 & n24562 ;
  assign n16511 = x115 | n16510 ;
  assign n16512 = x115 & n16510 ;
  assign n24563 = ~n15968 ;
  assign n16513 = n24563 & n15969 ;
  assign n16514 = n133 & n16513 ;
  assign n16515 = n15974 & n16514 ;
  assign n16516 = n15974 | n16514 ;
  assign n24564 = ~n16515 ;
  assign n16517 = n24564 & n16516 ;
  assign n24565 = ~n16512 ;
  assign n16518 = n24565 & n16517 ;
  assign n24566 = ~n16518 ;
  assign n16519 = n16511 & n24566 ;
  assign n16520 = x116 | n16519 ;
  assign n16521 = x116 & n16519 ;
  assign n24567 = ~n15977 ;
  assign n16522 = n24567 & n15978 ;
  assign n16523 = n133 & n16522 ;
  assign n16524 = n15983 & n16523 ;
  assign n16525 = n15983 | n16523 ;
  assign n24568 = ~n16524 ;
  assign n16526 = n24568 & n16525 ;
  assign n24569 = ~n16521 ;
  assign n16527 = n24569 & n16526 ;
  assign n24570 = ~n16527 ;
  assign n16528 = n16520 & n24570 ;
  assign n16529 = x117 | n16528 ;
  assign n16530 = x117 & n16528 ;
  assign n24571 = ~n15986 ;
  assign n16531 = n24571 & n15987 ;
  assign n16532 = n133 & n16531 ;
  assign n16533 = n15992 & n16532 ;
  assign n16534 = n15992 | n16532 ;
  assign n24572 = ~n16533 ;
  assign n16535 = n24572 & n16534 ;
  assign n24573 = ~n16530 ;
  assign n16536 = n24573 & n16535 ;
  assign n24574 = ~n16536 ;
  assign n16537 = n16529 & n24574 ;
  assign n16538 = x118 | n16537 ;
  assign n16539 = x118 & n16537 ;
  assign n24575 = ~n15995 ;
  assign n16540 = n24575 & n15996 ;
  assign n16541 = n133 & n16540 ;
  assign n16542 = n16001 & n16541 ;
  assign n16543 = n16001 | n16541 ;
  assign n24576 = ~n16542 ;
  assign n16544 = n24576 & n16543 ;
  assign n24577 = ~n16539 ;
  assign n16545 = n24577 & n16544 ;
  assign n24578 = ~n16545 ;
  assign n16546 = n16538 & n24578 ;
  assign n16547 = x119 | n16546 ;
  assign n16548 = x119 & n16546 ;
  assign n24579 = ~n16004 ;
  assign n16549 = n24579 & n16005 ;
  assign n16550 = n133 & n16549 ;
  assign n16551 = n16010 & n16550 ;
  assign n16552 = n16010 | n16550 ;
  assign n24580 = ~n16551 ;
  assign n16553 = n24580 & n16552 ;
  assign n24581 = ~n16548 ;
  assign n16554 = n24581 & n16553 ;
  assign n24582 = ~n16554 ;
  assign n16555 = n16547 & n24582 ;
  assign n16556 = x120 | n16555 ;
  assign n16557 = x120 & n16555 ;
  assign n24583 = ~n16013 ;
  assign n16558 = n24583 & n16014 ;
  assign n16559 = n133 & n16558 ;
  assign n16560 = n16019 & n16559 ;
  assign n16561 = n16019 | n16559 ;
  assign n24584 = ~n16560 ;
  assign n16562 = n24584 & n16561 ;
  assign n24585 = ~n16557 ;
  assign n16563 = n24585 & n16562 ;
  assign n24586 = ~n16563 ;
  assign n16564 = n16556 & n24586 ;
  assign n16565 = x121 | n16564 ;
  assign n16566 = x121 & n16564 ;
  assign n24587 = ~n16022 ;
  assign n16567 = n24587 & n16023 ;
  assign n16568 = n133 & n16567 ;
  assign n16569 = n24350 & n16568 ;
  assign n24588 = ~n16568 ;
  assign n16570 = n16028 & n24588 ;
  assign n16571 = n16569 | n16570 ;
  assign n24589 = ~n16566 ;
  assign n16572 = n24589 & n16571 ;
  assign n24590 = ~n16572 ;
  assign n16573 = n16565 & n24590 ;
  assign n16574 = x122 | n16573 ;
  assign n16575 = x122 & n16573 ;
  assign n24591 = ~n16031 ;
  assign n16576 = n24591 & n16032 ;
  assign n16577 = n133 & n16576 ;
  assign n16578 = n24353 & n16577 ;
  assign n24592 = ~n16577 ;
  assign n16579 = n16037 & n24592 ;
  assign n16580 = n16578 | n16579 ;
  assign n24593 = ~n16575 ;
  assign n16581 = n24593 & n16580 ;
  assign n24594 = ~n16581 ;
  assign n16582 = n16574 & n24594 ;
  assign n16589 = x123 & n16582 ;
  assign n24595 = ~n16589 ;
  assign n16590 = n16588 & n24595 ;
  assign n24596 = ~x124 ;
  assign n16059 = n24596 & n16057 ;
  assign n16583 = x123 | n16582 ;
  assign n24597 = ~n16059 ;
  assign n16591 = n24597 & n16583 ;
  assign n24598 = ~n16590 ;
  assign n16592 = n24598 & n16591 ;
  assign n16593 = n18273 | n16592 ;
  assign n24599 = ~n16057 ;
  assign n16595 = x124 & n24599 ;
  assign n16596 = n16593 | n16595 ;
  assign n132 = ~n16596 ;
  assign n16597 = x64 & n132 ;
  assign n16598 = x3 & n16597 ;
  assign n16599 = x3 | n16597 ;
  assign n24601 = ~n16598 ;
  assign n16600 = n24601 & n16599 ;
  assign n24602 = ~n5496 ;
  assign n16601 = n24602 & n16600 ;
  assign n24603 = ~n16601 ;
  assign n16602 = n5495 & n24603 ;
  assign n16604 = x66 | n16602 ;
  assign n16603 = x66 & n16602 ;
  assign n16605 = n24366 & n16062 ;
  assign n16606 = n132 & n16605 ;
  assign n16607 = n16067 & n16606 ;
  assign n16608 = n16067 | n16606 ;
  assign n24604 = ~n16607 ;
  assign n16609 = n24604 & n16608 ;
  assign n24605 = ~n16603 ;
  assign n16610 = n24605 & n16609 ;
  assign n24606 = ~n16610 ;
  assign n16611 = n16604 & n24606 ;
  assign n16612 = x67 | n16611 ;
  assign n16613 = x67 & n16611 ;
  assign n16614 = n16070 & n24369 ;
  assign n16615 = n132 & n16614 ;
  assign n24607 = ~n16076 ;
  assign n16616 = n24607 & n16615 ;
  assign n24608 = ~n16615 ;
  assign n16617 = n16076 & n24608 ;
  assign n16618 = n16616 | n16617 ;
  assign n24609 = ~n16613 ;
  assign n16619 = n24609 & n16618 ;
  assign n24610 = ~n16619 ;
  assign n16620 = n16612 & n24610 ;
  assign n16621 = x68 | n16620 ;
  assign n16622 = x68 & n16620 ;
  assign n16623 = n16079 & n24373 ;
  assign n16624 = n132 & n16623 ;
  assign n24611 = ~n16085 ;
  assign n16625 = n24611 & n16624 ;
  assign n24612 = ~n16624 ;
  assign n16626 = n16085 & n24612 ;
  assign n16627 = n16625 | n16626 ;
  assign n24613 = ~n16622 ;
  assign n16628 = n24613 & n16627 ;
  assign n24614 = ~n16628 ;
  assign n16629 = n16621 & n24614 ;
  assign n16630 = x69 | n16629 ;
  assign n16631 = x69 & n16629 ;
  assign n16632 = n16088 & n24377 ;
  assign n16633 = n132 & n16632 ;
  assign n24615 = ~n16094 ;
  assign n16634 = n24615 & n16633 ;
  assign n24616 = ~n16633 ;
  assign n16635 = n16094 & n24616 ;
  assign n16636 = n16634 | n16635 ;
  assign n24617 = ~n16631 ;
  assign n16637 = n24617 & n16636 ;
  assign n24618 = ~n16637 ;
  assign n16638 = n16630 & n24618 ;
  assign n16639 = x70 | n16638 ;
  assign n16640 = x70 & n16638 ;
  assign n16641 = n16097 & n24381 ;
  assign n16642 = n132 & n16641 ;
  assign n24619 = ~n16103 ;
  assign n16643 = n24619 & n16642 ;
  assign n24620 = ~n16642 ;
  assign n16644 = n16103 & n24620 ;
  assign n16645 = n16643 | n16644 ;
  assign n24621 = ~n16640 ;
  assign n16646 = n24621 & n16645 ;
  assign n24622 = ~n16646 ;
  assign n16647 = n16639 & n24622 ;
  assign n16648 = x71 | n16647 ;
  assign n16649 = x71 & n16647 ;
  assign n16650 = n16106 & n24385 ;
  assign n16651 = n132 & n16650 ;
  assign n16652 = n16112 & n16651 ;
  assign n16653 = n16112 | n16651 ;
  assign n24623 = ~n16652 ;
  assign n16654 = n24623 & n16653 ;
  assign n24624 = ~n16649 ;
  assign n16655 = n24624 & n16654 ;
  assign n24625 = ~n16655 ;
  assign n16656 = n16648 & n24625 ;
  assign n16657 = x72 | n16656 ;
  assign n16658 = x72 & n16656 ;
  assign n16659 = n16115 & n24389 ;
  assign n16660 = n132 & n16659 ;
  assign n16661 = n16121 & n16660 ;
  assign n16662 = n16121 | n16660 ;
  assign n24626 = ~n16661 ;
  assign n16663 = n24626 & n16662 ;
  assign n24627 = ~n16658 ;
  assign n16664 = n24627 & n16663 ;
  assign n24628 = ~n16664 ;
  assign n16665 = n16657 & n24628 ;
  assign n16666 = x73 | n16665 ;
  assign n16667 = x73 & n16665 ;
  assign n16668 = n16124 & n24393 ;
  assign n16669 = n132 & n16668 ;
  assign n16670 = n16130 & n16669 ;
  assign n16671 = n16130 | n16669 ;
  assign n24629 = ~n16670 ;
  assign n16672 = n24629 & n16671 ;
  assign n24630 = ~n16667 ;
  assign n16673 = n24630 & n16672 ;
  assign n24631 = ~n16673 ;
  assign n16674 = n16666 & n24631 ;
  assign n16675 = x74 | n16674 ;
  assign n16676 = x74 & n16674 ;
  assign n16677 = n16133 & n24397 ;
  assign n16678 = n132 & n16677 ;
  assign n24632 = ~n16139 ;
  assign n16679 = n24632 & n16678 ;
  assign n24633 = ~n16678 ;
  assign n16680 = n16139 & n24633 ;
  assign n16681 = n16679 | n16680 ;
  assign n24634 = ~n16676 ;
  assign n16682 = n24634 & n16681 ;
  assign n24635 = ~n16682 ;
  assign n16683 = n16675 & n24635 ;
  assign n16684 = x75 | n16683 ;
  assign n16685 = x75 & n16683 ;
  assign n16686 = n16142 & n24401 ;
  assign n16687 = n132 & n16686 ;
  assign n24636 = ~n16148 ;
  assign n16688 = n24636 & n16687 ;
  assign n24637 = ~n16687 ;
  assign n16689 = n16148 & n24637 ;
  assign n16690 = n16688 | n16689 ;
  assign n24638 = ~n16685 ;
  assign n16691 = n24638 & n16690 ;
  assign n24639 = ~n16691 ;
  assign n16692 = n16684 & n24639 ;
  assign n16693 = x76 | n16692 ;
  assign n16694 = x76 & n16692 ;
  assign n16695 = n16151 & n24405 ;
  assign n16696 = n132 & n16695 ;
  assign n24640 = ~n16157 ;
  assign n16697 = n24640 & n16696 ;
  assign n24641 = ~n16696 ;
  assign n16698 = n16157 & n24641 ;
  assign n16699 = n16697 | n16698 ;
  assign n24642 = ~n16694 ;
  assign n16700 = n24642 & n16699 ;
  assign n24643 = ~n16700 ;
  assign n16701 = n16693 & n24643 ;
  assign n16702 = x77 | n16701 ;
  assign n16703 = x77 & n16701 ;
  assign n16704 = n16160 & n24409 ;
  assign n16705 = n132 & n16704 ;
  assign n16706 = n16166 & n16705 ;
  assign n16707 = n16166 | n16705 ;
  assign n24644 = ~n16706 ;
  assign n16708 = n24644 & n16707 ;
  assign n24645 = ~n16703 ;
  assign n16709 = n24645 & n16708 ;
  assign n24646 = ~n16709 ;
  assign n16710 = n16702 & n24646 ;
  assign n16711 = x78 | n16710 ;
  assign n16712 = x78 & n16710 ;
  assign n16713 = n16169 & n24413 ;
  assign n16714 = n132 & n16713 ;
  assign n16715 = n16175 & n16714 ;
  assign n16716 = n16175 | n16714 ;
  assign n24647 = ~n16715 ;
  assign n16717 = n24647 & n16716 ;
  assign n24648 = ~n16712 ;
  assign n16718 = n24648 & n16717 ;
  assign n24649 = ~n16718 ;
  assign n16719 = n16711 & n24649 ;
  assign n16720 = x79 | n16719 ;
  assign n16721 = x79 & n16719 ;
  assign n16722 = n16178 & n24417 ;
  assign n16723 = n132 & n16722 ;
  assign n16724 = n16184 & n16723 ;
  assign n16725 = n16184 | n16723 ;
  assign n24650 = ~n16724 ;
  assign n16726 = n24650 & n16725 ;
  assign n24651 = ~n16721 ;
  assign n16727 = n24651 & n16726 ;
  assign n24652 = ~n16727 ;
  assign n16728 = n16720 & n24652 ;
  assign n16729 = x80 | n16728 ;
  assign n16730 = x80 & n16728 ;
  assign n16731 = n16187 & n24421 ;
  assign n16732 = n132 & n16731 ;
  assign n24653 = ~n16193 ;
  assign n16733 = n24653 & n16732 ;
  assign n24654 = ~n16732 ;
  assign n16734 = n16193 & n24654 ;
  assign n16735 = n16733 | n16734 ;
  assign n24655 = ~n16730 ;
  assign n16736 = n24655 & n16735 ;
  assign n24656 = ~n16736 ;
  assign n16737 = n16729 & n24656 ;
  assign n16738 = x81 | n16737 ;
  assign n16739 = x81 & n16737 ;
  assign n16740 = n16196 & n24425 ;
  assign n16741 = n132 & n16740 ;
  assign n24657 = ~n16202 ;
  assign n16742 = n24657 & n16741 ;
  assign n24658 = ~n16741 ;
  assign n16743 = n16202 & n24658 ;
  assign n16744 = n16742 | n16743 ;
  assign n24659 = ~n16739 ;
  assign n16745 = n24659 & n16744 ;
  assign n24660 = ~n16745 ;
  assign n16746 = n16738 & n24660 ;
  assign n16747 = x82 | n16746 ;
  assign n16748 = x82 & n16746 ;
  assign n16749 = n16205 & n24429 ;
  assign n16750 = n132 & n16749 ;
  assign n24661 = ~n16211 ;
  assign n16751 = n24661 & n16750 ;
  assign n24662 = ~n16750 ;
  assign n16752 = n16211 & n24662 ;
  assign n16753 = n16751 | n16752 ;
  assign n24663 = ~n16748 ;
  assign n16754 = n24663 & n16753 ;
  assign n24664 = ~n16754 ;
  assign n16755 = n16747 & n24664 ;
  assign n16756 = x83 | n16755 ;
  assign n16757 = x83 & n16755 ;
  assign n16758 = n16214 & n24433 ;
  assign n16759 = n132 & n16758 ;
  assign n16760 = n16220 & n16759 ;
  assign n16761 = n16220 | n16759 ;
  assign n24665 = ~n16760 ;
  assign n16762 = n24665 & n16761 ;
  assign n24666 = ~n16757 ;
  assign n16763 = n24666 & n16762 ;
  assign n24667 = ~n16763 ;
  assign n16764 = n16756 & n24667 ;
  assign n16765 = x84 | n16764 ;
  assign n16766 = x84 & n16764 ;
  assign n16767 = n16223 & n24437 ;
  assign n16768 = n132 & n16767 ;
  assign n24668 = ~n16229 ;
  assign n16769 = n24668 & n16768 ;
  assign n24669 = ~n16768 ;
  assign n16770 = n16229 & n24669 ;
  assign n16771 = n16769 | n16770 ;
  assign n24670 = ~n16766 ;
  assign n16772 = n24670 & n16771 ;
  assign n24671 = ~n16772 ;
  assign n16773 = n16765 & n24671 ;
  assign n16774 = x85 | n16773 ;
  assign n16775 = x85 & n16773 ;
  assign n16776 = n16232 & n24441 ;
  assign n16777 = n132 & n16776 ;
  assign n24672 = ~n16238 ;
  assign n16778 = n24672 & n16777 ;
  assign n24673 = ~n16777 ;
  assign n16779 = n16238 & n24673 ;
  assign n16780 = n16778 | n16779 ;
  assign n24674 = ~n16775 ;
  assign n16781 = n24674 & n16780 ;
  assign n24675 = ~n16781 ;
  assign n16782 = n16774 & n24675 ;
  assign n16783 = x86 | n16782 ;
  assign n16784 = x86 & n16782 ;
  assign n16785 = n16241 & n24445 ;
  assign n16786 = n132 & n16785 ;
  assign n16787 = n16247 & n16786 ;
  assign n16788 = n16247 | n16786 ;
  assign n24676 = ~n16787 ;
  assign n16789 = n24676 & n16788 ;
  assign n24677 = ~n16784 ;
  assign n16790 = n24677 & n16789 ;
  assign n24678 = ~n16790 ;
  assign n16791 = n16783 & n24678 ;
  assign n16792 = x87 | n16791 ;
  assign n16793 = x87 & n16791 ;
  assign n16794 = n16250 & n24449 ;
  assign n16795 = n132 & n16794 ;
  assign n16796 = n16256 & n16795 ;
  assign n16797 = n16256 | n16795 ;
  assign n24679 = ~n16796 ;
  assign n16798 = n24679 & n16797 ;
  assign n24680 = ~n16793 ;
  assign n16799 = n24680 & n16798 ;
  assign n24681 = ~n16799 ;
  assign n16800 = n16792 & n24681 ;
  assign n16801 = x88 | n16800 ;
  assign n16802 = x88 & n16800 ;
  assign n16803 = n16259 & n24453 ;
  assign n16804 = n132 & n16803 ;
  assign n24682 = ~n16265 ;
  assign n16805 = n24682 & n16804 ;
  assign n24683 = ~n16804 ;
  assign n16806 = n16265 & n24683 ;
  assign n16807 = n16805 | n16806 ;
  assign n24684 = ~n16802 ;
  assign n16808 = n24684 & n16807 ;
  assign n24685 = ~n16808 ;
  assign n16809 = n16801 & n24685 ;
  assign n16810 = x89 | n16809 ;
  assign n16811 = x89 & n16809 ;
  assign n16812 = n16268 & n24457 ;
  assign n16813 = n132 & n16812 ;
  assign n24686 = ~n16274 ;
  assign n16814 = n24686 & n16813 ;
  assign n24687 = ~n16813 ;
  assign n16815 = n16274 & n24687 ;
  assign n16816 = n16814 | n16815 ;
  assign n24688 = ~n16811 ;
  assign n16817 = n24688 & n16816 ;
  assign n24689 = ~n16817 ;
  assign n16818 = n16810 & n24689 ;
  assign n16819 = x90 | n16818 ;
  assign n16820 = x90 & n16818 ;
  assign n16821 = n16277 & n24461 ;
  assign n16822 = n132 & n16821 ;
  assign n24690 = ~n16283 ;
  assign n16823 = n24690 & n16822 ;
  assign n24691 = ~n16822 ;
  assign n16824 = n16283 & n24691 ;
  assign n16825 = n16823 | n16824 ;
  assign n24692 = ~n16820 ;
  assign n16826 = n24692 & n16825 ;
  assign n24693 = ~n16826 ;
  assign n16827 = n16819 & n24693 ;
  assign n16828 = x91 | n16827 ;
  assign n16829 = x91 & n16827 ;
  assign n16830 = n16286 & n24465 ;
  assign n16831 = n132 & n16830 ;
  assign n24694 = ~n16292 ;
  assign n16832 = n24694 & n16831 ;
  assign n24695 = ~n16831 ;
  assign n16833 = n16292 & n24695 ;
  assign n16834 = n16832 | n16833 ;
  assign n24696 = ~n16829 ;
  assign n16835 = n24696 & n16834 ;
  assign n24697 = ~n16835 ;
  assign n16836 = n16828 & n24697 ;
  assign n16837 = x92 | n16836 ;
  assign n16838 = x92 & n16836 ;
  assign n16839 = n16295 & n24469 ;
  assign n16840 = n132 & n16839 ;
  assign n24698 = ~n16301 ;
  assign n16841 = n24698 & n16840 ;
  assign n24699 = ~n16840 ;
  assign n16842 = n16301 & n24699 ;
  assign n16843 = n16841 | n16842 ;
  assign n24700 = ~n16838 ;
  assign n16844 = n24700 & n16843 ;
  assign n24701 = ~n16844 ;
  assign n16845 = n16837 & n24701 ;
  assign n16846 = x93 | n16845 ;
  assign n16847 = x93 & n16845 ;
  assign n16848 = n16304 & n24473 ;
  assign n16849 = n132 & n16848 ;
  assign n24702 = ~n16310 ;
  assign n16850 = n24702 & n16849 ;
  assign n24703 = ~n16849 ;
  assign n16851 = n16310 & n24703 ;
  assign n16852 = n16850 | n16851 ;
  assign n24704 = ~n16847 ;
  assign n16853 = n24704 & n16852 ;
  assign n24705 = ~n16853 ;
  assign n16854 = n16846 & n24705 ;
  assign n16855 = x94 | n16854 ;
  assign n16856 = x94 & n16854 ;
  assign n16857 = n16313 & n24477 ;
  assign n16858 = n132 & n16857 ;
  assign n16859 = n16319 & n16858 ;
  assign n16860 = n16319 | n16858 ;
  assign n24706 = ~n16859 ;
  assign n16861 = n24706 & n16860 ;
  assign n24707 = ~n16856 ;
  assign n16862 = n24707 & n16861 ;
  assign n24708 = ~n16862 ;
  assign n16863 = n16855 & n24708 ;
  assign n16864 = x95 | n16863 ;
  assign n16865 = x95 & n16863 ;
  assign n16866 = n16322 & n24481 ;
  assign n16867 = n132 & n16866 ;
  assign n24709 = ~n16328 ;
  assign n16868 = n24709 & n16867 ;
  assign n24710 = ~n16867 ;
  assign n16869 = n16328 & n24710 ;
  assign n16870 = n16868 | n16869 ;
  assign n24711 = ~n16865 ;
  assign n16871 = n24711 & n16870 ;
  assign n24712 = ~n16871 ;
  assign n16872 = n16864 & n24712 ;
  assign n16873 = x96 | n16872 ;
  assign n16874 = x96 & n16872 ;
  assign n16875 = n16331 & n24485 ;
  assign n16876 = n132 & n16875 ;
  assign n24713 = ~n16337 ;
  assign n16877 = n24713 & n16876 ;
  assign n24714 = ~n16876 ;
  assign n16878 = n16337 & n24714 ;
  assign n16879 = n16877 | n16878 ;
  assign n24715 = ~n16874 ;
  assign n16880 = n24715 & n16879 ;
  assign n24716 = ~n16880 ;
  assign n16881 = n16873 & n24716 ;
  assign n16882 = x97 | n16881 ;
  assign n16883 = x97 & n16881 ;
  assign n16884 = n16340 & n24489 ;
  assign n16885 = n132 & n16884 ;
  assign n24717 = ~n16346 ;
  assign n16886 = n24717 & n16885 ;
  assign n24718 = ~n16885 ;
  assign n16887 = n16346 & n24718 ;
  assign n16888 = n16886 | n16887 ;
  assign n24719 = ~n16883 ;
  assign n16889 = n24719 & n16888 ;
  assign n24720 = ~n16889 ;
  assign n16890 = n16882 & n24720 ;
  assign n16891 = x98 | n16890 ;
  assign n16892 = x98 & n16890 ;
  assign n16893 = n16349 & n24493 ;
  assign n16894 = n132 & n16893 ;
  assign n24721 = ~n16355 ;
  assign n16895 = n24721 & n16894 ;
  assign n24722 = ~n16894 ;
  assign n16896 = n16355 & n24722 ;
  assign n16897 = n16895 | n16896 ;
  assign n24723 = ~n16892 ;
  assign n16898 = n24723 & n16897 ;
  assign n24724 = ~n16898 ;
  assign n16899 = n16891 & n24724 ;
  assign n16900 = x99 | n16899 ;
  assign n16901 = x99 & n16899 ;
  assign n16902 = n16358 & n24497 ;
  assign n16903 = n132 & n16902 ;
  assign n24725 = ~n16364 ;
  assign n16904 = n24725 & n16903 ;
  assign n24726 = ~n16903 ;
  assign n16905 = n16364 & n24726 ;
  assign n16906 = n16904 | n16905 ;
  assign n24727 = ~n16901 ;
  assign n16907 = n24727 & n16906 ;
  assign n24728 = ~n16907 ;
  assign n16908 = n16900 & n24728 ;
  assign n16909 = x100 | n16908 ;
  assign n16910 = x100 & n16908 ;
  assign n16911 = n16367 & n24501 ;
  assign n16912 = n132 & n16911 ;
  assign n16913 = n16373 & n16912 ;
  assign n16914 = n16373 | n16912 ;
  assign n24729 = ~n16913 ;
  assign n16915 = n24729 & n16914 ;
  assign n24730 = ~n16910 ;
  assign n16916 = n24730 & n16915 ;
  assign n24731 = ~n16916 ;
  assign n16917 = n16909 & n24731 ;
  assign n16918 = x101 | n16917 ;
  assign n16919 = x101 & n16917 ;
  assign n16920 = n16376 & n24505 ;
  assign n16921 = n132 & n16920 ;
  assign n24732 = ~n16382 ;
  assign n16922 = n24732 & n16921 ;
  assign n24733 = ~n16921 ;
  assign n16923 = n16382 & n24733 ;
  assign n16924 = n16922 | n16923 ;
  assign n24734 = ~n16919 ;
  assign n16925 = n24734 & n16924 ;
  assign n24735 = ~n16925 ;
  assign n16926 = n16918 & n24735 ;
  assign n16927 = x102 | n16926 ;
  assign n16928 = x102 & n16926 ;
  assign n16929 = n16385 & n24509 ;
  assign n16930 = n132 & n16929 ;
  assign n24736 = ~n16391 ;
  assign n16931 = n24736 & n16930 ;
  assign n24737 = ~n16930 ;
  assign n16932 = n16391 & n24737 ;
  assign n16933 = n16931 | n16932 ;
  assign n24738 = ~n16928 ;
  assign n16934 = n24738 & n16933 ;
  assign n24739 = ~n16934 ;
  assign n16935 = n16927 & n24739 ;
  assign n16936 = x103 | n16935 ;
  assign n16937 = x103 & n16935 ;
  assign n16938 = n16394 & n24513 ;
  assign n16939 = n132 & n16938 ;
  assign n16940 = n16400 & n16939 ;
  assign n16941 = n16400 | n16939 ;
  assign n24740 = ~n16940 ;
  assign n16942 = n24740 & n16941 ;
  assign n24741 = ~n16937 ;
  assign n16943 = n24741 & n16942 ;
  assign n24742 = ~n16943 ;
  assign n16944 = n16936 & n24742 ;
  assign n16945 = x104 | n16944 ;
  assign n16946 = x104 & n16944 ;
  assign n16947 = n16403 & n24517 ;
  assign n16948 = n132 & n16947 ;
  assign n16949 = n16409 & n16948 ;
  assign n16950 = n16409 | n16948 ;
  assign n24743 = ~n16949 ;
  assign n16951 = n24743 & n16950 ;
  assign n24744 = ~n16946 ;
  assign n16952 = n24744 & n16951 ;
  assign n24745 = ~n16952 ;
  assign n16953 = n16945 & n24745 ;
  assign n16954 = x105 | n16953 ;
  assign n16955 = x105 & n16953 ;
  assign n16956 = n16412 & n24521 ;
  assign n16957 = n132 & n16956 ;
  assign n24746 = ~n16418 ;
  assign n16958 = n24746 & n16957 ;
  assign n24747 = ~n16957 ;
  assign n16959 = n16418 & n24747 ;
  assign n16960 = n16958 | n16959 ;
  assign n24748 = ~n16955 ;
  assign n16961 = n24748 & n16960 ;
  assign n24749 = ~n16961 ;
  assign n16962 = n16954 & n24749 ;
  assign n16963 = x106 | n16962 ;
  assign n16964 = x106 & n16962 ;
  assign n16965 = n16421 & n24525 ;
  assign n16966 = n132 & n16965 ;
  assign n24750 = ~n16427 ;
  assign n16967 = n24750 & n16966 ;
  assign n24751 = ~n16966 ;
  assign n16968 = n16427 & n24751 ;
  assign n16969 = n16967 | n16968 ;
  assign n24752 = ~n16964 ;
  assign n16970 = n24752 & n16969 ;
  assign n24753 = ~n16970 ;
  assign n16971 = n16963 & n24753 ;
  assign n16972 = x107 | n16971 ;
  assign n16973 = x107 & n16971 ;
  assign n16974 = n16430 & n24529 ;
  assign n16975 = n132 & n16974 ;
  assign n24754 = ~n16436 ;
  assign n16976 = n24754 & n16975 ;
  assign n24755 = ~n16975 ;
  assign n16977 = n16436 & n24755 ;
  assign n16978 = n16976 | n16977 ;
  assign n24756 = ~n16973 ;
  assign n16979 = n24756 & n16978 ;
  assign n24757 = ~n16979 ;
  assign n16980 = n16972 & n24757 ;
  assign n16981 = x108 | n16980 ;
  assign n16982 = x108 & n16980 ;
  assign n16983 = n16439 & n24533 ;
  assign n16984 = n132 & n16983 ;
  assign n24758 = ~n16445 ;
  assign n16985 = n24758 & n16984 ;
  assign n24759 = ~n16984 ;
  assign n16986 = n16445 & n24759 ;
  assign n16987 = n16985 | n16986 ;
  assign n24760 = ~n16982 ;
  assign n16988 = n24760 & n16987 ;
  assign n24761 = ~n16988 ;
  assign n16989 = n16981 & n24761 ;
  assign n16990 = x109 | n16989 ;
  assign n16991 = x109 & n16989 ;
  assign n16992 = n16448 & n24537 ;
  assign n16993 = n132 & n16992 ;
  assign n24762 = ~n16454 ;
  assign n16994 = n24762 & n16993 ;
  assign n24763 = ~n16993 ;
  assign n16995 = n16454 & n24763 ;
  assign n16996 = n16994 | n16995 ;
  assign n24764 = ~n16991 ;
  assign n16997 = n24764 & n16996 ;
  assign n24765 = ~n16997 ;
  assign n16998 = n16990 & n24765 ;
  assign n16999 = x110 | n16998 ;
  assign n17000 = x110 & n16998 ;
  assign n17001 = n16457 & n24541 ;
  assign n17002 = n132 & n17001 ;
  assign n17003 = n16463 & n17002 ;
  assign n17004 = n16463 | n17002 ;
  assign n24766 = ~n17003 ;
  assign n17005 = n24766 & n17004 ;
  assign n24767 = ~n17000 ;
  assign n17006 = n24767 & n17005 ;
  assign n24768 = ~n17006 ;
  assign n17007 = n16999 & n24768 ;
  assign n17008 = x111 | n17007 ;
  assign n17009 = x111 & n17007 ;
  assign n17010 = n16466 & n24545 ;
  assign n17011 = n132 & n17010 ;
  assign n17012 = n16472 & n17011 ;
  assign n17013 = n16472 | n17011 ;
  assign n24769 = ~n17012 ;
  assign n17014 = n24769 & n17013 ;
  assign n24770 = ~n17009 ;
  assign n17015 = n24770 & n17014 ;
  assign n24771 = ~n17015 ;
  assign n17016 = n17008 & n24771 ;
  assign n17017 = x112 | n17016 ;
  assign n17018 = x112 & n17016 ;
  assign n17019 = n16475 & n24549 ;
  assign n17020 = n132 & n17019 ;
  assign n24772 = ~n16481 ;
  assign n17021 = n24772 & n17020 ;
  assign n24773 = ~n17020 ;
  assign n17022 = n16481 & n24773 ;
  assign n17023 = n17021 | n17022 ;
  assign n24774 = ~n17018 ;
  assign n17024 = n24774 & n17023 ;
  assign n24775 = ~n17024 ;
  assign n17025 = n17017 & n24775 ;
  assign n17026 = x113 | n17025 ;
  assign n17027 = x113 & n17025 ;
  assign n17028 = n16484 & n24553 ;
  assign n17029 = n132 & n17028 ;
  assign n24776 = ~n16490 ;
  assign n17030 = n24776 & n17029 ;
  assign n24777 = ~n17029 ;
  assign n17031 = n16490 & n24777 ;
  assign n17032 = n17030 | n17031 ;
  assign n24778 = ~n17027 ;
  assign n17033 = n24778 & n17032 ;
  assign n24779 = ~n17033 ;
  assign n17034 = n17026 & n24779 ;
  assign n17035 = x114 | n17034 ;
  assign n17036 = x114 & n17034 ;
  assign n17037 = n16493 & n24557 ;
  assign n17038 = n132 & n17037 ;
  assign n17039 = n16499 & n17038 ;
  assign n17040 = n16499 | n17038 ;
  assign n24780 = ~n17039 ;
  assign n17041 = n24780 & n17040 ;
  assign n24781 = ~n17036 ;
  assign n17042 = n24781 & n17041 ;
  assign n24782 = ~n17042 ;
  assign n17043 = n17035 & n24782 ;
  assign n17044 = x115 | n17043 ;
  assign n17045 = x115 & n17043 ;
  assign n17046 = n16502 & n24561 ;
  assign n17047 = n132 & n17046 ;
  assign n17048 = n16508 & n17047 ;
  assign n17049 = n16508 | n17047 ;
  assign n24783 = ~n17048 ;
  assign n17050 = n24783 & n17049 ;
  assign n24784 = ~n17045 ;
  assign n17051 = n24784 & n17050 ;
  assign n24785 = ~n17051 ;
  assign n17052 = n17044 & n24785 ;
  assign n17053 = x116 | n17052 ;
  assign n17054 = x116 & n17052 ;
  assign n17055 = n16511 & n24565 ;
  assign n17056 = n132 & n17055 ;
  assign n17057 = n16517 & n17056 ;
  assign n17058 = n16517 | n17056 ;
  assign n24786 = ~n17057 ;
  assign n17059 = n24786 & n17058 ;
  assign n24787 = ~n17054 ;
  assign n17060 = n24787 & n17059 ;
  assign n24788 = ~n17060 ;
  assign n17061 = n17053 & n24788 ;
  assign n17062 = x117 | n17061 ;
  assign n17063 = x117 & n17061 ;
  assign n17064 = n16520 & n24569 ;
  assign n17065 = n132 & n17064 ;
  assign n17066 = n16526 & n17065 ;
  assign n17067 = n16526 | n17065 ;
  assign n24789 = ~n17066 ;
  assign n17068 = n24789 & n17067 ;
  assign n24790 = ~n17063 ;
  assign n17069 = n24790 & n17068 ;
  assign n24791 = ~n17069 ;
  assign n17070 = n17062 & n24791 ;
  assign n17071 = x118 | n17070 ;
  assign n17072 = x118 & n17070 ;
  assign n17073 = n16529 & n24573 ;
  assign n17074 = n132 & n17073 ;
  assign n17075 = n16535 & n17074 ;
  assign n17076 = n16535 | n17074 ;
  assign n24792 = ~n17075 ;
  assign n17077 = n24792 & n17076 ;
  assign n24793 = ~n17072 ;
  assign n17078 = n24793 & n17077 ;
  assign n24794 = ~n17078 ;
  assign n17079 = n17071 & n24794 ;
  assign n17080 = x119 | n17079 ;
  assign n17081 = x119 & n17079 ;
  assign n17082 = n16538 & n24577 ;
  assign n17083 = n132 & n17082 ;
  assign n17084 = n16544 & n17083 ;
  assign n17085 = n16544 | n17083 ;
  assign n24795 = ~n17084 ;
  assign n17086 = n24795 & n17085 ;
  assign n24796 = ~n17081 ;
  assign n17087 = n24796 & n17086 ;
  assign n24797 = ~n17087 ;
  assign n17088 = n17080 & n24797 ;
  assign n17089 = x120 | n17088 ;
  assign n17090 = x120 & n17088 ;
  assign n17091 = n16547 & n24581 ;
  assign n17092 = n132 & n17091 ;
  assign n24798 = ~n16553 ;
  assign n17093 = n24798 & n17092 ;
  assign n24799 = ~n17092 ;
  assign n17094 = n16553 & n24799 ;
  assign n17095 = n17093 | n17094 ;
  assign n24800 = ~n17090 ;
  assign n17096 = n24800 & n17095 ;
  assign n24801 = ~n17096 ;
  assign n17097 = n17089 & n24801 ;
  assign n17098 = x121 | n17097 ;
  assign n17099 = x121 & n17097 ;
  assign n17100 = n16556 & n24585 ;
  assign n17101 = n132 & n17100 ;
  assign n24802 = ~n16562 ;
  assign n17102 = n24802 & n17101 ;
  assign n24803 = ~n17101 ;
  assign n17103 = n16562 & n24803 ;
  assign n17104 = n17102 | n17103 ;
  assign n24804 = ~n17099 ;
  assign n17105 = n24804 & n17104 ;
  assign n24805 = ~n17105 ;
  assign n17106 = n17098 & n24805 ;
  assign n17107 = x122 | n17106 ;
  assign n17108 = x122 & n17106 ;
  assign n17109 = n16565 & n24589 ;
  assign n17110 = n132 & n17109 ;
  assign n24806 = ~n16571 ;
  assign n17111 = n24806 & n17110 ;
  assign n24807 = ~n17110 ;
  assign n17112 = n16571 & n24807 ;
  assign n17113 = n17111 | n17112 ;
  assign n24808 = ~n17108 ;
  assign n17114 = n24808 & n17113 ;
  assign n24809 = ~n17114 ;
  assign n17115 = n17107 & n24809 ;
  assign n17116 = x123 | n17115 ;
  assign n17117 = x123 & n17115 ;
  assign n17118 = n16574 & n24593 ;
  assign n17119 = n132 & n17118 ;
  assign n24810 = ~n16580 ;
  assign n17120 = n24810 & n17119 ;
  assign n24811 = ~n17119 ;
  assign n17121 = n16580 & n24811 ;
  assign n17122 = n17120 | n17121 ;
  assign n24812 = ~n17117 ;
  assign n17123 = n24812 & n17122 ;
  assign n24813 = ~n17123 ;
  assign n17124 = n17116 & n24813 ;
  assign n17126 = x124 | n17124 ;
  assign n17127 = n16583 & n24595 ;
  assign n17128 = n132 & n17127 ;
  assign n17129 = n16588 & n17128 ;
  assign n17130 = n16588 | n17128 ;
  assign n24814 = ~n17129 ;
  assign n17131 = n24814 & n17130 ;
  assign n24815 = ~n17131 ;
  assign n17132 = n17126 & n24815 ;
  assign n16594 = n21884 | n16593 ;
  assign n17133 = n16057 & n16594 ;
  assign n24816 = ~n18268 ;
  assign n17134 = x125 & n24816 ;
  assign n24817 = ~n17134 ;
  assign n17135 = n17133 & n24817 ;
  assign n17136 = x124 & n17124 ;
  assign n17137 = n17135 | n17136 ;
  assign n17138 = n17132 | n17137 ;
  assign n17139 = n16058 & n17138 ;
  assign n17140 = n21884 | n17139 ;
  assign n24818 = ~x0 ;
  assign n5489 = n24818 & x64 ;
  assign n5490 = x65 | n5489 ;
  assign n5491 = x65 & n5489 ;
  assign n24819 = ~x1 ;
  assign n5492 = n24819 & x64 ;
  assign n17141 = x65 | n5492 ;
  assign n5493 = x65 & n5492 ;
  assign n24820 = ~n18273 ;
  assign n17142 = n24820 & n17133 ;
  assign n17143 = n18273 & n24599 ;
  assign n17144 = n17138 | n17143 ;
  assign n24821 = ~n17142 ;
  assign n17145 = n24821 & n17144 ;
  assign n131 = ~n17145 ;
  assign n17146 = x64 & n131 ;
  assign n17147 = x2 & n17146 ;
  assign n17148 = x2 | n17146 ;
  assign n24823 = ~n17147 ;
  assign n17149 = n24823 & n17148 ;
  assign n24824 = ~n5493 ;
  assign n17150 = n24824 & n17149 ;
  assign n24825 = ~n17150 ;
  assign n17151 = n17141 & n24825 ;
  assign n17152 = x66 | n17151 ;
  assign n17153 = x66 & n17151 ;
  assign n17154 = n5495 & n24602 ;
  assign n17155 = n131 & n17154 ;
  assign n17156 = n16600 & n17155 ;
  assign n17157 = n16600 | n17155 ;
  assign n24826 = ~n17156 ;
  assign n17158 = n24826 & n17157 ;
  assign n24827 = ~n17153 ;
  assign n17159 = n24827 & n17158 ;
  assign n24828 = ~n17159 ;
  assign n17160 = n17152 & n24828 ;
  assign n17162 = x67 & n17160 ;
  assign n17161 = x67 | n17160 ;
  assign n17163 = n16604 & n131 ;
  assign n17164 = n16610 & n17163 ;
  assign n17165 = n24605 & n17163 ;
  assign n17166 = n16609 | n17165 ;
  assign n24829 = ~n17164 ;
  assign n17167 = n24829 & n17166 ;
  assign n24830 = ~n17167 ;
  assign n17168 = n17161 & n24830 ;
  assign n17169 = n17162 | n17168 ;
  assign n17170 = x68 & n17169 ;
  assign n17171 = x68 | n17169 ;
  assign n17172 = n16612 & n131 ;
  assign n17173 = n16619 & n17172 ;
  assign n17174 = n24609 & n17172 ;
  assign n17175 = n16618 | n17174 ;
  assign n24831 = ~n17173 ;
  assign n17176 = n24831 & n17175 ;
  assign n24832 = ~n17176 ;
  assign n17177 = n17171 & n24832 ;
  assign n17178 = n17170 | n17177 ;
  assign n17179 = x69 & n17178 ;
  assign n17180 = x69 | n17178 ;
  assign n17181 = n16621 & n24613 ;
  assign n17182 = n131 & n17181 ;
  assign n24833 = ~n16627 ;
  assign n17183 = n24833 & n17182 ;
  assign n24834 = ~n17182 ;
  assign n17184 = n16627 & n24834 ;
  assign n17185 = n17183 | n17184 ;
  assign n24835 = ~n17185 ;
  assign n17186 = n17180 & n24835 ;
  assign n17187 = n17179 | n17186 ;
  assign n17188 = x70 & n17187 ;
  assign n17189 = x70 | n17187 ;
  assign n17190 = n16630 & n24617 ;
  assign n17191 = n131 & n17190 ;
  assign n24836 = ~n16636 ;
  assign n17192 = n24836 & n17191 ;
  assign n24837 = ~n17191 ;
  assign n17193 = n16636 & n24837 ;
  assign n17194 = n17192 | n17193 ;
  assign n24838 = ~n17194 ;
  assign n17195 = n17189 & n24838 ;
  assign n17196 = n17188 | n17195 ;
  assign n17197 = x71 & n17196 ;
  assign n17198 = x71 | n17196 ;
  assign n17199 = n16639 & n24621 ;
  assign n17200 = n131 & n17199 ;
  assign n17201 = n16645 & n17200 ;
  assign n17202 = n16645 | n17200 ;
  assign n24839 = ~n17201 ;
  assign n17203 = n24839 & n17202 ;
  assign n24840 = ~n17203 ;
  assign n17204 = n17198 & n24840 ;
  assign n17205 = n17197 | n17204 ;
  assign n17206 = x72 & n17205 ;
  assign n17207 = x72 | n17205 ;
  assign n17208 = n16648 & n24624 ;
  assign n17209 = n131 & n17208 ;
  assign n17210 = n16654 & n17209 ;
  assign n17211 = n16654 | n17209 ;
  assign n24841 = ~n17210 ;
  assign n17212 = n24841 & n17211 ;
  assign n24842 = ~n17212 ;
  assign n17213 = n17207 & n24842 ;
  assign n17214 = n17206 | n17213 ;
  assign n17215 = x73 & n17214 ;
  assign n17216 = x73 | n17214 ;
  assign n17217 = n16657 & n24627 ;
  assign n17218 = n131 & n17217 ;
  assign n24843 = ~n16663 ;
  assign n17219 = n24843 & n17218 ;
  assign n24844 = ~n17218 ;
  assign n17220 = n16663 & n24844 ;
  assign n17221 = n17219 | n17220 ;
  assign n24845 = ~n17221 ;
  assign n17222 = n17216 & n24845 ;
  assign n17223 = n17215 | n17222 ;
  assign n17224 = x74 & n17223 ;
  assign n17225 = x74 | n17223 ;
  assign n17226 = n16666 & n24630 ;
  assign n17227 = n131 & n17226 ;
  assign n17228 = n16672 & n17227 ;
  assign n17229 = n16672 | n17227 ;
  assign n24846 = ~n17228 ;
  assign n17230 = n24846 & n17229 ;
  assign n24847 = ~n17230 ;
  assign n17231 = n17225 & n24847 ;
  assign n17232 = n17224 | n17231 ;
  assign n17233 = x75 & n17232 ;
  assign n17234 = x75 | n17232 ;
  assign n17235 = n16675 & n24634 ;
  assign n17236 = n131 & n17235 ;
  assign n24848 = ~n16681 ;
  assign n17237 = n24848 & n17236 ;
  assign n24849 = ~n17236 ;
  assign n17238 = n16681 & n24849 ;
  assign n17239 = n17237 | n17238 ;
  assign n24850 = ~n17239 ;
  assign n17240 = n17234 & n24850 ;
  assign n17241 = n17233 | n17240 ;
  assign n17242 = x76 & n17241 ;
  assign n17243 = x76 | n17241 ;
  assign n17244 = n16684 & n24638 ;
  assign n17245 = n131 & n17244 ;
  assign n17246 = n16690 & n17245 ;
  assign n17247 = n16690 | n17245 ;
  assign n24851 = ~n17246 ;
  assign n17248 = n24851 & n17247 ;
  assign n24852 = ~n17248 ;
  assign n17249 = n17243 & n24852 ;
  assign n17250 = n17242 | n17249 ;
  assign n17251 = x77 & n17250 ;
  assign n17252 = x77 | n17250 ;
  assign n17253 = n16693 & n24642 ;
  assign n17254 = n131 & n17253 ;
  assign n24853 = ~n16699 ;
  assign n17255 = n24853 & n17254 ;
  assign n24854 = ~n17254 ;
  assign n17256 = n16699 & n24854 ;
  assign n17257 = n17255 | n17256 ;
  assign n24855 = ~n17257 ;
  assign n17258 = n17252 & n24855 ;
  assign n17259 = n17251 | n17258 ;
  assign n17260 = x78 & n17259 ;
  assign n17261 = x78 | n17259 ;
  assign n17262 = n16702 & n24645 ;
  assign n17263 = n131 & n17262 ;
  assign n24856 = ~n16708 ;
  assign n17264 = n24856 & n17263 ;
  assign n24857 = ~n17263 ;
  assign n17265 = n16708 & n24857 ;
  assign n17266 = n17264 | n17265 ;
  assign n24858 = ~n17266 ;
  assign n17267 = n17261 & n24858 ;
  assign n17268 = n17260 | n17267 ;
  assign n17269 = x79 & n17268 ;
  assign n17270 = x79 | n17268 ;
  assign n17271 = n16711 & n24648 ;
  assign n17272 = n131 & n17271 ;
  assign n17273 = n16717 & n17272 ;
  assign n17274 = n16717 | n17272 ;
  assign n24859 = ~n17273 ;
  assign n17275 = n24859 & n17274 ;
  assign n24860 = ~n17275 ;
  assign n17276 = n17270 & n24860 ;
  assign n17277 = n17269 | n17276 ;
  assign n17278 = x80 & n17277 ;
  assign n17279 = x80 | n17277 ;
  assign n17280 = n16720 & n24651 ;
  assign n17281 = n131 & n17280 ;
  assign n17282 = n16726 & n17281 ;
  assign n17283 = n16726 | n17281 ;
  assign n24861 = ~n17282 ;
  assign n17284 = n24861 & n17283 ;
  assign n24862 = ~n17284 ;
  assign n17285 = n17279 & n24862 ;
  assign n17286 = n17278 | n17285 ;
  assign n17287 = x81 & n17286 ;
  assign n17288 = x81 | n17286 ;
  assign n17289 = n16729 & n24655 ;
  assign n17290 = n131 & n17289 ;
  assign n24863 = ~n16735 ;
  assign n17291 = n24863 & n17290 ;
  assign n24864 = ~n17290 ;
  assign n17292 = n16735 & n24864 ;
  assign n17293 = n17291 | n17292 ;
  assign n24865 = ~n17293 ;
  assign n17294 = n17288 & n24865 ;
  assign n17295 = n17287 | n17294 ;
  assign n17296 = x82 & n17295 ;
  assign n17297 = x82 | n17295 ;
  assign n17298 = n16738 & n24659 ;
  assign n17299 = n131 & n17298 ;
  assign n24866 = ~n16744 ;
  assign n17300 = n24866 & n17299 ;
  assign n24867 = ~n17299 ;
  assign n17301 = n16744 & n24867 ;
  assign n17302 = n17300 | n17301 ;
  assign n24868 = ~n17302 ;
  assign n17303 = n17297 & n24868 ;
  assign n17304 = n17296 | n17303 ;
  assign n17305 = x83 & n17304 ;
  assign n17306 = x83 | n17304 ;
  assign n17307 = n16747 & n24663 ;
  assign n17308 = n131 & n17307 ;
  assign n17309 = n16753 & n17308 ;
  assign n17310 = n16753 | n17308 ;
  assign n24869 = ~n17309 ;
  assign n17311 = n24869 & n17310 ;
  assign n24870 = ~n17311 ;
  assign n17312 = n17306 & n24870 ;
  assign n17313 = n17305 | n17312 ;
  assign n17314 = x84 & n17313 ;
  assign n17315 = x84 | n17313 ;
  assign n17316 = n16756 & n24666 ;
  assign n17317 = n131 & n17316 ;
  assign n24871 = ~n16762 ;
  assign n17318 = n24871 & n17317 ;
  assign n24872 = ~n17317 ;
  assign n17319 = n16762 & n24872 ;
  assign n17320 = n17318 | n17319 ;
  assign n24873 = ~n17320 ;
  assign n17321 = n17315 & n24873 ;
  assign n17322 = n17314 | n17321 ;
  assign n17323 = x85 & n17322 ;
  assign n17324 = x85 | n17322 ;
  assign n17325 = n16765 & n24670 ;
  assign n17326 = n131 & n17325 ;
  assign n17327 = n16771 & n17326 ;
  assign n17328 = n16771 | n17326 ;
  assign n24874 = ~n17327 ;
  assign n17329 = n24874 & n17328 ;
  assign n24875 = ~n17329 ;
  assign n17330 = n17324 & n24875 ;
  assign n17331 = n17323 | n17330 ;
  assign n17332 = x86 & n17331 ;
  assign n17333 = x86 | n17331 ;
  assign n17334 = n16774 & n24674 ;
  assign n17335 = n131 & n17334 ;
  assign n24876 = ~n16780 ;
  assign n17336 = n24876 & n17335 ;
  assign n24877 = ~n17335 ;
  assign n17337 = n16780 & n24877 ;
  assign n17338 = n17336 | n17337 ;
  assign n24878 = ~n17338 ;
  assign n17339 = n17333 & n24878 ;
  assign n17340 = n17332 | n17339 ;
  assign n17341 = x87 & n17340 ;
  assign n17342 = x87 | n17340 ;
  assign n17343 = n16783 & n24677 ;
  assign n17344 = n131 & n17343 ;
  assign n24879 = ~n16789 ;
  assign n17345 = n24879 & n17344 ;
  assign n24880 = ~n17344 ;
  assign n17346 = n16789 & n24880 ;
  assign n17347 = n17345 | n17346 ;
  assign n24881 = ~n17347 ;
  assign n17348 = n17342 & n24881 ;
  assign n17349 = n17341 | n17348 ;
  assign n17350 = x88 & n17349 ;
  assign n17351 = x88 | n17349 ;
  assign n17352 = n16792 & n24680 ;
  assign n17353 = n131 & n17352 ;
  assign n17354 = n16798 & n17353 ;
  assign n17355 = n16798 | n17353 ;
  assign n24882 = ~n17354 ;
  assign n17356 = n24882 & n17355 ;
  assign n24883 = ~n17356 ;
  assign n17357 = n17351 & n24883 ;
  assign n17358 = n17350 | n17357 ;
  assign n17359 = x89 & n17358 ;
  assign n17360 = x89 | n17358 ;
  assign n17361 = n16801 & n24684 ;
  assign n17362 = n131 & n17361 ;
  assign n24884 = ~n16807 ;
  assign n17363 = n24884 & n17362 ;
  assign n24885 = ~n17362 ;
  assign n17364 = n16807 & n24885 ;
  assign n17365 = n17363 | n17364 ;
  assign n24886 = ~n17365 ;
  assign n17366 = n17360 & n24886 ;
  assign n17367 = n17359 | n17366 ;
  assign n17368 = x90 & n17367 ;
  assign n17369 = x90 | n17367 ;
  assign n17370 = n16810 & n24688 ;
  assign n17371 = n131 & n17370 ;
  assign n24887 = ~n16816 ;
  assign n17372 = n24887 & n17371 ;
  assign n24888 = ~n17371 ;
  assign n17373 = n16816 & n24888 ;
  assign n17374 = n17372 | n17373 ;
  assign n24889 = ~n17374 ;
  assign n17375 = n17369 & n24889 ;
  assign n17376 = n17368 | n17375 ;
  assign n17377 = x91 & n17376 ;
  assign n17378 = x91 | n17376 ;
  assign n17379 = n16819 & n24692 ;
  assign n17380 = n131 & n17379 ;
  assign n24890 = ~n16825 ;
  assign n17381 = n24890 & n17380 ;
  assign n24891 = ~n17380 ;
  assign n17382 = n16825 & n24891 ;
  assign n17383 = n17381 | n17382 ;
  assign n24892 = ~n17383 ;
  assign n17384 = n17378 & n24892 ;
  assign n17385 = n17377 | n17384 ;
  assign n17386 = x92 & n17385 ;
  assign n17387 = x92 | n17385 ;
  assign n17388 = n16828 & n24696 ;
  assign n17389 = n131 & n17388 ;
  assign n24893 = ~n16834 ;
  assign n17390 = n24893 & n17389 ;
  assign n24894 = ~n17389 ;
  assign n17391 = n16834 & n24894 ;
  assign n17392 = n17390 | n17391 ;
  assign n24895 = ~n17392 ;
  assign n17393 = n17387 & n24895 ;
  assign n17394 = n17386 | n17393 ;
  assign n17395 = x93 & n17394 ;
  assign n17396 = x93 | n17394 ;
  assign n17397 = n16837 & n24700 ;
  assign n17398 = n131 & n17397 ;
  assign n24896 = ~n16843 ;
  assign n17399 = n24896 & n17398 ;
  assign n24897 = ~n17398 ;
  assign n17400 = n16843 & n24897 ;
  assign n17401 = n17399 | n17400 ;
  assign n24898 = ~n17401 ;
  assign n17402 = n17396 & n24898 ;
  assign n17403 = n17395 | n17402 ;
  assign n17404 = x94 & n17403 ;
  assign n17405 = x94 | n17403 ;
  assign n17406 = n16846 & n24704 ;
  assign n17407 = n131 & n17406 ;
  assign n24899 = ~n16852 ;
  assign n17408 = n24899 & n17407 ;
  assign n24900 = ~n17407 ;
  assign n17409 = n16852 & n24900 ;
  assign n17410 = n17408 | n17409 ;
  assign n24901 = ~n17410 ;
  assign n17411 = n17405 & n24901 ;
  assign n17412 = n17404 | n17411 ;
  assign n17413 = x95 & n17412 ;
  assign n17414 = x95 | n17412 ;
  assign n17415 = n16855 & n24707 ;
  assign n17416 = n131 & n17415 ;
  assign n17417 = n16861 & n17416 ;
  assign n17418 = n16861 | n17416 ;
  assign n24902 = ~n17417 ;
  assign n17419 = n24902 & n17418 ;
  assign n24903 = ~n17419 ;
  assign n17420 = n17414 & n24903 ;
  assign n17421 = n17413 | n17420 ;
  assign n17422 = x96 & n17421 ;
  assign n17423 = x96 | n17421 ;
  assign n17424 = n16864 & n24711 ;
  assign n17425 = n131 & n17424 ;
  assign n24904 = ~n16870 ;
  assign n17426 = n24904 & n17425 ;
  assign n24905 = ~n17425 ;
  assign n17427 = n16870 & n24905 ;
  assign n17428 = n17426 | n17427 ;
  assign n24906 = ~n17428 ;
  assign n17429 = n17423 & n24906 ;
  assign n17430 = n17422 | n17429 ;
  assign n17431 = x97 & n17430 ;
  assign n17432 = x97 | n17430 ;
  assign n17433 = n16873 & n24715 ;
  assign n17434 = n131 & n17433 ;
  assign n24907 = ~n16879 ;
  assign n17435 = n24907 & n17434 ;
  assign n24908 = ~n17434 ;
  assign n17436 = n16879 & n24908 ;
  assign n17437 = n17435 | n17436 ;
  assign n24909 = ~n17437 ;
  assign n17438 = n17432 & n24909 ;
  assign n17439 = n17431 | n17438 ;
  assign n17440 = x98 & n17439 ;
  assign n17441 = x98 | n17439 ;
  assign n17442 = n16882 & n24719 ;
  assign n17443 = n131 & n17442 ;
  assign n24910 = ~n16888 ;
  assign n17444 = n24910 & n17443 ;
  assign n24911 = ~n17443 ;
  assign n17445 = n16888 & n24911 ;
  assign n17446 = n17444 | n17445 ;
  assign n24912 = ~n17446 ;
  assign n17447 = n17441 & n24912 ;
  assign n17448 = n17440 | n17447 ;
  assign n17449 = x99 & n17448 ;
  assign n17450 = x99 | n17448 ;
  assign n17451 = n16891 & n24723 ;
  assign n17452 = n131 & n17451 ;
  assign n24913 = ~n16897 ;
  assign n17453 = n24913 & n17452 ;
  assign n24914 = ~n17452 ;
  assign n17454 = n16897 & n24914 ;
  assign n17455 = n17453 | n17454 ;
  assign n24915 = ~n17455 ;
  assign n17456 = n17450 & n24915 ;
  assign n17457 = n17449 | n17456 ;
  assign n17458 = x100 & n17457 ;
  assign n17459 = x100 | n17457 ;
  assign n17460 = n16900 & n24727 ;
  assign n17461 = n131 & n17460 ;
  assign n24916 = ~n16906 ;
  assign n17462 = n24916 & n17461 ;
  assign n24917 = ~n17461 ;
  assign n17463 = n16906 & n24917 ;
  assign n17464 = n17462 | n17463 ;
  assign n24918 = ~n17464 ;
  assign n17465 = n17459 & n24918 ;
  assign n17466 = n17458 | n17465 ;
  assign n17467 = x101 & n17466 ;
  assign n17468 = x101 | n17466 ;
  assign n17469 = n16909 & n24730 ;
  assign n17470 = n131 & n17469 ;
  assign n24919 = ~n16915 ;
  assign n17471 = n24919 & n17470 ;
  assign n24920 = ~n17470 ;
  assign n17472 = n16915 & n24920 ;
  assign n17473 = n17471 | n17472 ;
  assign n24921 = ~n17473 ;
  assign n17474 = n17468 & n24921 ;
  assign n17475 = n17467 | n17474 ;
  assign n17476 = x102 & n17475 ;
  assign n17477 = x102 | n17475 ;
  assign n17478 = n16918 & n24734 ;
  assign n17479 = n131 & n17478 ;
  assign n24922 = ~n16924 ;
  assign n17480 = n24922 & n17479 ;
  assign n24923 = ~n17479 ;
  assign n17481 = n16924 & n24923 ;
  assign n17482 = n17480 | n17481 ;
  assign n24924 = ~n17482 ;
  assign n17483 = n17477 & n24924 ;
  assign n17484 = n17476 | n17483 ;
  assign n17485 = x103 & n17484 ;
  assign n17486 = x103 | n17484 ;
  assign n17487 = n16927 & n24738 ;
  assign n17488 = n131 & n17487 ;
  assign n24925 = ~n16933 ;
  assign n17489 = n24925 & n17488 ;
  assign n24926 = ~n17488 ;
  assign n17490 = n16933 & n24926 ;
  assign n17491 = n17489 | n17490 ;
  assign n24927 = ~n17491 ;
  assign n17492 = n17486 & n24927 ;
  assign n17493 = n17485 | n17492 ;
  assign n17494 = x104 & n17493 ;
  assign n17495 = x104 | n17493 ;
  assign n17496 = n16936 & n24741 ;
  assign n17497 = n131 & n17496 ;
  assign n17498 = n16942 & n17497 ;
  assign n17499 = n16942 | n17497 ;
  assign n24928 = ~n17498 ;
  assign n17500 = n24928 & n17499 ;
  assign n24929 = ~n17500 ;
  assign n17501 = n17495 & n24929 ;
  assign n17502 = n17494 | n17501 ;
  assign n17503 = x105 & n17502 ;
  assign n17504 = x105 | n17502 ;
  assign n17505 = n16945 & n24744 ;
  assign n17506 = n131 & n17505 ;
  assign n24930 = ~n16951 ;
  assign n17507 = n24930 & n17506 ;
  assign n24931 = ~n17506 ;
  assign n17508 = n16951 & n24931 ;
  assign n17509 = n17507 | n17508 ;
  assign n24932 = ~n17509 ;
  assign n17510 = n17504 & n24932 ;
  assign n17511 = n17503 | n17510 ;
  assign n17512 = x106 & n17511 ;
  assign n17513 = x106 | n17511 ;
  assign n17514 = n16954 & n24748 ;
  assign n17515 = n131 & n17514 ;
  assign n24933 = ~n16960 ;
  assign n17516 = n24933 & n17515 ;
  assign n24934 = ~n17515 ;
  assign n17517 = n16960 & n24934 ;
  assign n17518 = n17516 | n17517 ;
  assign n24935 = ~n17518 ;
  assign n17519 = n17513 & n24935 ;
  assign n17520 = n17512 | n17519 ;
  assign n17521 = x107 & n17520 ;
  assign n17522 = x107 | n17520 ;
  assign n17523 = n16963 & n24752 ;
  assign n17524 = n131 & n17523 ;
  assign n24936 = ~n16969 ;
  assign n17525 = n24936 & n17524 ;
  assign n24937 = ~n17524 ;
  assign n17526 = n16969 & n24937 ;
  assign n17527 = n17525 | n17526 ;
  assign n24938 = ~n17527 ;
  assign n17528 = n17522 & n24938 ;
  assign n17529 = n17521 | n17528 ;
  assign n17530 = x108 & n17529 ;
  assign n17531 = x108 | n17529 ;
  assign n17532 = n16972 & n24756 ;
  assign n17533 = n131 & n17532 ;
  assign n24939 = ~n16978 ;
  assign n17534 = n24939 & n17533 ;
  assign n24940 = ~n17533 ;
  assign n17535 = n16978 & n24940 ;
  assign n17536 = n17534 | n17535 ;
  assign n24941 = ~n17536 ;
  assign n17537 = n17531 & n24941 ;
  assign n17538 = n17530 | n17537 ;
  assign n17539 = x109 & n17538 ;
  assign n17540 = x109 | n17538 ;
  assign n17541 = n16981 & n24760 ;
  assign n17542 = n131 & n17541 ;
  assign n24942 = ~n16987 ;
  assign n17543 = n24942 & n17542 ;
  assign n24943 = ~n17542 ;
  assign n17544 = n16987 & n24943 ;
  assign n17545 = n17543 | n17544 ;
  assign n24944 = ~n17545 ;
  assign n17546 = n17540 & n24944 ;
  assign n17547 = n17539 | n17546 ;
  assign n17548 = x110 & n17547 ;
  assign n17549 = x110 | n17547 ;
  assign n17550 = n16990 & n24764 ;
  assign n17551 = n131 & n17550 ;
  assign n17552 = n16996 & n17551 ;
  assign n17553 = n16996 | n17551 ;
  assign n24945 = ~n17552 ;
  assign n17554 = n24945 & n17553 ;
  assign n24946 = ~n17554 ;
  assign n17555 = n17549 & n24946 ;
  assign n17556 = n17548 | n17555 ;
  assign n17557 = x111 & n17556 ;
  assign n17558 = x111 | n17556 ;
  assign n17559 = n16999 & n24767 ;
  assign n17560 = n131 & n17559 ;
  assign n24947 = ~n17005 ;
  assign n17561 = n24947 & n17560 ;
  assign n24948 = ~n17560 ;
  assign n17562 = n17005 & n24948 ;
  assign n17563 = n17561 | n17562 ;
  assign n24949 = ~n17563 ;
  assign n17564 = n17558 & n24949 ;
  assign n17565 = n17557 | n17564 ;
  assign n17566 = x112 & n17565 ;
  assign n17567 = x112 | n17565 ;
  assign n17568 = n17008 & n24770 ;
  assign n17569 = n131 & n17568 ;
  assign n24950 = ~n17014 ;
  assign n17570 = n24950 & n17569 ;
  assign n24951 = ~n17569 ;
  assign n17571 = n17014 & n24951 ;
  assign n17572 = n17570 | n17571 ;
  assign n24952 = ~n17572 ;
  assign n17573 = n17567 & n24952 ;
  assign n17574 = n17566 | n17573 ;
  assign n17575 = x113 & n17574 ;
  assign n17576 = x113 | n17574 ;
  assign n17577 = n17017 & n24774 ;
  assign n17578 = n131 & n17577 ;
  assign n24953 = ~n17023 ;
  assign n17579 = n24953 & n17578 ;
  assign n24954 = ~n17578 ;
  assign n17580 = n17023 & n24954 ;
  assign n17581 = n17579 | n17580 ;
  assign n24955 = ~n17581 ;
  assign n17582 = n17576 & n24955 ;
  assign n17583 = n17575 | n17582 ;
  assign n17584 = x114 & n17583 ;
  assign n17585 = x114 | n17583 ;
  assign n17586 = n17026 & n24778 ;
  assign n17587 = n131 & n17586 ;
  assign n24956 = ~n17032 ;
  assign n17588 = n24956 & n17587 ;
  assign n24957 = ~n17587 ;
  assign n17589 = n17032 & n24957 ;
  assign n17590 = n17588 | n17589 ;
  assign n24958 = ~n17590 ;
  assign n17591 = n17585 & n24958 ;
  assign n17592 = n17584 | n17591 ;
  assign n17593 = x115 & n17592 ;
  assign n17594 = x115 | n17592 ;
  assign n17595 = n17035 & n24781 ;
  assign n17596 = n131 & n17595 ;
  assign n17597 = n17041 & n17596 ;
  assign n17598 = n17041 | n17596 ;
  assign n24959 = ~n17597 ;
  assign n17599 = n24959 & n17598 ;
  assign n24960 = ~n17599 ;
  assign n17600 = n17594 & n24960 ;
  assign n17601 = n17593 | n17600 ;
  assign n17602 = x116 & n17601 ;
  assign n17603 = x116 | n17601 ;
  assign n17604 = n17044 & n24784 ;
  assign n17605 = n131 & n17604 ;
  assign n17606 = n17050 & n17605 ;
  assign n17607 = n17050 | n17605 ;
  assign n24961 = ~n17606 ;
  assign n17608 = n24961 & n17607 ;
  assign n24962 = ~n17608 ;
  assign n17609 = n17603 & n24962 ;
  assign n17610 = n17602 | n17609 ;
  assign n17611 = x117 & n17610 ;
  assign n17612 = x117 | n17610 ;
  assign n17613 = n17053 & n24787 ;
  assign n17614 = n131 & n17613 ;
  assign n24963 = ~n17059 ;
  assign n17615 = n24963 & n17614 ;
  assign n24964 = ~n17614 ;
  assign n17616 = n17059 & n24964 ;
  assign n17617 = n17615 | n17616 ;
  assign n24965 = ~n17617 ;
  assign n17618 = n17612 & n24965 ;
  assign n17619 = n17611 | n17618 ;
  assign n17620 = x118 & n17619 ;
  assign n17621 = x118 | n17619 ;
  assign n17622 = n17062 & n24790 ;
  assign n17623 = n131 & n17622 ;
  assign n17624 = n17068 & n17623 ;
  assign n17625 = n17068 | n17623 ;
  assign n24966 = ~n17624 ;
  assign n17626 = n24966 & n17625 ;
  assign n24967 = ~n17626 ;
  assign n17627 = n17621 & n24967 ;
  assign n17628 = n17620 | n17627 ;
  assign n17629 = x119 & n17628 ;
  assign n17630 = x119 | n17628 ;
  assign n17631 = n17071 & n24793 ;
  assign n17632 = n131 & n17631 ;
  assign n24968 = ~n17077 ;
  assign n17633 = n24968 & n17632 ;
  assign n24969 = ~n17632 ;
  assign n17634 = n17077 & n24969 ;
  assign n17635 = n17633 | n17634 ;
  assign n24970 = ~n17635 ;
  assign n17636 = n17630 & n24970 ;
  assign n17637 = n17629 | n17636 ;
  assign n17638 = x120 & n17637 ;
  assign n17639 = x120 | n17637 ;
  assign n17640 = n17080 & n24796 ;
  assign n17641 = n131 & n17640 ;
  assign n17642 = n17086 & n17641 ;
  assign n17643 = n17086 | n17641 ;
  assign n24971 = ~n17642 ;
  assign n17644 = n24971 & n17643 ;
  assign n24972 = ~n17644 ;
  assign n17645 = n17639 & n24972 ;
  assign n17646 = n17638 | n17645 ;
  assign n17647 = x121 & n17646 ;
  assign n17648 = x121 | n17646 ;
  assign n17649 = n17089 & n24800 ;
  assign n17650 = n131 & n17649 ;
  assign n24973 = ~n17095 ;
  assign n17651 = n24973 & n17650 ;
  assign n24974 = ~n17650 ;
  assign n17652 = n17095 & n24974 ;
  assign n17653 = n17651 | n17652 ;
  assign n24975 = ~n17653 ;
  assign n17654 = n17648 & n24975 ;
  assign n17655 = n17647 | n17654 ;
  assign n17656 = x122 & n17655 ;
  assign n17657 = x122 | n17655 ;
  assign n17658 = n17098 & n24804 ;
  assign n17659 = n131 & n17658 ;
  assign n24976 = ~n17104 ;
  assign n17660 = n24976 & n17659 ;
  assign n24977 = ~n17659 ;
  assign n17661 = n17104 & n24977 ;
  assign n17662 = n17660 | n17661 ;
  assign n24978 = ~n17662 ;
  assign n17663 = n17657 & n24978 ;
  assign n17664 = n17656 | n17663 ;
  assign n17665 = x123 & n17664 ;
  assign n17666 = x123 | n17664 ;
  assign n17667 = n17107 & n24808 ;
  assign n17668 = n131 & n17667 ;
  assign n24979 = ~n17113 ;
  assign n17669 = n24979 & n17668 ;
  assign n24980 = ~n17668 ;
  assign n17670 = n17113 & n24980 ;
  assign n17671 = n17669 | n17670 ;
  assign n24981 = ~n17671 ;
  assign n17672 = n17666 & n24981 ;
  assign n17673 = n17665 | n17672 ;
  assign n17674 = x124 & n17673 ;
  assign n17675 = x124 | n17673 ;
  assign n17676 = n17116 & n24812 ;
  assign n17677 = n131 & n17676 ;
  assign n24982 = ~n17122 ;
  assign n17678 = n24982 & n17677 ;
  assign n24983 = ~n17677 ;
  assign n17679 = n17122 & n24983 ;
  assign n17680 = n17678 | n17679 ;
  assign n24984 = ~n17680 ;
  assign n17681 = n17675 & n24984 ;
  assign n17682 = n17674 | n17681 ;
  assign n17683 = x125 & n17682 ;
  assign n17684 = x125 | n17682 ;
  assign n17125 = n24596 & n17124 ;
  assign n24985 = ~n17124 ;
  assign n17685 = x124 & n24985 ;
  assign n17686 = n17125 | n17685 ;
  assign n17687 = n131 & n17686 ;
  assign n17688 = n17131 & n17687 ;
  assign n17689 = n17131 | n17687 ;
  assign n24986 = ~n17688 ;
  assign n17690 = n24986 & n17689 ;
  assign n24987 = ~n17690 ;
  assign n17691 = n17684 & n24987 ;
  assign n17692 = n17683 | n17691 ;
  assign n17693 = x126 | n17692 ;
  assign n24988 = ~n17140 ;
  assign n17694 = n24988 & n17693 ;
  assign n17695 = x126 & n17692 ;
  assign n17696 = x127 | n17695 ;
  assign n17697 = n17694 | n17696 ;
  assign n130 = ~n17697 ;
  assign n17699 = n5492 & n130 ;
  assign n17698 = x64 & n130 ;
  assign n24990 = ~n17698 ;
  assign n17700 = x1 & n24990 ;
  assign n17701 = n17699 | n17700 ;
  assign n24991 = ~n5491 ;
  assign n17702 = n24991 & n17701 ;
  assign n24992 = ~n17702 ;
  assign n17703 = n5490 & n24992 ;
  assign n17704 = x66 | n17703 ;
  assign n17705 = n24824 & n17141 ;
  assign n17706 = n130 & n17705 ;
  assign n17707 = n17149 & n17706 ;
  assign n17708 = n17149 | n17706 ;
  assign n24993 = ~n17707 ;
  assign n17709 = n24993 & n17708 ;
  assign n17710 = x66 & n17703 ;
  assign n24994 = ~n17710 ;
  assign n17711 = n17709 & n24994 ;
  assign n24995 = ~n17711 ;
  assign n17712 = n17704 & n24995 ;
  assign n17713 = x67 | n17712 ;
  assign n17714 = n17152 & n24827 ;
  assign n17715 = n130 & n17714 ;
  assign n17716 = n17158 | n17715 ;
  assign n17717 = n17158 & n17715 ;
  assign n24996 = ~n17717 ;
  assign n17718 = n17716 & n24996 ;
  assign n17719 = x67 & n17712 ;
  assign n24997 = ~n17719 ;
  assign n17720 = n17718 & n24997 ;
  assign n24998 = ~n17720 ;
  assign n17721 = n17713 & n24998 ;
  assign n17722 = x68 | n17721 ;
  assign n17723 = x68 & n17721 ;
  assign n17724 = n17162 | n17697 ;
  assign n24999 = ~n17724 ;
  assign n17725 = n17168 & n24999 ;
  assign n17726 = n17161 & n24999 ;
  assign n25000 = ~n17726 ;
  assign n17727 = n17167 & n25000 ;
  assign n17728 = n17725 | n17727 ;
  assign n25001 = ~n17723 ;
  assign n17729 = n25001 & n17728 ;
  assign n25002 = ~n17729 ;
  assign n17730 = n17722 & n25002 ;
  assign n17731 = x69 | n17730 ;
  assign n17732 = x69 & n17730 ;
  assign n25003 = ~n17170 ;
  assign n17733 = n25003 & n17171 ;
  assign n17734 = n130 & n17733 ;
  assign n17735 = n17176 & n17734 ;
  assign n17736 = n17176 | n17734 ;
  assign n25004 = ~n17735 ;
  assign n17737 = n25004 & n17736 ;
  assign n25005 = ~n17732 ;
  assign n17738 = n25005 & n17737 ;
  assign n25006 = ~n17738 ;
  assign n17739 = n17731 & n25006 ;
  assign n17740 = x70 | n17739 ;
  assign n17741 = x70 & n17739 ;
  assign n25007 = ~n17179 ;
  assign n17742 = n25007 & n17180 ;
  assign n17743 = n130 & n17742 ;
  assign n17744 = n17185 & n17743 ;
  assign n17745 = n17185 | n17743 ;
  assign n25008 = ~n17744 ;
  assign n17746 = n25008 & n17745 ;
  assign n25009 = ~n17741 ;
  assign n17747 = n25009 & n17746 ;
  assign n25010 = ~n17747 ;
  assign n17748 = n17740 & n25010 ;
  assign n17749 = x71 | n17748 ;
  assign n17750 = x71 & n17748 ;
  assign n25011 = ~n17188 ;
  assign n17751 = n25011 & n17189 ;
  assign n17752 = n130 & n17751 ;
  assign n17753 = n24838 & n17752 ;
  assign n25012 = ~n17752 ;
  assign n17754 = n17194 & n25012 ;
  assign n17755 = n17753 | n17754 ;
  assign n25013 = ~n17750 ;
  assign n17756 = n25013 & n17755 ;
  assign n25014 = ~n17756 ;
  assign n17757 = n17749 & n25014 ;
  assign n17758 = x72 | n17757 ;
  assign n17759 = x72 & n17757 ;
  assign n25015 = ~n17197 ;
  assign n17760 = n25015 & n17198 ;
  assign n17761 = n130 & n17760 ;
  assign n17762 = n17203 & n17761 ;
  assign n17763 = n17203 | n17761 ;
  assign n25016 = ~n17762 ;
  assign n17764 = n25016 & n17763 ;
  assign n25017 = ~n17759 ;
  assign n17765 = n25017 & n17764 ;
  assign n25018 = ~n17765 ;
  assign n17766 = n17758 & n25018 ;
  assign n17767 = x73 | n17766 ;
  assign n17768 = x73 & n17766 ;
  assign n25019 = ~n17206 ;
  assign n17769 = n25019 & n17207 ;
  assign n17770 = n130 & n17769 ;
  assign n17771 = n17212 & n17770 ;
  assign n17772 = n17212 | n17770 ;
  assign n25020 = ~n17771 ;
  assign n17773 = n25020 & n17772 ;
  assign n25021 = ~n17768 ;
  assign n17774 = n25021 & n17773 ;
  assign n25022 = ~n17774 ;
  assign n17775 = n17767 & n25022 ;
  assign n17776 = x74 | n17775 ;
  assign n17777 = x74 & n17775 ;
  assign n25023 = ~n17215 ;
  assign n17778 = n25023 & n17216 ;
  assign n17779 = n130 & n17778 ;
  assign n17780 = n24845 & n17779 ;
  assign n25024 = ~n17779 ;
  assign n17781 = n17221 & n25024 ;
  assign n17782 = n17780 | n17781 ;
  assign n25025 = ~n17777 ;
  assign n17783 = n25025 & n17782 ;
  assign n25026 = ~n17783 ;
  assign n17784 = n17776 & n25026 ;
  assign n17785 = x75 | n17784 ;
  assign n17786 = x75 & n17784 ;
  assign n25027 = ~n17224 ;
  assign n17787 = n25027 & n17225 ;
  assign n17788 = n130 & n17787 ;
  assign n17789 = n17230 & n17788 ;
  assign n17790 = n17230 | n17788 ;
  assign n25028 = ~n17789 ;
  assign n17791 = n25028 & n17790 ;
  assign n25029 = ~n17786 ;
  assign n17792 = n25029 & n17791 ;
  assign n25030 = ~n17792 ;
  assign n17793 = n17785 & n25030 ;
  assign n17794 = x76 | n17793 ;
  assign n17795 = x76 & n17793 ;
  assign n25031 = ~n17233 ;
  assign n17796 = n25031 & n17234 ;
  assign n17797 = n130 & n17796 ;
  assign n17798 = n17239 & n17797 ;
  assign n17799 = n17239 | n17797 ;
  assign n25032 = ~n17798 ;
  assign n17800 = n25032 & n17799 ;
  assign n25033 = ~n17795 ;
  assign n17801 = n25033 & n17800 ;
  assign n25034 = ~n17801 ;
  assign n17802 = n17794 & n25034 ;
  assign n17803 = x77 | n17802 ;
  assign n17804 = x77 & n17802 ;
  assign n25035 = ~n17242 ;
  assign n17805 = n25035 & n17243 ;
  assign n17806 = n130 & n17805 ;
  assign n17807 = n17248 & n17806 ;
  assign n17808 = n17248 | n17806 ;
  assign n25036 = ~n17807 ;
  assign n17809 = n25036 & n17808 ;
  assign n25037 = ~n17804 ;
  assign n17810 = n25037 & n17809 ;
  assign n25038 = ~n17810 ;
  assign n17811 = n17803 & n25038 ;
  assign n17812 = x78 | n17811 ;
  assign n17813 = x78 & n17811 ;
  assign n25039 = ~n17251 ;
  assign n17814 = n25039 & n17252 ;
  assign n17815 = n130 & n17814 ;
  assign n17816 = n17257 & n17815 ;
  assign n17817 = n17257 | n17815 ;
  assign n25040 = ~n17816 ;
  assign n17818 = n25040 & n17817 ;
  assign n25041 = ~n17813 ;
  assign n17819 = n25041 & n17818 ;
  assign n25042 = ~n17819 ;
  assign n17820 = n17812 & n25042 ;
  assign n17821 = x79 | n17820 ;
  assign n17822 = x79 & n17820 ;
  assign n25043 = ~n17260 ;
  assign n17823 = n25043 & n17261 ;
  assign n17824 = n130 & n17823 ;
  assign n17825 = n24858 & n17824 ;
  assign n25044 = ~n17824 ;
  assign n17826 = n17266 & n25044 ;
  assign n17827 = n17825 | n17826 ;
  assign n25045 = ~n17822 ;
  assign n17828 = n25045 & n17827 ;
  assign n25046 = ~n17828 ;
  assign n17829 = n17821 & n25046 ;
  assign n17830 = x80 | n17829 ;
  assign n17831 = x80 & n17829 ;
  assign n25047 = ~n17269 ;
  assign n17832 = n25047 & n17270 ;
  assign n17833 = n130 & n17832 ;
  assign n17834 = n17275 & n17833 ;
  assign n17835 = n17275 | n17833 ;
  assign n25048 = ~n17834 ;
  assign n17836 = n25048 & n17835 ;
  assign n25049 = ~n17831 ;
  assign n17837 = n25049 & n17836 ;
  assign n25050 = ~n17837 ;
  assign n17838 = n17830 & n25050 ;
  assign n17839 = x81 | n17838 ;
  assign n17840 = x81 & n17838 ;
  assign n25051 = ~n17278 ;
  assign n17841 = n25051 & n17279 ;
  assign n17842 = n130 & n17841 ;
  assign n17843 = n17284 & n17842 ;
  assign n17844 = n17284 | n17842 ;
  assign n25052 = ~n17843 ;
  assign n17845 = n25052 & n17844 ;
  assign n25053 = ~n17840 ;
  assign n17846 = n25053 & n17845 ;
  assign n25054 = ~n17846 ;
  assign n17847 = n17839 & n25054 ;
  assign n17848 = x82 | n17847 ;
  assign n17849 = x82 & n17847 ;
  assign n25055 = ~n17287 ;
  assign n17850 = n25055 & n17288 ;
  assign n17851 = n130 & n17850 ;
  assign n17852 = n24865 & n17851 ;
  assign n25056 = ~n17851 ;
  assign n17853 = n17293 & n25056 ;
  assign n17854 = n17852 | n17853 ;
  assign n25057 = ~n17849 ;
  assign n17855 = n25057 & n17854 ;
  assign n25058 = ~n17855 ;
  assign n17856 = n17848 & n25058 ;
  assign n17857 = x83 | n17856 ;
  assign n17858 = x83 & n17856 ;
  assign n25059 = ~n17296 ;
  assign n17859 = n25059 & n17297 ;
  assign n17860 = n130 & n17859 ;
  assign n17861 = n17302 & n17860 ;
  assign n17862 = n17302 | n17860 ;
  assign n25060 = ~n17861 ;
  assign n17863 = n25060 & n17862 ;
  assign n25061 = ~n17858 ;
  assign n17864 = n25061 & n17863 ;
  assign n25062 = ~n17864 ;
  assign n17865 = n17857 & n25062 ;
  assign n17866 = x84 | n17865 ;
  assign n17867 = x84 & n17865 ;
  assign n25063 = ~n17305 ;
  assign n17868 = n25063 & n17306 ;
  assign n17869 = n130 & n17868 ;
  assign n17870 = n17311 & n17869 ;
  assign n17871 = n17311 | n17869 ;
  assign n25064 = ~n17870 ;
  assign n17872 = n25064 & n17871 ;
  assign n25065 = ~n17867 ;
  assign n17873 = n25065 & n17872 ;
  assign n25066 = ~n17873 ;
  assign n17874 = n17866 & n25066 ;
  assign n17875 = x85 | n17874 ;
  assign n17876 = x85 & n17874 ;
  assign n25067 = ~n17314 ;
  assign n17877 = n25067 & n17315 ;
  assign n17878 = n130 & n17877 ;
  assign n17879 = n24873 & n17878 ;
  assign n25068 = ~n17878 ;
  assign n17880 = n17320 & n25068 ;
  assign n17881 = n17879 | n17880 ;
  assign n25069 = ~n17876 ;
  assign n17882 = n25069 & n17881 ;
  assign n25070 = ~n17882 ;
  assign n17883 = n17875 & n25070 ;
  assign n17884 = x86 | n17883 ;
  assign n17885 = x86 & n17883 ;
  assign n25071 = ~n17323 ;
  assign n17886 = n25071 & n17324 ;
  assign n17887 = n130 & n17886 ;
  assign n17888 = n17329 & n17887 ;
  assign n17889 = n17329 | n17887 ;
  assign n25072 = ~n17888 ;
  assign n17890 = n25072 & n17889 ;
  assign n25073 = ~n17885 ;
  assign n17891 = n25073 & n17890 ;
  assign n25074 = ~n17891 ;
  assign n17892 = n17884 & n25074 ;
  assign n17893 = x87 | n17892 ;
  assign n17894 = x87 & n17892 ;
  assign n25075 = ~n17332 ;
  assign n17895 = n25075 & n17333 ;
  assign n17896 = n130 & n17895 ;
  assign n17897 = n24878 & n17896 ;
  assign n25076 = ~n17896 ;
  assign n17898 = n17338 & n25076 ;
  assign n17899 = n17897 | n17898 ;
  assign n25077 = ~n17894 ;
  assign n17900 = n25077 & n17899 ;
  assign n25078 = ~n17900 ;
  assign n17901 = n17893 & n25078 ;
  assign n17902 = x88 | n17901 ;
  assign n17903 = x88 & n17901 ;
  assign n25079 = ~n17341 ;
  assign n17904 = n25079 & n17342 ;
  assign n17905 = n130 & n17904 ;
  assign n17906 = n24881 & n17905 ;
  assign n25080 = ~n17905 ;
  assign n17907 = n17347 & n25080 ;
  assign n17908 = n17906 | n17907 ;
  assign n25081 = ~n17903 ;
  assign n17909 = n25081 & n17908 ;
  assign n25082 = ~n17909 ;
  assign n17910 = n17902 & n25082 ;
  assign n17911 = x89 | n17910 ;
  assign n17912 = x89 & n17910 ;
  assign n25083 = ~n17350 ;
  assign n17913 = n25083 & n17351 ;
  assign n17914 = n130 & n17913 ;
  assign n17915 = n17356 & n17914 ;
  assign n17916 = n17356 | n17914 ;
  assign n25084 = ~n17915 ;
  assign n17917 = n25084 & n17916 ;
  assign n25085 = ~n17912 ;
  assign n17918 = n25085 & n17917 ;
  assign n25086 = ~n17918 ;
  assign n17919 = n17911 & n25086 ;
  assign n17920 = x90 | n17919 ;
  assign n17921 = x90 & n17919 ;
  assign n25087 = ~n17359 ;
  assign n17922 = n25087 & n17360 ;
  assign n17923 = n130 & n17922 ;
  assign n17924 = n17365 & n17923 ;
  assign n17925 = n17365 | n17923 ;
  assign n25088 = ~n17924 ;
  assign n17926 = n25088 & n17925 ;
  assign n25089 = ~n17921 ;
  assign n17927 = n25089 & n17926 ;
  assign n25090 = ~n17927 ;
  assign n17928 = n17920 & n25090 ;
  assign n17929 = x91 | n17928 ;
  assign n17930 = x91 & n17928 ;
  assign n25091 = ~n17368 ;
  assign n17931 = n25091 & n17369 ;
  assign n17932 = n130 & n17931 ;
  assign n17933 = n24889 & n17932 ;
  assign n25092 = ~n17932 ;
  assign n17934 = n17374 & n25092 ;
  assign n17935 = n17933 | n17934 ;
  assign n25093 = ~n17930 ;
  assign n17936 = n25093 & n17935 ;
  assign n25094 = ~n17936 ;
  assign n17937 = n17929 & n25094 ;
  assign n17938 = x92 | n17937 ;
  assign n17939 = x92 & n17937 ;
  assign n25095 = ~n17377 ;
  assign n17940 = n25095 & n17378 ;
  assign n17941 = n130 & n17940 ;
  assign n17942 = n24892 & n17941 ;
  assign n25096 = ~n17941 ;
  assign n17943 = n17383 & n25096 ;
  assign n17944 = n17942 | n17943 ;
  assign n25097 = ~n17939 ;
  assign n17945 = n25097 & n17944 ;
  assign n25098 = ~n17945 ;
  assign n17946 = n17938 & n25098 ;
  assign n17947 = x93 | n17946 ;
  assign n17948 = x93 & n17946 ;
  assign n25099 = ~n17386 ;
  assign n17949 = n25099 & n17387 ;
  assign n17950 = n130 & n17949 ;
  assign n17951 = n17392 & n17950 ;
  assign n17952 = n17392 | n17950 ;
  assign n25100 = ~n17951 ;
  assign n17953 = n25100 & n17952 ;
  assign n25101 = ~n17948 ;
  assign n17954 = n25101 & n17953 ;
  assign n25102 = ~n17954 ;
  assign n17955 = n17947 & n25102 ;
  assign n17956 = x94 | n17955 ;
  assign n17957 = x94 & n17955 ;
  assign n25103 = ~n17395 ;
  assign n17958 = n25103 & n17396 ;
  assign n17959 = n130 & n17958 ;
  assign n17960 = n24898 & n17959 ;
  assign n25104 = ~n17959 ;
  assign n17961 = n17401 & n25104 ;
  assign n17962 = n17960 | n17961 ;
  assign n25105 = ~n17957 ;
  assign n17963 = n25105 & n17962 ;
  assign n25106 = ~n17963 ;
  assign n17964 = n17956 & n25106 ;
  assign n17965 = x95 | n17964 ;
  assign n17966 = x95 & n17964 ;
  assign n25107 = ~n17404 ;
  assign n17967 = n25107 & n17405 ;
  assign n17968 = n130 & n17967 ;
  assign n17969 = n24901 & n17968 ;
  assign n25108 = ~n17968 ;
  assign n17970 = n17410 & n25108 ;
  assign n17971 = n17969 | n17970 ;
  assign n25109 = ~n17966 ;
  assign n17972 = n25109 & n17971 ;
  assign n25110 = ~n17972 ;
  assign n17973 = n17965 & n25110 ;
  assign n17974 = x96 | n17973 ;
  assign n17975 = x96 & n17973 ;
  assign n25111 = ~n17413 ;
  assign n17976 = n25111 & n17414 ;
  assign n17977 = n130 & n17976 ;
  assign n17978 = n17419 & n17977 ;
  assign n17979 = n17419 | n17977 ;
  assign n25112 = ~n17978 ;
  assign n17980 = n25112 & n17979 ;
  assign n25113 = ~n17975 ;
  assign n17981 = n25113 & n17980 ;
  assign n25114 = ~n17981 ;
  assign n17982 = n17974 & n25114 ;
  assign n17983 = x97 | n17982 ;
  assign n17984 = x97 & n17982 ;
  assign n25115 = ~n17422 ;
  assign n17985 = n25115 & n17423 ;
  assign n17986 = n130 & n17985 ;
  assign n17987 = n24906 & n17986 ;
  assign n25116 = ~n17986 ;
  assign n17988 = n17428 & n25116 ;
  assign n17989 = n17987 | n17988 ;
  assign n25117 = ~n17984 ;
  assign n17990 = n25117 & n17989 ;
  assign n25118 = ~n17990 ;
  assign n17991 = n17983 & n25118 ;
  assign n17992 = x98 | n17991 ;
  assign n17993 = x98 & n17991 ;
  assign n25119 = ~n17431 ;
  assign n17994 = n25119 & n17432 ;
  assign n17995 = n130 & n17994 ;
  assign n17996 = n17437 & n17995 ;
  assign n17997 = n17437 | n17995 ;
  assign n25120 = ~n17996 ;
  assign n17998 = n25120 & n17997 ;
  assign n25121 = ~n17993 ;
  assign n17999 = n25121 & n17998 ;
  assign n25122 = ~n17999 ;
  assign n18000 = n17992 & n25122 ;
  assign n18001 = x99 | n18000 ;
  assign n18002 = x99 & n18000 ;
  assign n25123 = ~n17440 ;
  assign n18003 = n25123 & n17441 ;
  assign n18004 = n130 & n18003 ;
  assign n18005 = n24912 & n18004 ;
  assign n25124 = ~n18004 ;
  assign n18006 = n17446 & n25124 ;
  assign n18007 = n18005 | n18006 ;
  assign n25125 = ~n18002 ;
  assign n18008 = n25125 & n18007 ;
  assign n25126 = ~n18008 ;
  assign n18009 = n18001 & n25126 ;
  assign n18010 = x100 | n18009 ;
  assign n18011 = x100 & n18009 ;
  assign n25127 = ~n17449 ;
  assign n18012 = n25127 & n17450 ;
  assign n18013 = n130 & n18012 ;
  assign n18014 = n24915 & n18013 ;
  assign n25128 = ~n18013 ;
  assign n18015 = n17455 & n25128 ;
  assign n18016 = n18014 | n18015 ;
  assign n25129 = ~n18011 ;
  assign n18017 = n25129 & n18016 ;
  assign n25130 = ~n18017 ;
  assign n18018 = n18010 & n25130 ;
  assign n18019 = x101 | n18018 ;
  assign n18020 = x101 & n18018 ;
  assign n25131 = ~n17458 ;
  assign n18021 = n25131 & n17459 ;
  assign n18022 = n130 & n18021 ;
  assign n18023 = n17464 & n18022 ;
  assign n18024 = n17464 | n18022 ;
  assign n25132 = ~n18023 ;
  assign n18025 = n25132 & n18024 ;
  assign n25133 = ~n18020 ;
  assign n18026 = n25133 & n18025 ;
  assign n25134 = ~n18026 ;
  assign n18027 = n18019 & n25134 ;
  assign n18028 = x102 | n18027 ;
  assign n18029 = x102 & n18027 ;
  assign n25135 = ~n17467 ;
  assign n18030 = n25135 & n17468 ;
  assign n18031 = n130 & n18030 ;
  assign n18032 = n24921 & n18031 ;
  assign n25136 = ~n18031 ;
  assign n18033 = n17473 & n25136 ;
  assign n18034 = n18032 | n18033 ;
  assign n25137 = ~n18029 ;
  assign n18035 = n25137 & n18034 ;
  assign n25138 = ~n18035 ;
  assign n18036 = n18028 & n25138 ;
  assign n18037 = x103 | n18036 ;
  assign n18038 = x103 & n18036 ;
  assign n25139 = ~n17476 ;
  assign n18039 = n25139 & n17477 ;
  assign n18040 = n130 & n18039 ;
  assign n18041 = n24924 & n18040 ;
  assign n25140 = ~n18040 ;
  assign n18042 = n17482 & n25140 ;
  assign n18043 = n18041 | n18042 ;
  assign n25141 = ~n18038 ;
  assign n18044 = n25141 & n18043 ;
  assign n25142 = ~n18044 ;
  assign n18045 = n18037 & n25142 ;
  assign n18046 = x104 | n18045 ;
  assign n18047 = x104 & n18045 ;
  assign n25143 = ~n17485 ;
  assign n18048 = n25143 & n17486 ;
  assign n18049 = n130 & n18048 ;
  assign n18050 = n24927 & n18049 ;
  assign n25144 = ~n18049 ;
  assign n18051 = n17491 & n25144 ;
  assign n18052 = n18050 | n18051 ;
  assign n25145 = ~n18047 ;
  assign n18053 = n25145 & n18052 ;
  assign n25146 = ~n18053 ;
  assign n18054 = n18046 & n25146 ;
  assign n18055 = x105 | n18054 ;
  assign n18056 = x105 & n18054 ;
  assign n25147 = ~n17494 ;
  assign n18057 = n25147 & n17495 ;
  assign n18058 = n130 & n18057 ;
  assign n18059 = n17500 & n18058 ;
  assign n18060 = n17500 | n18058 ;
  assign n25148 = ~n18059 ;
  assign n18061 = n25148 & n18060 ;
  assign n25149 = ~n18056 ;
  assign n18062 = n25149 & n18061 ;
  assign n25150 = ~n18062 ;
  assign n18063 = n18055 & n25150 ;
  assign n18064 = x106 | n18063 ;
  assign n18065 = x106 & n18063 ;
  assign n25151 = ~n17503 ;
  assign n18066 = n25151 & n17504 ;
  assign n18067 = n130 & n18066 ;
  assign n18068 = n24932 & n18067 ;
  assign n25152 = ~n18067 ;
  assign n18069 = n17509 & n25152 ;
  assign n18070 = n18068 | n18069 ;
  assign n25153 = ~n18065 ;
  assign n18071 = n25153 & n18070 ;
  assign n25154 = ~n18071 ;
  assign n18072 = n18064 & n25154 ;
  assign n18073 = x107 | n18072 ;
  assign n18074 = x107 & n18072 ;
  assign n25155 = ~n17512 ;
  assign n18075 = n25155 & n17513 ;
  assign n18076 = n130 & n18075 ;
  assign n18077 = n17518 & n18076 ;
  assign n18078 = n17518 | n18076 ;
  assign n25156 = ~n18077 ;
  assign n18079 = n25156 & n18078 ;
  assign n25157 = ~n18074 ;
  assign n18080 = n25157 & n18079 ;
  assign n25158 = ~n18080 ;
  assign n18081 = n18073 & n25158 ;
  assign n18082 = x108 | n18081 ;
  assign n18083 = x108 & n18081 ;
  assign n25159 = ~n17521 ;
  assign n18084 = n25159 & n17522 ;
  assign n18085 = n130 & n18084 ;
  assign n18086 = n24938 & n18085 ;
  assign n25160 = ~n18085 ;
  assign n18087 = n17527 & n25160 ;
  assign n18088 = n18086 | n18087 ;
  assign n25161 = ~n18083 ;
  assign n18089 = n25161 & n18088 ;
  assign n25162 = ~n18089 ;
  assign n18090 = n18082 & n25162 ;
  assign n18091 = x109 | n18090 ;
  assign n18092 = x109 & n18090 ;
  assign n25163 = ~n17530 ;
  assign n18093 = n25163 & n17531 ;
  assign n18094 = n130 & n18093 ;
  assign n18095 = n24941 & n18094 ;
  assign n25164 = ~n18094 ;
  assign n18096 = n17536 & n25164 ;
  assign n18097 = n18095 | n18096 ;
  assign n25165 = ~n18092 ;
  assign n18098 = n25165 & n18097 ;
  assign n25166 = ~n18098 ;
  assign n18099 = n18091 & n25166 ;
  assign n18100 = x110 | n18099 ;
  assign n18101 = x110 & n18099 ;
  assign n25167 = ~n17539 ;
  assign n18102 = n25167 & n17540 ;
  assign n18103 = n130 & n18102 ;
  assign n18104 = n17545 & n18103 ;
  assign n18105 = n17545 | n18103 ;
  assign n25168 = ~n18104 ;
  assign n18106 = n25168 & n18105 ;
  assign n25169 = ~n18101 ;
  assign n18107 = n25169 & n18106 ;
  assign n25170 = ~n18107 ;
  assign n18108 = n18100 & n25170 ;
  assign n18109 = x111 | n18108 ;
  assign n18110 = x111 & n18108 ;
  assign n25171 = ~n17548 ;
  assign n18111 = n25171 & n17549 ;
  assign n18112 = n130 & n18111 ;
  assign n18113 = n17554 & n18112 ;
  assign n18114 = n17554 | n18112 ;
  assign n25172 = ~n18113 ;
  assign n18115 = n25172 & n18114 ;
  assign n25173 = ~n18110 ;
  assign n18116 = n25173 & n18115 ;
  assign n25174 = ~n18116 ;
  assign n18117 = n18109 & n25174 ;
  assign n18118 = x112 | n18117 ;
  assign n18119 = x112 & n18117 ;
  assign n25175 = ~n17557 ;
  assign n18120 = n25175 & n17558 ;
  assign n18121 = n130 & n18120 ;
  assign n18122 = n24949 & n18121 ;
  assign n25176 = ~n18121 ;
  assign n18123 = n17563 & n25176 ;
  assign n18124 = n18122 | n18123 ;
  assign n25177 = ~n18119 ;
  assign n18125 = n25177 & n18124 ;
  assign n25178 = ~n18125 ;
  assign n18126 = n18118 & n25178 ;
  assign n18127 = x113 | n18126 ;
  assign n18128 = x113 & n18126 ;
  assign n25179 = ~n17566 ;
  assign n18129 = n25179 & n17567 ;
  assign n18130 = n130 & n18129 ;
  assign n18131 = n24952 & n18130 ;
  assign n25180 = ~n18130 ;
  assign n18132 = n17572 & n25180 ;
  assign n18133 = n18131 | n18132 ;
  assign n25181 = ~n18128 ;
  assign n18134 = n25181 & n18133 ;
  assign n25182 = ~n18134 ;
  assign n18135 = n18127 & n25182 ;
  assign n18136 = x114 | n18135 ;
  assign n18137 = x114 & n18135 ;
  assign n25183 = ~n17575 ;
  assign n18138 = n25183 & n17576 ;
  assign n18139 = n130 & n18138 ;
  assign n18140 = n17581 & n18139 ;
  assign n18141 = n17581 | n18139 ;
  assign n25184 = ~n18140 ;
  assign n18142 = n25184 & n18141 ;
  assign n25185 = ~n18137 ;
  assign n18143 = n25185 & n18142 ;
  assign n25186 = ~n18143 ;
  assign n18144 = n18136 & n25186 ;
  assign n18145 = x115 | n18144 ;
  assign n18146 = x115 & n18144 ;
  assign n25187 = ~n17584 ;
  assign n18147 = n25187 & n17585 ;
  assign n18148 = n130 & n18147 ;
  assign n18149 = n17590 & n18148 ;
  assign n18150 = n17590 | n18148 ;
  assign n25188 = ~n18149 ;
  assign n18151 = n25188 & n18150 ;
  assign n25189 = ~n18146 ;
  assign n18152 = n25189 & n18151 ;
  assign n25190 = ~n18152 ;
  assign n18153 = n18145 & n25190 ;
  assign n18154 = x116 | n18153 ;
  assign n18155 = x116 & n18153 ;
  assign n25191 = ~n17593 ;
  assign n18156 = n25191 & n17594 ;
  assign n18157 = n130 & n18156 ;
  assign n18158 = n17599 & n18157 ;
  assign n18159 = n17599 | n18157 ;
  assign n25192 = ~n18158 ;
  assign n18160 = n25192 & n18159 ;
  assign n25193 = ~n18155 ;
  assign n18161 = n25193 & n18160 ;
  assign n25194 = ~n18161 ;
  assign n18162 = n18154 & n25194 ;
  assign n18163 = x117 | n18162 ;
  assign n18164 = x117 & n18162 ;
  assign n25195 = ~n17602 ;
  assign n18165 = n25195 & n17603 ;
  assign n18166 = n130 & n18165 ;
  assign n18167 = n17608 & n18166 ;
  assign n18168 = n17608 | n18166 ;
  assign n25196 = ~n18167 ;
  assign n18169 = n25196 & n18168 ;
  assign n25197 = ~n18164 ;
  assign n18170 = n25197 & n18169 ;
  assign n25198 = ~n18170 ;
  assign n18171 = n18163 & n25198 ;
  assign n18172 = x118 | n18171 ;
  assign n18173 = x118 & n18171 ;
  assign n25199 = ~n17611 ;
  assign n18174 = n25199 & n17612 ;
  assign n18175 = n130 & n18174 ;
  assign n18176 = n24965 & n18175 ;
  assign n25200 = ~n18175 ;
  assign n18177 = n17617 & n25200 ;
  assign n18178 = n18176 | n18177 ;
  assign n25201 = ~n18173 ;
  assign n18179 = n25201 & n18178 ;
  assign n25202 = ~n18179 ;
  assign n18180 = n18172 & n25202 ;
  assign n18181 = x119 | n18180 ;
  assign n18182 = x119 & n18180 ;
  assign n25203 = ~n17620 ;
  assign n18183 = n25203 & n17621 ;
  assign n18184 = n130 & n18183 ;
  assign n18185 = n17626 & n18184 ;
  assign n18186 = n17626 | n18184 ;
  assign n25204 = ~n18185 ;
  assign n18187 = n25204 & n18186 ;
  assign n25205 = ~n18182 ;
  assign n18188 = n25205 & n18187 ;
  assign n25206 = ~n18188 ;
  assign n18189 = n18181 & n25206 ;
  assign n18190 = x120 | n18189 ;
  assign n18191 = x120 & n18189 ;
  assign n25207 = ~n17629 ;
  assign n18192 = n25207 & n17630 ;
  assign n18193 = n130 & n18192 ;
  assign n18194 = n24970 & n18193 ;
  assign n25208 = ~n18193 ;
  assign n18195 = n17635 & n25208 ;
  assign n18196 = n18194 | n18195 ;
  assign n25209 = ~n18191 ;
  assign n18197 = n25209 & n18196 ;
  assign n25210 = ~n18197 ;
  assign n18198 = n18190 & n25210 ;
  assign n18199 = x121 | n18198 ;
  assign n18200 = x121 & n18198 ;
  assign n25211 = ~n17638 ;
  assign n18201 = n25211 & n17639 ;
  assign n18202 = n130 & n18201 ;
  assign n18203 = n17644 & n18202 ;
  assign n18204 = n17644 | n18202 ;
  assign n25212 = ~n18203 ;
  assign n18205 = n25212 & n18204 ;
  assign n25213 = ~n18200 ;
  assign n18206 = n25213 & n18205 ;
  assign n25214 = ~n18206 ;
  assign n18207 = n18199 & n25214 ;
  assign n18208 = x122 | n18207 ;
  assign n18209 = x122 & n18207 ;
  assign n25215 = ~n17647 ;
  assign n18210 = n25215 & n17648 ;
  assign n18211 = n130 & n18210 ;
  assign n18212 = n24975 & n18211 ;
  assign n25216 = ~n18211 ;
  assign n18213 = n17653 & n25216 ;
  assign n18214 = n18212 | n18213 ;
  assign n25217 = ~n18209 ;
  assign n18215 = n25217 & n18214 ;
  assign n25218 = ~n18215 ;
  assign n18216 = n18208 & n25218 ;
  assign n18217 = x123 | n18216 ;
  assign n18218 = x123 & n18216 ;
  assign n25219 = ~n17656 ;
  assign n18219 = n25219 & n17657 ;
  assign n18220 = n130 & n18219 ;
  assign n18221 = n24978 & n18220 ;
  assign n25220 = ~n18220 ;
  assign n18222 = n17662 & n25220 ;
  assign n18223 = n18221 | n18222 ;
  assign n25221 = ~n18218 ;
  assign n18224 = n25221 & n18223 ;
  assign n25222 = ~n18224 ;
  assign n18225 = n18217 & n25222 ;
  assign n18226 = x124 | n18225 ;
  assign n18227 = x124 & n18225 ;
  assign n25223 = ~n17665 ;
  assign n18228 = n25223 & n17666 ;
  assign n18229 = n130 & n18228 ;
  assign n18230 = n24981 & n18229 ;
  assign n25224 = ~n18229 ;
  assign n18231 = n17671 & n25224 ;
  assign n18232 = n18230 | n18231 ;
  assign n25225 = ~n18227 ;
  assign n18233 = n25225 & n18232 ;
  assign n25226 = ~n18233 ;
  assign n18234 = n18226 & n25226 ;
  assign n18235 = x125 | n18234 ;
  assign n18236 = x125 & n18234 ;
  assign n25227 = ~n17674 ;
  assign n18237 = n25227 & n17675 ;
  assign n18238 = n130 & n18237 ;
  assign n18239 = n24984 & n18238 ;
  assign n25228 = ~n18238 ;
  assign n18240 = n17680 & n25228 ;
  assign n18241 = n18239 | n18240 ;
  assign n25229 = ~n18236 ;
  assign n18242 = n25229 & n18241 ;
  assign n25230 = ~n18242 ;
  assign n18243 = n18235 & n25230 ;
  assign n18244 = x126 | n18243 ;
  assign n25231 = ~n17683 ;
  assign n18245 = n25231 & n17684 ;
  assign n18246 = n130 & n18245 ;
  assign n18247 = n17690 & n18246 ;
  assign n18248 = n17690 | n18246 ;
  assign n25232 = ~n18247 ;
  assign n18249 = n25232 & n18248 ;
  assign n18250 = x126 & n18243 ;
  assign n25233 = ~n18250 ;
  assign n18251 = n18249 & n25233 ;
  assign n25234 = ~n18251 ;
  assign n18252 = n18244 & n25234 ;
  assign n25235 = ~n18252 ;
  assign n18253 = n17140 & n25235 ;
  assign n25236 = ~n18253 ;
  assign n18256 = x127 & n25236 ;
  assign n25237 = ~n17696 ;
  assign n18254 = n17693 & n25237 ;
  assign n25238 = ~n18254 ;
  assign n18255 = n17140 & n25238 ;
  assign n25239 = ~n18255 ;
  assign n18257 = n18252 & n25239 ;
  assign n18258 = n18256 | n18257 ;
  assign n18358 = x65 | x66 ;
  assign n18359 = n18585 & x64 ;
  assign n18360 = n18358 | n18359 ;
  assign n18361 = n18563 | n18360 ;
  assign n129 = ~n18258 ;
  assign n18354 = x64 & n129 ;
  assign n18355 = x0 & n18354 ;
  assign n18356 = x0 | n18354 ;
  assign n25241 = ~n18355 ;
  assign n193 = n25241 & n18356 ;
  assign n18349 = n5490 & n24991 ;
  assign n18350 = n129 & n18349 ;
  assign n18351 = n17701 | n18350 ;
  assign n18352 = n17701 & n18350 ;
  assign n25242 = ~n18352 ;
  assign n194 = n18351 & n25242 ;
  assign n18344 = n17704 & n129 ;
  assign n18345 = n17711 & n18344 ;
  assign n18346 = n24994 & n18344 ;
  assign n18347 = n17709 | n18346 ;
  assign n25243 = ~n18345 ;
  assign n195 = n25243 & n18347 ;
  assign n18339 = n17713 & n129 ;
  assign n18340 = n17720 & n18339 ;
  assign n18341 = n24997 & n18339 ;
  assign n18342 = n17718 | n18341 ;
  assign n25244 = ~n18340 ;
  assign n196 = n25244 & n18342 ;
  assign n18334 = n17722 & n25001 ;
  assign n18335 = n129 & n18334 ;
  assign n18336 = n17728 | n18335 ;
  assign n18337 = n17728 & n18335 ;
  assign n25245 = ~n18337 ;
  assign n197 = n18336 & n25245 ;
  assign n18574 = n17731 & n25005 ;
  assign n18575 = n129 & n18574 ;
  assign n18576 = n17737 | n18575 ;
  assign n18577 = n17737 & n18575 ;
  assign n25246 = ~n18577 ;
  assign n198 = n18576 & n25246 ;
  assign n18329 = n17740 & n25009 ;
  assign n18330 = n129 & n18329 ;
  assign n18331 = n17746 & n18330 ;
  assign n18332 = n17746 | n18330 ;
  assign n25247 = ~n18331 ;
  assign n199 = n25247 & n18332 ;
  assign n18569 = n17749 & n25013 ;
  assign n18570 = n129 & n18569 ;
  assign n18571 = n17755 | n18570 ;
  assign n18572 = n17755 & n18570 ;
  assign n25248 = ~n18572 ;
  assign n200 = n18571 & n25248 ;
  assign n18564 = n17758 & n25017 ;
  assign n18565 = n129 & n18564 ;
  assign n18566 = n17764 & n18565 ;
  assign n18567 = n17764 | n18565 ;
  assign n25249 = ~n18566 ;
  assign n201 = n25249 & n18567 ;
  assign n18559 = n17767 & n25021 ;
  assign n18560 = n129 & n18559 ;
  assign n18561 = n17773 | n18560 ;
  assign n18562 = n17773 & n18560 ;
  assign n25250 = ~n18562 ;
  assign n202 = n18561 & n25250 ;
  assign n18554 = n17776 & n25025 ;
  assign n18555 = n129 & n18554 ;
  assign n18556 = n17782 | n18555 ;
  assign n18557 = n17782 & n18555 ;
  assign n25251 = ~n18557 ;
  assign n203 = n18556 & n25251 ;
  assign n18549 = n17785 & n25029 ;
  assign n18550 = n129 & n18549 ;
  assign n18551 = n17791 | n18550 ;
  assign n18552 = n17791 & n18550 ;
  assign n25252 = ~n18552 ;
  assign n204 = n18551 & n25252 ;
  assign n18324 = n17794 & n25033 ;
  assign n18325 = n129 & n18324 ;
  assign n18326 = n17800 & n18325 ;
  assign n18327 = n17800 | n18325 ;
  assign n25253 = ~n18326 ;
  assign n205 = n25253 & n18327 ;
  assign n18544 = n17803 & n25037 ;
  assign n18545 = n129 & n18544 ;
  assign n18546 = n17809 & n18545 ;
  assign n18547 = n17809 | n18545 ;
  assign n25254 = ~n18546 ;
  assign n206 = n25254 & n18547 ;
  assign n18319 = n17812 & n25041 ;
  assign n18320 = n129 & n18319 ;
  assign n18321 = n17818 & n18320 ;
  assign n18322 = n17818 | n18320 ;
  assign n25255 = ~n18321 ;
  assign n207 = n25255 & n18322 ;
  assign n18539 = n17821 & n25045 ;
  assign n18540 = n129 & n18539 ;
  assign n18541 = n17827 | n18540 ;
  assign n18542 = n17827 & n18540 ;
  assign n25256 = ~n18542 ;
  assign n208 = n18541 & n25256 ;
  assign n18534 = n17830 & n25049 ;
  assign n18535 = n129 & n18534 ;
  assign n18536 = n17836 | n18535 ;
  assign n18537 = n17836 & n18535 ;
  assign n25257 = ~n18537 ;
  assign n209 = n18536 & n25257 ;
  assign n18529 = n17839 & n25053 ;
  assign n18530 = n129 & n18529 ;
  assign n18531 = n17845 | n18530 ;
  assign n18532 = n17845 & n18530 ;
  assign n25258 = ~n18532 ;
  assign n210 = n18531 & n25258 ;
  assign n18524 = n17848 & n25057 ;
  assign n18525 = n129 & n18524 ;
  assign n18526 = n17854 | n18525 ;
  assign n18527 = n17854 & n18525 ;
  assign n25259 = ~n18527 ;
  assign n211 = n18526 & n25259 ;
  assign n18314 = n17857 & n25061 ;
  assign n18315 = n129 & n18314 ;
  assign n18316 = n17863 & n18315 ;
  assign n18317 = n17863 | n18315 ;
  assign n25260 = ~n18316 ;
  assign n212 = n25260 & n18317 ;
  assign n18519 = n17866 & n25065 ;
  assign n18520 = n129 & n18519 ;
  assign n18521 = n17872 & n18520 ;
  assign n18522 = n17872 | n18520 ;
  assign n25261 = ~n18521 ;
  assign n213 = n25261 & n18522 ;
  assign n18514 = n17875 & n25069 ;
  assign n18515 = n129 & n18514 ;
  assign n18516 = n17881 | n18515 ;
  assign n18517 = n17881 & n18515 ;
  assign n25262 = ~n18517 ;
  assign n214 = n18516 & n25262 ;
  assign n18509 = n17884 & n25073 ;
  assign n18510 = n129 & n18509 ;
  assign n18511 = n17890 & n18510 ;
  assign n18512 = n17890 | n18510 ;
  assign n25263 = ~n18511 ;
  assign n215 = n25263 & n18512 ;
  assign n18309 = n17893 & n25077 ;
  assign n18310 = n129 & n18309 ;
  assign n18311 = n17899 | n18310 ;
  assign n18312 = n17899 & n18310 ;
  assign n25264 = ~n18312 ;
  assign n216 = n18311 & n25264 ;
  assign n18504 = n17902 & n25081 ;
  assign n18505 = n129 & n18504 ;
  assign n18506 = n17908 | n18505 ;
  assign n18507 = n17908 & n18505 ;
  assign n25265 = ~n18507 ;
  assign n217 = n18506 & n25265 ;
  assign n18499 = n17911 & n25085 ;
  assign n18500 = n129 & n18499 ;
  assign n18501 = n17917 | n18500 ;
  assign n18502 = n17917 & n18500 ;
  assign n25266 = ~n18502 ;
  assign n218 = n18501 & n25266 ;
  assign n18304 = n17920 & n25089 ;
  assign n18305 = n129 & n18304 ;
  assign n18306 = n17926 & n18305 ;
  assign n18307 = n17926 | n18305 ;
  assign n25267 = ~n18306 ;
  assign n219 = n25267 & n18307 ;
  assign n18494 = n17929 & n25093 ;
  assign n18495 = n129 & n18494 ;
  assign n18496 = n17935 | n18495 ;
  assign n18497 = n17935 & n18495 ;
  assign n25268 = ~n18497 ;
  assign n220 = n18496 & n25268 ;
  assign n18489 = n17938 & n25097 ;
  assign n18490 = n129 & n18489 ;
  assign n18491 = n17944 | n18490 ;
  assign n18492 = n17944 & n18490 ;
  assign n25269 = ~n18492 ;
  assign n221 = n18491 & n25269 ;
  assign n18299 = n17947 & n25101 ;
  assign n18300 = n129 & n18299 ;
  assign n18301 = n17953 & n18300 ;
  assign n18302 = n17953 | n18300 ;
  assign n25270 = ~n18301 ;
  assign n222 = n25270 & n18302 ;
  assign n18484 = n17956 & n25105 ;
  assign n18485 = n129 & n18484 ;
  assign n18486 = n17962 | n18485 ;
  assign n18487 = n17962 & n18485 ;
  assign n25271 = ~n18487 ;
  assign n223 = n18486 & n25271 ;
  assign n18479 = n17965 & n25109 ;
  assign n18480 = n129 & n18479 ;
  assign n18481 = n17971 | n18480 ;
  assign n18482 = n17971 & n18480 ;
  assign n25272 = ~n18482 ;
  assign n224 = n18481 & n25272 ;
  assign n18474 = n17974 & n25113 ;
  assign n18475 = n129 & n18474 ;
  assign n18476 = n17980 | n18475 ;
  assign n18477 = n17980 & n18475 ;
  assign n25273 = ~n18477 ;
  assign n225 = n18476 & n25273 ;
  assign n18294 = n17983 & n25117 ;
  assign n18295 = n129 & n18294 ;
  assign n18296 = n17989 | n18295 ;
  assign n18297 = n17989 & n18295 ;
  assign n25274 = ~n18297 ;
  assign n226 = n18296 & n25274 ;
  assign n18289 = n17992 & n25121 ;
  assign n18290 = n129 & n18289 ;
  assign n18291 = n17998 & n18290 ;
  assign n18292 = n17998 | n18290 ;
  assign n25275 = ~n18291 ;
  assign n227 = n25275 & n18292 ;
  assign n18469 = n18001 & n25125 ;
  assign n18470 = n129 & n18469 ;
  assign n18471 = n18007 | n18470 ;
  assign n18472 = n18007 & n18470 ;
  assign n25276 = ~n18472 ;
  assign n228 = n18471 & n25276 ;
  assign n18464 = n18010 & n25129 ;
  assign n18465 = n129 & n18464 ;
  assign n18466 = n18016 | n18465 ;
  assign n18467 = n18016 & n18465 ;
  assign n25277 = ~n18467 ;
  assign n229 = n18466 & n25277 ;
  assign n18284 = n18019 & n25133 ;
  assign n18285 = n129 & n18284 ;
  assign n18286 = n18025 & n18285 ;
  assign n18287 = n18025 | n18285 ;
  assign n25278 = ~n18286 ;
  assign n230 = n25278 & n18287 ;
  assign n18459 = n18028 & n25137 ;
  assign n18460 = n129 & n18459 ;
  assign n18461 = n18034 | n18460 ;
  assign n18462 = n18034 & n18460 ;
  assign n25279 = ~n18462 ;
  assign n231 = n18461 & n25279 ;
  assign n18454 = n18037 & n25141 ;
  assign n18455 = n129 & n18454 ;
  assign n18456 = n18043 | n18455 ;
  assign n18457 = n18043 & n18455 ;
  assign n25280 = ~n18457 ;
  assign n232 = n18456 & n25280 ;
  assign n18449 = n18046 & n25145 ;
  assign n18450 = n129 & n18449 ;
  assign n18451 = n18052 | n18450 ;
  assign n18452 = n18052 & n18450 ;
  assign n25281 = ~n18452 ;
  assign n233 = n18451 & n25281 ;
  assign n18444 = n18055 & n25149 ;
  assign n18445 = n129 & n18444 ;
  assign n18446 = n18061 | n18445 ;
  assign n18447 = n18061 & n18445 ;
  assign n25282 = ~n18447 ;
  assign n234 = n18446 & n25282 ;
  assign n18439 = n18064 & n25153 ;
  assign n18440 = n129 & n18439 ;
  assign n18441 = n18070 | n18440 ;
  assign n18442 = n18070 & n18440 ;
  assign n25283 = ~n18442 ;
  assign n235 = n18441 & n25283 ;
  assign n18279 = n18073 & n25157 ;
  assign n18280 = n129 & n18279 ;
  assign n18281 = n18079 & n18280 ;
  assign n18282 = n18079 | n18280 ;
  assign n25284 = ~n18281 ;
  assign n236 = n25284 & n18282 ;
  assign n18434 = n18082 & n25161 ;
  assign n18435 = n129 & n18434 ;
  assign n18436 = n18088 | n18435 ;
  assign n18437 = n18088 & n18435 ;
  assign n25285 = ~n18437 ;
  assign n237 = n18436 & n25285 ;
  assign n18429 = n18091 & n25165 ;
  assign n18430 = n129 & n18429 ;
  assign n18431 = n18097 | n18430 ;
  assign n18432 = n18097 & n18430 ;
  assign n25286 = ~n18432 ;
  assign n238 = n18431 & n25286 ;
  assign n18274 = n18100 & n25169 ;
  assign n18275 = n129 & n18274 ;
  assign n18276 = n18106 & n18275 ;
  assign n18277 = n18106 | n18275 ;
  assign n25287 = ~n18276 ;
  assign n239 = n25287 & n18277 ;
  assign n18424 = n18109 & n25173 ;
  assign n18425 = n129 & n18424 ;
  assign n18426 = n18115 & n18425 ;
  assign n18427 = n18115 | n18425 ;
  assign n25288 = ~n18426 ;
  assign n240 = n25288 & n18427 ;
  assign n18419 = n18118 & n25177 ;
  assign n18420 = n129 & n18419 ;
  assign n18421 = n18124 | n18420 ;
  assign n18422 = n18124 & n18420 ;
  assign n25289 = ~n18422 ;
  assign n241 = n18421 & n25289 ;
  assign n18414 = n18127 & n25181 ;
  assign n18415 = n129 & n18414 ;
  assign n18416 = n18133 | n18415 ;
  assign n18417 = n18133 & n18415 ;
  assign n25290 = ~n18417 ;
  assign n242 = n18416 & n25290 ;
  assign n18269 = n18136 & n25185 ;
  assign n18270 = n129 & n18269 ;
  assign n18271 = n18142 & n18270 ;
  assign n18272 = n18142 | n18270 ;
  assign n25291 = ~n18271 ;
  assign n243 = n25291 & n18272 ;
  assign n18264 = n18145 & n25189 ;
  assign n18265 = n129 & n18264 ;
  assign n18266 = n18151 & n18265 ;
  assign n18267 = n18151 | n18265 ;
  assign n25292 = ~n18266 ;
  assign n244 = n25292 & n18267 ;
  assign n18409 = n18154 & n25193 ;
  assign n18410 = n129 & n18409 ;
  assign n18411 = n18160 | n18410 ;
  assign n18412 = n18160 & n18410 ;
  assign n25293 = ~n18412 ;
  assign n245 = n18411 & n25293 ;
  assign n18404 = n18163 & n25197 ;
  assign n18405 = n129 & n18404 ;
  assign n18406 = n18169 | n18405 ;
  assign n18407 = n18169 & n18405 ;
  assign n25294 = ~n18407 ;
  assign n246 = n18406 & n25294 ;
  assign n18399 = n18172 & n25201 ;
  assign n18400 = n129 & n18399 ;
  assign n18401 = n18178 | n18400 ;
  assign n18402 = n18178 & n18400 ;
  assign n25295 = ~n18402 ;
  assign n247 = n18401 & n25295 ;
  assign n18394 = n18181 & n25205 ;
  assign n18395 = n129 & n18394 ;
  assign n18396 = n18187 | n18395 ;
  assign n18397 = n18187 & n18395 ;
  assign n25296 = ~n18397 ;
  assign n248 = n18396 & n25296 ;
  assign n18389 = n18190 & n25209 ;
  assign n18390 = n129 & n18389 ;
  assign n18391 = n18196 | n18390 ;
  assign n18392 = n18196 & n18390 ;
  assign n25297 = ~n18392 ;
  assign n249 = n18391 & n25297 ;
  assign n18384 = n18199 & n25213 ;
  assign n18385 = n129 & n18384 ;
  assign n18386 = n18205 | n18385 ;
  assign n18387 = n18205 & n18385 ;
  assign n25298 = ~n18387 ;
  assign n250 = n18386 & n25298 ;
  assign n18379 = n18208 & n25217 ;
  assign n18380 = n129 & n18379 ;
  assign n18381 = n18214 | n18380 ;
  assign n18382 = n18214 & n18380 ;
  assign n25299 = ~n18382 ;
  assign n251 = n18381 & n25299 ;
  assign n18374 = n18217 & n25221 ;
  assign n18375 = n129 & n18374 ;
  assign n18376 = n18223 | n18375 ;
  assign n18377 = n18223 & n18375 ;
  assign n25300 = ~n18377 ;
  assign n252 = n18376 & n25300 ;
  assign n18259 = n18226 & n25225 ;
  assign n18260 = n129 & n18259 ;
  assign n18261 = n18232 | n18260 ;
  assign n18262 = n18232 & n18260 ;
  assign n25301 = ~n18262 ;
  assign n253 = n18261 & n25301 ;
  assign n18369 = n18235 & n25229 ;
  assign n18370 = n129 & n18369 ;
  assign n18371 = n18241 | n18370 ;
  assign n18372 = n18241 & n18370 ;
  assign n25302 = ~n18372 ;
  assign n254 = n18371 & n25302 ;
  assign n18364 = n18244 & n25233 ;
  assign n18365 = n129 & n18364 ;
  assign n18366 = n18249 & n18365 ;
  assign n18367 = n18249 | n18365 ;
  assign n25303 = ~n18366 ;
  assign n255 = n25303 & n18367 ;
  assign n18362 = n18255 & n18256 ;
  assign n256 = n21884 | n18362 ;
  assign n192 = ~n18361 ;
  assign y0 = n129 ;
  assign y1 = n130 ;
  assign y2 = n131 ;
  assign y3 = n132 ;
  assign y4 = n133 ;
  assign y5 = n134 ;
  assign y6 = n135 ;
  assign y7 = n136 ;
  assign y8 = n137 ;
  assign y9 = n138 ;
  assign y10 = n139 ;
  assign y11 = n140 ;
  assign y12 = n141 ;
  assign y13 = n142 ;
  assign y14 = n143 ;
  assign y15 = n144 ;
  assign y16 = n145 ;
  assign y17 = n146 ;
  assign y18 = n147 ;
  assign y19 = n148 ;
  assign y20 = n149 ;
  assign y21 = n150 ;
  assign y22 = n151 ;
  assign y23 = n152 ;
  assign y24 = n153 ;
  assign y25 = n154 ;
  assign y26 = n155 ;
  assign y27 = n156 ;
  assign y28 = n157 ;
  assign y29 = n158 ;
  assign y30 = n159 ;
  assign y31 = n160 ;
  assign y32 = n161 ;
  assign y33 = n162 ;
  assign y34 = n163 ;
  assign y35 = n164 ;
  assign y36 = n165 ;
  assign y37 = n166 ;
  assign y38 = n167 ;
  assign y39 = n168 ;
  assign y40 = n169 ;
  assign y41 = n170 ;
  assign y42 = n171 ;
  assign y43 = n172 ;
  assign y44 = n173 ;
  assign y45 = n174 ;
  assign y46 = n175 ;
  assign y47 = n176 ;
  assign y48 = n177 ;
  assign y49 = n178 ;
  assign y50 = n179 ;
  assign y51 = n180 ;
  assign y52 = n181 ;
  assign y53 = n182 ;
  assign y54 = n183 ;
  assign y55 = n184 ;
  assign y56 = n185 ;
  assign y57 = n186 ;
  assign y58 = n187 ;
  assign y59 = n188 ;
  assign y60 = n189 ;
  assign y61 = n190 ;
  assign y62 = n191 ;
  assign y63 = n192 ;
  assign y64 = n193 ;
  assign y65 = n194 ;
  assign y66 = n195 ;
  assign y67 = n196 ;
  assign y68 = n197 ;
  assign y69 = n198 ;
  assign y70 = n199 ;
  assign y71 = n200 ;
  assign y72 = n201 ;
  assign y73 = n202 ;
  assign y74 = n203 ;
  assign y75 = n204 ;
  assign y76 = n205 ;
  assign y77 = n206 ;
  assign y78 = n207 ;
  assign y79 = n208 ;
  assign y80 = n209 ;
  assign y81 = n210 ;
  assign y82 = n211 ;
  assign y83 = n212 ;
  assign y84 = n213 ;
  assign y85 = n214 ;
  assign y86 = n215 ;
  assign y87 = n216 ;
  assign y88 = n217 ;
  assign y89 = n218 ;
  assign y90 = n219 ;
  assign y91 = n220 ;
  assign y92 = n221 ;
  assign y93 = n222 ;
  assign y94 = n223 ;
  assign y95 = n224 ;
  assign y96 = n225 ;
  assign y97 = n226 ;
  assign y98 = n227 ;
  assign y99 = n228 ;
  assign y100 = n229 ;
  assign y101 = n230 ;
  assign y102 = n231 ;
  assign y103 = n232 ;
  assign y104 = n233 ;
  assign y105 = n234 ;
  assign y106 = n235 ;
  assign y107 = n236 ;
  assign y108 = n237 ;
  assign y109 = n238 ;
  assign y110 = n239 ;
  assign y111 = n240 ;
  assign y112 = n241 ;
  assign y113 = n242 ;
  assign y114 = n243 ;
  assign y115 = n244 ;
  assign y116 = n245 ;
  assign y117 = n246 ;
  assign y118 = n247 ;
  assign y119 = n248 ;
  assign y120 = n249 ;
  assign y121 = n250 ;
  assign y122 = n251 ;
  assign y123 = n252 ;
  assign y124 = n253 ;
  assign y125 = n254 ;
  assign y126 = n255 ;
  assign y127 = n256 ;
endmodule
