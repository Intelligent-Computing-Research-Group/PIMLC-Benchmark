module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 ;
  assign n3384 = ~x255 ;
  assign n1134 = x127 & n3384 ;
  assign n3385 = ~x126 ;
  assign n3295 = n3385 & x254 ;
  assign n3386 = ~x125 ;
  assign n3297 = n3386 & x253 ;
  assign n1601 = n3295 | n3297 ;
  assign n3387 = ~x251 ;
  assign n1135 = x123 & n3387 ;
  assign n3388 = ~x122 ;
  assign n1594 = n3388 & x250 ;
  assign n3389 = ~x119 ;
  assign n1136 = n3389 & x247 ;
  assign n3390 = ~x246 ;
  assign n1137 = x118 & n3390 ;
  assign n3391 = ~x244 ;
  assign n1578 = x116 & n3391 ;
  assign n3392 = ~x245 ;
  assign n1579 = x117 & n3392 ;
  assign n1580 = n1578 | n1579 ;
  assign n3393 = ~x243 ;
  assign n1138 = x115 & n3393 ;
  assign n3394 = ~x114 ;
  assign n1139 = n3394 & x242 ;
  assign n3395 = ~x241 ;
  assign n1568 = x113 & n3395 ;
  assign n3396 = ~x242 ;
  assign n1569 = x114 & n3396 ;
  assign n1570 = n1568 | n1569 ;
  assign n3397 = ~x240 ;
  assign n1140 = x112 & n3397 ;
  assign n3398 = ~x111 ;
  assign n1141 = n3398 & x239 ;
  assign n3399 = ~x238 ;
  assign n1558 = x110 & n3399 ;
  assign n3400 = ~x239 ;
  assign n1559 = x111 & n3400 ;
  assign n1560 = n1558 | n1559 ;
  assign n3401 = ~x110 ;
  assign n1142 = n3401 & x238 ;
  assign n3402 = ~x237 ;
  assign n1143 = x109 & n3402 ;
  assign n3403 = ~x236 ;
  assign n1548 = x108 & n3403 ;
  assign n3404 = ~x235 ;
  assign n1549 = x107 & n3404 ;
  assign n1550 = n1548 | n1549 ;
  assign n3405 = ~x107 ;
  assign n1144 = n3405 & x235 ;
  assign n3406 = ~x234 ;
  assign n1145 = x106 & n3406 ;
  assign n3407 = ~x233 ;
  assign n1538 = x105 & n3407 ;
  assign n3408 = ~x232 ;
  assign n1539 = x104 & n3408 ;
  assign n1540 = n1538 | n1539 ;
  assign n3409 = ~x102 ;
  assign n1146 = n3409 & x230 ;
  assign n3410 = ~x229 ;
  assign n1527 = x101 & n3410 ;
  assign n3411 = ~x99 ;
  assign n1147 = n3411 & x227 ;
  assign n3412 = ~x226 ;
  assign n1517 = x98 & n3412 ;
  assign n3413 = ~x225 ;
  assign n1148 = x97 & n3413 ;
  assign n3414 = ~x96 ;
  assign n1149 = n3414 & x224 ;
  assign n3415 = ~x223 ;
  assign n1508 = x95 & n3415 ;
  assign n3416 = ~x224 ;
  assign n1509 = x96 & n3416 ;
  assign n1510 = n1508 | n1509 ;
  assign n3417 = ~x220 ;
  assign n1492 = x92 & n3417 ;
  assign n3418 = ~x219 ;
  assign n1493 = x91 & n3418 ;
  assign n1494 = n1492 | n1493 ;
  assign n3419 = ~x91 ;
  assign n1150 = n3419 & x219 ;
  assign n3420 = ~x218 ;
  assign n1151 = x90 & n3420 ;
  assign n3421 = ~x216 ;
  assign n1482 = x88 & n3421 ;
  assign n3422 = ~x217 ;
  assign n1483 = x89 & n3422 ;
  assign n1484 = n1482 | n1483 ;
  assign n3423 = ~x215 ;
  assign n1152 = x87 & n3423 ;
  assign n3424 = ~x86 ;
  assign n1153 = n3424 & x214 ;
  assign n3425 = ~x213 ;
  assign n1472 = x85 & n3425 ;
  assign n3426 = ~x214 ;
  assign n1473 = x86 & n3426 ;
  assign n1474 = n1472 | n1473 ;
  assign n3427 = ~x212 ;
  assign n1154 = x84 & n3427 ;
  assign n3428 = ~x83 ;
  assign n1155 = n3428 & x211 ;
  assign n3429 = ~x211 ;
  assign n1462 = x83 & n3429 ;
  assign n3430 = ~x210 ;
  assign n1463 = x82 & n3430 ;
  assign n1464 = n1462 | n1463 ;
  assign n3431 = ~x209 ;
  assign n1156 = x81 & n3431 ;
  assign n3432 = ~x80 ;
  assign n1157 = n3432 & x208 ;
  assign n3433 = ~x208 ;
  assign n1452 = x80 & n3433 ;
  assign n3434 = ~x207 ;
  assign n1453 = x79 & n3434 ;
  assign n1454 = n1452 | n1453 ;
  assign n3435 = ~x206 ;
  assign n1158 = x78 & n3435 ;
  assign n3436 = ~x77 ;
  assign n1159 = n3436 & x205 ;
  assign n3437 = ~x205 ;
  assign n1442 = x77 & n3437 ;
  assign n3438 = ~x204 ;
  assign n1443 = x76 & n3438 ;
  assign n1444 = n1442 | n1443 ;
  assign n3439 = ~x203 ;
  assign n1160 = x75 & n3439 ;
  assign n3440 = ~x74 ;
  assign n1161 = n3440 & x202 ;
  assign n3441 = ~x202 ;
  assign n1432 = x74 & n3441 ;
  assign n3442 = ~x201 ;
  assign n1433 = x73 & n3442 ;
  assign n1434 = n1432 | n1433 ;
  assign n3443 = ~x69 ;
  assign n1409 = n3443 & x197 ;
  assign n3444 = ~x196 ;
  assign n1413 = x68 & n3444 ;
  assign n3445 = ~n1409 ;
  assign n1414 = n3445 & n1413 ;
  assign n3446 = ~x197 ;
  assign n1415 = x69 & n3446 ;
  assign n3447 = ~x198 ;
  assign n1416 = x70 & n3447 ;
  assign n1417 = n1415 | n1416 ;
  assign n1418 = n1414 | n1417 ;
  assign n3448 = ~x193 ;
  assign n1396 = x65 & n3448 ;
  assign n3449 = ~x192 ;
  assign n1397 = x64 & n3449 ;
  assign n1398 = n1396 | n1397 ;
  assign n3450 = ~x191 ;
  assign n1162 = x63 & n3450 ;
  assign n3451 = ~x62 ;
  assign n1163 = n3451 & x190 ;
  assign n3452 = ~x190 ;
  assign n1164 = x62 & n3452 ;
  assign n3453 = ~x61 ;
  assign n1165 = n3453 & x189 ;
  assign n3454 = ~x186 ;
  assign n1376 = x58 & n3454 ;
  assign n3455 = ~x187 ;
  assign n1377 = x59 & n3455 ;
  assign n1378 = n1376 | n1377 ;
  assign n3456 = ~x58 ;
  assign n1166 = n3456 & x186 ;
  assign n3457 = ~x185 ;
  assign n1167 = x57 & n3457 ;
  assign n3458 = ~x184 ;
  assign n1369 = x56 & n3458 ;
  assign n3459 = ~x55 ;
  assign n1168 = n3459 & x183 ;
  assign n3460 = ~x181 ;
  assign n1359 = x53 & n3460 ;
  assign n3461 = ~x52 ;
  assign n1169 = n3461 & x180 ;
  assign n3462 = ~x51 ;
  assign n1170 = n3462 & x179 ;
  assign n3463 = ~x178 ;
  assign n1351 = x50 & n3463 ;
  assign n3464 = ~x177 ;
  assign n1171 = x49 & n3464 ;
  assign n3465 = ~x48 ;
  assign n1172 = n3465 & x176 ;
  assign n3466 = ~x175 ;
  assign n1342 = x47 & n3466 ;
  assign n3467 = ~x176 ;
  assign n1343 = x48 & n3467 ;
  assign n1344 = n1342 | n1343 ;
  assign n3468 = ~x47 ;
  assign n1173 = n3468 & x175 ;
  assign n3469 = ~x174 ;
  assign n1174 = x46 & n3469 ;
  assign n3470 = ~x173 ;
  assign n1332 = x45 & n3470 ;
  assign n3471 = ~x172 ;
  assign n1333 = x44 & n3471 ;
  assign n1334 = n1332 | n1333 ;
  assign n3472 = ~x44 ;
  assign n1175 = n3472 & x172 ;
  assign n3473 = ~x171 ;
  assign n1176 = x43 & n3473 ;
  assign n3474 = ~x41 ;
  assign n1315 = n3474 & x169 ;
  assign n3475 = ~x168 ;
  assign n1319 = x40 & n3475 ;
  assign n3476 = ~n1315 ;
  assign n1320 = n3476 & n1319 ;
  assign n3477 = ~x169 ;
  assign n1321 = x41 & n3477 ;
  assign n3478 = ~x170 ;
  assign n1322 = x42 & n3478 ;
  assign n1323 = n1321 | n1322 ;
  assign n1324 = n1320 | n1323 ;
  assign n3479 = ~x165 ;
  assign n1302 = x37 & n3479 ;
  assign n3480 = ~x164 ;
  assign n1303 = x36 & n3480 ;
  assign n1304 = n1302 | n1303 ;
  assign n3481 = ~x163 ;
  assign n1177 = x35 & n3481 ;
  assign n3482 = ~x34 ;
  assign n1178 = n3482 & x162 ;
  assign n3483 = ~x162 ;
  assign n1179 = x34 & n3483 ;
  assign n3484 = ~x33 ;
  assign n1180 = n3484 & x161 ;
  assign n3485 = ~x159 ;
  assign n1282 = x31 & n3485 ;
  assign n3486 = ~x158 ;
  assign n1283 = x30 & n3486 ;
  assign n1284 = n1282 | n1283 ;
  assign n3487 = ~x30 ;
  assign n1181 = n3487 & x158 ;
  assign n3488 = ~x157 ;
  assign n1182 = x29 & n3488 ;
  assign n3489 = ~x156 ;
  assign n1272 = x28 & n3489 ;
  assign n3490 = ~x155 ;
  assign n1273 = x27 & n3490 ;
  assign n1274 = n1272 | n1273 ;
  assign n3491 = ~x154 ;
  assign n1183 = x26 & n3491 ;
  assign n3492 = ~x25 ;
  assign n1184 = n3492 & x153 ;
  assign n3493 = ~x153 ;
  assign n1262 = x25 & n3493 ;
  assign n3494 = ~x152 ;
  assign n1263 = x24 & n3494 ;
  assign n1264 = n1262 | n1263 ;
  assign n3495 = ~x22 ;
  assign n1185 = n3495 & x150 ;
  assign n3496 = ~x149 ;
  assign n1251 = x21 & n3496 ;
  assign n3497 = ~x145 ;
  assign n1236 = x17 & n3497 ;
  assign n3498 = ~x146 ;
  assign n1237 = x18 & n3498 ;
  assign n1238 = n1236 | n1237 ;
  assign n3499 = ~x17 ;
  assign n1186 = n3499 & x145 ;
  assign n3500 = ~x144 ;
  assign n1187 = x16 & n3500 ;
  assign n3501 = ~x143 ;
  assign n1229 = x15 & n3501 ;
  assign n3502 = ~x14 ;
  assign n1188 = n3502 & x142 ;
  assign n3503 = ~x13 ;
  assign n1189 = n3503 & x141 ;
  assign n3504 = ~x140 ;
  assign n1221 = x12 & n3504 ;
  assign n3505 = ~x10 ;
  assign n1190 = n3505 & x138 ;
  assign n3506 = ~x137 ;
  assign n1214 = x9 & n3506 ;
  assign n3507 = ~x136 ;
  assign n3243 = x8 & n3507 ;
  assign n3508 = ~x7 ;
  assign n1191 = n3508 & x135 ;
  assign n3509 = ~x134 ;
  assign n3239 = x6 & n3509 ;
  assign n3510 = ~x135 ;
  assign n3241 = x7 & n3510 ;
  assign n1208 = n3239 | n3241 ;
  assign n3511 = ~x131 ;
  assign n3229 = x3 & n3511 ;
  assign n3512 = ~x130 ;
  assign n3233 = x2 & n3512 ;
  assign n1196 = n3229 | n3233 ;
  assign n3513 = ~x2 ;
  assign n1192 = n3513 & x130 ;
  assign n3514 = ~x129 ;
  assign n3227 = x1 & n3514 ;
  assign n3515 = ~x1 ;
  assign n3225 = n3515 & x129 ;
  assign n3516 = ~x128 ;
  assign n1193 = x0 & n3516 ;
  assign n3517 = ~n3225 ;
  assign n1194 = n3517 & n1193 ;
  assign n1195 = n3227 | n1194 ;
  assign n3518 = ~n1192 ;
  assign n1197 = n3518 & n1195 ;
  assign n1198 = n1196 | n1197 ;
  assign n3519 = ~x4 ;
  assign n3235 = n3519 & x132 ;
  assign n3520 = ~x3 ;
  assign n3237 = n3520 & x131 ;
  assign n1199 = n3235 | n3237 ;
  assign n3521 = ~n1199 ;
  assign n1200 = n1198 & n3521 ;
  assign n3522 = ~x133 ;
  assign n1201 = x5 & n3522 ;
  assign n3523 = ~x132 ;
  assign n1202 = x4 & n3523 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = n1200 | n1203 ;
  assign n3524 = ~x6 ;
  assign n1205 = n3524 & x134 ;
  assign n3525 = ~x5 ;
  assign n1206 = n3525 & x133 ;
  assign n1207 = n1205 | n1206 ;
  assign n3526 = ~n1207 ;
  assign n1209 = n1204 & n3526 ;
  assign n1210 = n1208 | n1209 ;
  assign n3527 = ~n1191 ;
  assign n1211 = n3527 & n1210 ;
  assign n1212 = n3243 | n1211 ;
  assign n3528 = ~x8 ;
  assign n3245 = n3528 & x136 ;
  assign n3529 = ~x9 ;
  assign n3247 = n3529 & x137 ;
  assign n1213 = n3245 | n3247 ;
  assign n3530 = ~n1213 ;
  assign n1215 = n1212 & n3530 ;
  assign n1216 = n1214 | n1215 ;
  assign n3531 = ~n1190 ;
  assign n1217 = n3531 & n1216 ;
  assign n3532 = ~x139 ;
  assign n3249 = x11 & n3532 ;
  assign n3533 = ~x138 ;
  assign n3251 = x10 & n3533 ;
  assign n1218 = n3249 | n3251 ;
  assign n1219 = n1217 | n1218 ;
  assign n3534 = ~x11 ;
  assign n3253 = n3534 & x139 ;
  assign n3535 = ~x12 ;
  assign n3255 = n3535 & x140 ;
  assign n1220 = n3253 | n3255 ;
  assign n3536 = ~n1220 ;
  assign n1222 = n1219 & n3536 ;
  assign n1223 = n1221 | n1222 ;
  assign n3537 = ~n1189 ;
  assign n1224 = n3537 & n1223 ;
  assign n3538 = ~x141 ;
  assign n1225 = x13 & n3538 ;
  assign n3539 = ~x142 ;
  assign n1226 = x14 & n3539 ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = n1224 | n1227 ;
  assign n3540 = ~n1188 ;
  assign n1230 = n3540 & n1228 ;
  assign n1231 = n1229 | n1230 ;
  assign n3541 = ~x15 ;
  assign n3257 = n3541 & x143 ;
  assign n3542 = ~x16 ;
  assign n1232 = n3542 & x144 ;
  assign n1233 = n3257 | n1232 ;
  assign n3543 = ~n1233 ;
  assign n1234 = n1231 & n3543 ;
  assign n1235 = n1187 | n1234 ;
  assign n3544 = ~n1186 ;
  assign n1239 = n3544 & n1235 ;
  assign n1240 = n1238 | n1239 ;
  assign n3545 = ~x18 ;
  assign n1241 = n3545 & x146 ;
  assign n3546 = ~x19 ;
  assign n1242 = n3546 & x147 ;
  assign n1243 = n1241 | n1242 ;
  assign n3547 = ~n1243 ;
  assign n1244 = n1240 & n3547 ;
  assign n3548 = ~x148 ;
  assign n1245 = x20 & n3548 ;
  assign n3549 = ~x147 ;
  assign n1246 = x19 & n3549 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = n1244 | n1247 ;
  assign n3550 = ~x21 ;
  assign n3259 = n3550 & x149 ;
  assign n3551 = ~x20 ;
  assign n1249 = n3551 & x148 ;
  assign n1250 = n3259 | n1249 ;
  assign n3552 = ~n1250 ;
  assign n1252 = n1248 & n3552 ;
  assign n1253 = n1251 | n1252 ;
  assign n3553 = ~n1185 ;
  assign n1254 = n3553 & n1253 ;
  assign n3554 = ~x150 ;
  assign n1255 = x22 & n3554 ;
  assign n3555 = ~x151 ;
  assign n1256 = x23 & n3555 ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = n1254 | n1257 ;
  assign n3556 = ~x23 ;
  assign n1259 = n3556 & x151 ;
  assign n3557 = ~x24 ;
  assign n1260 = n3557 & x152 ;
  assign n1261 = n1259 | n1260 ;
  assign n3558 = ~n1261 ;
  assign n1265 = n1258 & n3558 ;
  assign n1266 = n1264 | n1265 ;
  assign n3559 = ~n1184 ;
  assign n1267 = n3559 & n1266 ;
  assign n1268 = n1183 | n1267 ;
  assign n3560 = ~x27 ;
  assign n1269 = n3560 & x155 ;
  assign n3561 = ~x26 ;
  assign n1270 = n3561 & x154 ;
  assign n1271 = n1269 | n1270 ;
  assign n3562 = ~n1271 ;
  assign n1275 = n1268 & n3562 ;
  assign n1276 = n1274 | n1275 ;
  assign n3563 = ~x28 ;
  assign n1277 = n3563 & x156 ;
  assign n3564 = ~x29 ;
  assign n1278 = n3564 & x157 ;
  assign n1279 = n1277 | n1278 ;
  assign n3565 = ~n1279 ;
  assign n1280 = n1276 & n3565 ;
  assign n1281 = n1182 | n1280 ;
  assign n3566 = ~n1181 ;
  assign n1285 = n3566 & n1281 ;
  assign n1286 = n1284 | n1285 ;
  assign n3567 = ~x31 ;
  assign n1287 = n3567 & x159 ;
  assign n3568 = ~x32 ;
  assign n1288 = n3568 & x160 ;
  assign n1289 = n1287 | n1288 ;
  assign n3569 = ~n1289 ;
  assign n1290 = n1286 & n3569 ;
  assign n3570 = ~x161 ;
  assign n1291 = x33 & n3570 ;
  assign n3571 = ~x160 ;
  assign n1292 = x32 & n3571 ;
  assign n1293 = n1291 | n1292 ;
  assign n1294 = n1290 | n1293 ;
  assign n3572 = ~n1180 ;
  assign n1295 = n3572 & n1294 ;
  assign n1296 = n1179 | n1295 ;
  assign n3573 = ~n1178 ;
  assign n1297 = n3573 & n1296 ;
  assign n1298 = n1177 | n1297 ;
  assign n3574 = ~x36 ;
  assign n1299 = n3574 & x164 ;
  assign n3575 = ~x35 ;
  assign n1300 = n3575 & x163 ;
  assign n1301 = n1299 | n1300 ;
  assign n3576 = ~n1301 ;
  assign n1305 = n1298 & n3576 ;
  assign n1306 = n1304 | n1305 ;
  assign n3577 = ~x37 ;
  assign n1307 = n3577 & x165 ;
  assign n3578 = ~x38 ;
  assign n1308 = n3578 & x166 ;
  assign n1309 = n1307 | n1308 ;
  assign n3579 = ~n1309 ;
  assign n1310 = n1306 & n3579 ;
  assign n3580 = ~x167 ;
  assign n3261 = x39 & n3580 ;
  assign n3581 = ~x166 ;
  assign n1311 = x38 & n3581 ;
  assign n1312 = n3261 | n1311 ;
  assign n1313 = n1310 | n1312 ;
  assign n3582 = ~x40 ;
  assign n1314 = n3582 & x168 ;
  assign n1316 = n1314 | n1315 ;
  assign n3583 = ~x39 ;
  assign n1317 = n3583 & x167 ;
  assign n1318 = n1316 | n1317 ;
  assign n3584 = ~n1318 ;
  assign n1325 = n1313 & n3584 ;
  assign n1326 = n1324 | n1325 ;
  assign n3585 = ~x43 ;
  assign n1327 = n3585 & x171 ;
  assign n3586 = ~x42 ;
  assign n1328 = n3586 & x170 ;
  assign n1329 = n1327 | n1328 ;
  assign n3587 = ~n1329 ;
  assign n1330 = n1326 & n3587 ;
  assign n1331 = n1176 | n1330 ;
  assign n3588 = ~n1175 ;
  assign n1335 = n3588 & n1331 ;
  assign n1336 = n1334 | n1335 ;
  assign n3589 = ~x46 ;
  assign n1337 = n3589 & x174 ;
  assign n3590 = ~x45 ;
  assign n1338 = n3590 & x173 ;
  assign n1339 = n1337 | n1338 ;
  assign n3591 = ~n1339 ;
  assign n1340 = n1336 & n3591 ;
  assign n1341 = n1174 | n1340 ;
  assign n3592 = ~n1173 ;
  assign n1345 = n3592 & n1341 ;
  assign n1346 = n1344 | n1345 ;
  assign n3593 = ~n1172 ;
  assign n1347 = n3593 & n1346 ;
  assign n1348 = n1171 | n1347 ;
  assign n3594 = ~x50 ;
  assign n3263 = n3594 & x178 ;
  assign n3595 = ~x49 ;
  assign n1349 = n3595 & x177 ;
  assign n1350 = n3263 | n1349 ;
  assign n3596 = ~n1350 ;
  assign n1352 = n1348 & n3596 ;
  assign n1353 = n1351 | n1352 ;
  assign n3597 = ~n1170 ;
  assign n1354 = n3597 & n1353 ;
  assign n3598 = ~x179 ;
  assign n1355 = x51 & n3598 ;
  assign n3599 = ~x180 ;
  assign n1356 = x52 & n3599 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = n1354 | n1357 ;
  assign n3600 = ~n1169 ;
  assign n1360 = n3600 & n1358 ;
  assign n1361 = n1359 | n1360 ;
  assign n3601 = ~x53 ;
  assign n3265 = n3601 & x181 ;
  assign n3602 = ~x54 ;
  assign n1362 = n3602 & x182 ;
  assign n1363 = n3265 | n1362 ;
  assign n3603 = ~n1363 ;
  assign n1364 = n1361 & n3603 ;
  assign n3604 = ~x183 ;
  assign n1365 = x55 & n3604 ;
  assign n3605 = ~x182 ;
  assign n1366 = x54 & n3605 ;
  assign n1367 = n1365 | n1366 ;
  assign n1368 = n1364 | n1367 ;
  assign n3606 = ~n1168 ;
  assign n1370 = n3606 & n1368 ;
  assign n1371 = n1369 | n1370 ;
  assign n3607 = ~x56 ;
  assign n3267 = n3607 & x184 ;
  assign n3608 = ~x57 ;
  assign n1372 = n3608 & x185 ;
  assign n1373 = n3267 | n1372 ;
  assign n3609 = ~n1373 ;
  assign n1374 = n1371 & n3609 ;
  assign n1375 = n1167 | n1374 ;
  assign n3610 = ~n1166 ;
  assign n1379 = n3610 & n1375 ;
  assign n1380 = n1378 | n1379 ;
  assign n3611 = ~x59 ;
  assign n1381 = n3611 & x187 ;
  assign n3612 = ~x60 ;
  assign n1382 = n3612 & x188 ;
  assign n1383 = n1381 | n1382 ;
  assign n3613 = ~n1383 ;
  assign n1384 = n1380 & n3613 ;
  assign n3614 = ~x189 ;
  assign n1385 = x61 & n3614 ;
  assign n3615 = ~x188 ;
  assign n1386 = x60 & n3615 ;
  assign n1387 = n1385 | n1386 ;
  assign n1388 = n1384 | n1387 ;
  assign n3616 = ~n1165 ;
  assign n1389 = n3616 & n1388 ;
  assign n1390 = n1164 | n1389 ;
  assign n3617 = ~n1163 ;
  assign n1391 = n3617 & n1390 ;
  assign n1392 = n1162 | n1391 ;
  assign n3618 = ~x64 ;
  assign n1393 = n3618 & x192 ;
  assign n3619 = ~x63 ;
  assign n1394 = n3619 & x191 ;
  assign n1395 = n1393 | n1394 ;
  assign n3620 = ~n1395 ;
  assign n1399 = n1392 & n3620 ;
  assign n1400 = n1398 | n1399 ;
  assign n3621 = ~x65 ;
  assign n1401 = n3621 & x193 ;
  assign n3622 = ~x66 ;
  assign n1402 = n3622 & x194 ;
  assign n1403 = n1401 | n1402 ;
  assign n3623 = ~n1403 ;
  assign n1404 = n1400 & n3623 ;
  assign n3624 = ~x195 ;
  assign n3269 = x67 & n3624 ;
  assign n3625 = ~x194 ;
  assign n1405 = x66 & n3625 ;
  assign n1406 = n3269 | n1405 ;
  assign n1407 = n1404 | n1406 ;
  assign n3626 = ~x68 ;
  assign n1408 = n3626 & x196 ;
  assign n1410 = n1408 | n1409 ;
  assign n3627 = ~x67 ;
  assign n1411 = n3627 & x195 ;
  assign n1412 = n1410 | n1411 ;
  assign n3628 = ~n1412 ;
  assign n1419 = n1407 & n3628 ;
  assign n1420 = n1418 | n1419 ;
  assign n3629 = ~x70 ;
  assign n1421 = n3629 & x198 ;
  assign n3630 = ~x71 ;
  assign n1422 = n3630 & x199 ;
  assign n1423 = n1421 | n1422 ;
  assign n3631 = ~n1423 ;
  assign n1424 = n1420 & n3631 ;
  assign n3632 = ~x200 ;
  assign n1425 = x72 & n3632 ;
  assign n3633 = ~x199 ;
  assign n1426 = x71 & n3633 ;
  assign n1427 = n1425 | n1426 ;
  assign n1428 = n1424 | n1427 ;
  assign n3634 = ~x72 ;
  assign n1429 = n3634 & x200 ;
  assign n3635 = ~x73 ;
  assign n1430 = n3635 & x201 ;
  assign n1431 = n1429 | n1430 ;
  assign n3636 = ~n1431 ;
  assign n1435 = n1428 & n3636 ;
  assign n1436 = n1434 | n1435 ;
  assign n3637 = ~n1161 ;
  assign n1437 = n3637 & n1436 ;
  assign n1438 = n1160 | n1437 ;
  assign n3638 = ~x76 ;
  assign n1439 = n3638 & x204 ;
  assign n3639 = ~x75 ;
  assign n1440 = n3639 & x203 ;
  assign n1441 = n1439 | n1440 ;
  assign n3640 = ~n1441 ;
  assign n1445 = n1438 & n3640 ;
  assign n1446 = n1444 | n1445 ;
  assign n3641 = ~n1159 ;
  assign n1447 = n3641 & n1446 ;
  assign n1448 = n1158 | n1447 ;
  assign n3642 = ~x79 ;
  assign n1449 = n3642 & x207 ;
  assign n3643 = ~x78 ;
  assign n1450 = n3643 & x206 ;
  assign n1451 = n1449 | n1450 ;
  assign n3644 = ~n1451 ;
  assign n1455 = n1448 & n3644 ;
  assign n1456 = n1454 | n1455 ;
  assign n3645 = ~n1157 ;
  assign n1457 = n3645 & n1456 ;
  assign n1458 = n1156 | n1457 ;
  assign n3646 = ~x82 ;
  assign n1459 = n3646 & x210 ;
  assign n3647 = ~x81 ;
  assign n1460 = n3647 & x209 ;
  assign n1461 = n1459 | n1460 ;
  assign n3648 = ~n1461 ;
  assign n1465 = n1458 & n3648 ;
  assign n1466 = n1464 | n1465 ;
  assign n3649 = ~n1155 ;
  assign n1467 = n3649 & n1466 ;
  assign n1468 = n1154 | n1467 ;
  assign n3650 = ~x84 ;
  assign n1469 = n3650 & x212 ;
  assign n3651 = ~x85 ;
  assign n1470 = n3651 & x213 ;
  assign n1471 = n1469 | n1470 ;
  assign n3652 = ~n1471 ;
  assign n1475 = n1468 & n3652 ;
  assign n1476 = n1474 | n1475 ;
  assign n3653 = ~n1153 ;
  assign n1477 = n3653 & n1476 ;
  assign n1478 = n1152 | n1477 ;
  assign n3654 = ~x88 ;
  assign n1479 = n3654 & x216 ;
  assign n3655 = ~x87 ;
  assign n1480 = n3655 & x215 ;
  assign n1481 = n1479 | n1480 ;
  assign n3656 = ~n1481 ;
  assign n1485 = n1478 & n3656 ;
  assign n1486 = n1484 | n1485 ;
  assign n3657 = ~x89 ;
  assign n1487 = n3657 & x217 ;
  assign n3658 = ~x90 ;
  assign n1488 = n3658 & x218 ;
  assign n1489 = n1487 | n1488 ;
  assign n3659 = ~n1489 ;
  assign n1490 = n1486 & n3659 ;
  assign n1491 = n1151 | n1490 ;
  assign n3660 = ~n1150 ;
  assign n1495 = n3660 & n1491 ;
  assign n1496 = n1494 | n1495 ;
  assign n3661 = ~x92 ;
  assign n1497 = n3661 & x220 ;
  assign n3662 = ~x93 ;
  assign n1498 = n3662 & x221 ;
  assign n1499 = n1497 | n1498 ;
  assign n3663 = ~n1499 ;
  assign n1500 = n1496 & n3663 ;
  assign n3664 = ~x221 ;
  assign n1501 = x93 & n3664 ;
  assign n3665 = ~x222 ;
  assign n1502 = x94 & n3665 ;
  assign n1503 = n1501 | n1502 ;
  assign n1504 = n1500 | n1503 ;
  assign n3666 = ~x95 ;
  assign n1505 = n3666 & x223 ;
  assign n3667 = ~x94 ;
  assign n1506 = n3667 & x222 ;
  assign n1507 = n1505 | n1506 ;
  assign n3668 = ~n1507 ;
  assign n1511 = n1504 & n3668 ;
  assign n1512 = n1510 | n1511 ;
  assign n3669 = ~n1149 ;
  assign n1513 = n3669 & n1512 ;
  assign n1514 = n1148 | n1513 ;
  assign n3670 = ~x98 ;
  assign n3271 = n3670 & x226 ;
  assign n3671 = ~x97 ;
  assign n1515 = n3671 & x225 ;
  assign n1516 = n3271 | n1515 ;
  assign n3672 = ~n1516 ;
  assign n1518 = n1514 & n3672 ;
  assign n1519 = n1517 | n1518 ;
  assign n3673 = ~n1147 ;
  assign n1520 = n3673 & n1519 ;
  assign n3674 = ~x228 ;
  assign n1521 = x100 & n3674 ;
  assign n3675 = ~x227 ;
  assign n1522 = x99 & n3675 ;
  assign n1523 = n1521 | n1522 ;
  assign n1524 = n1520 | n1523 ;
  assign n3676 = ~x101 ;
  assign n3273 = n3676 & x229 ;
  assign n3677 = ~x100 ;
  assign n1525 = n3677 & x228 ;
  assign n1526 = n3273 | n1525 ;
  assign n3678 = ~n1526 ;
  assign n1528 = n1524 & n3678 ;
  assign n1529 = n1527 | n1528 ;
  assign n3679 = ~n1146 ;
  assign n1530 = n3679 & n1529 ;
  assign n3680 = ~x230 ;
  assign n1531 = x102 & n3680 ;
  assign n3681 = ~x231 ;
  assign n1532 = x103 & n3681 ;
  assign n1533 = n1531 | n1532 ;
  assign n1534 = n1530 | n1533 ;
  assign n3682 = ~x103 ;
  assign n1535 = n3682 & x231 ;
  assign n3683 = ~x104 ;
  assign n1536 = n3683 & x232 ;
  assign n1537 = n1535 | n1536 ;
  assign n3684 = ~n1537 ;
  assign n1541 = n1534 & n3684 ;
  assign n1542 = n1540 | n1541 ;
  assign n3685 = ~x105 ;
  assign n1543 = n3685 & x233 ;
  assign n3686 = ~x106 ;
  assign n1544 = n3686 & x234 ;
  assign n1545 = n1543 | n1544 ;
  assign n3687 = ~n1545 ;
  assign n1546 = n1542 & n3687 ;
  assign n1547 = n1145 | n1546 ;
  assign n3688 = ~n1144 ;
  assign n1551 = n3688 & n1547 ;
  assign n1552 = n1550 | n1551 ;
  assign n3689 = ~x109 ;
  assign n1553 = n3689 & x237 ;
  assign n3690 = ~x108 ;
  assign n1554 = n3690 & x236 ;
  assign n1555 = n1553 | n1554 ;
  assign n3691 = ~n1555 ;
  assign n1556 = n1552 & n3691 ;
  assign n1557 = n1143 | n1556 ;
  assign n3692 = ~n1142 ;
  assign n1561 = n3692 & n1557 ;
  assign n1562 = n1560 | n1561 ;
  assign n3693 = ~n1141 ;
  assign n1563 = n3693 & n1562 ;
  assign n1564 = n1140 | n1563 ;
  assign n3694 = ~x112 ;
  assign n1565 = n3694 & x240 ;
  assign n3695 = ~x113 ;
  assign n1566 = n3695 & x241 ;
  assign n1567 = n1565 | n1566 ;
  assign n3696 = ~n1567 ;
  assign n1571 = n1564 & n3696 ;
  assign n1572 = n1570 | n1571 ;
  assign n3697 = ~n1139 ;
  assign n1573 = n3697 & n1572 ;
  assign n1574 = n1138 | n1573 ;
  assign n3698 = ~x116 ;
  assign n1575 = n3698 & x244 ;
  assign n3699 = ~x115 ;
  assign n1576 = n3699 & x243 ;
  assign n1577 = n1575 | n1576 ;
  assign n3700 = ~n1577 ;
  assign n1581 = n1574 & n3700 ;
  assign n1582 = n1580 | n1581 ;
  assign n3701 = ~x117 ;
  assign n1583 = n3701 & x245 ;
  assign n3702 = ~x118 ;
  assign n1584 = n3702 & x246 ;
  assign n1585 = n1583 | n1584 ;
  assign n3703 = ~n1585 ;
  assign n1586 = n1582 & n3703 ;
  assign n1587 = n1137 | n1586 ;
  assign n3704 = ~n1136 ;
  assign n1588 = n3704 & n1587 ;
  assign n3705 = ~x248 ;
  assign n3275 = x120 & n3705 ;
  assign n3706 = ~x247 ;
  assign n3277 = x119 & n3706 ;
  assign n1589 = n3275 | n3277 ;
  assign n1590 = n1588 | n1589 ;
  assign n3707 = ~x121 ;
  assign n3279 = n3707 & x249 ;
  assign n3708 = ~x120 ;
  assign n3281 = n3708 & x248 ;
  assign n1591 = n3279 | n3281 ;
  assign n3709 = ~n1591 ;
  assign n1592 = n1590 & n3709 ;
  assign n3710 = ~x249 ;
  assign n3283 = x121 & n3710 ;
  assign n3711 = ~x250 ;
  assign n3285 = x122 & n3711 ;
  assign n1593 = n3283 | n3285 ;
  assign n1595 = n1592 | n1593 ;
  assign n3712 = ~n1594 ;
  assign n1596 = n3712 & n1595 ;
  assign n1597 = n1135 | n1596 ;
  assign n3713 = ~x124 ;
  assign n3287 = n3713 & x252 ;
  assign n3714 = ~x123 ;
  assign n3289 = n3714 & x251 ;
  assign n1598 = n3287 | n3289 ;
  assign n3715 = ~n1598 ;
  assign n1599 = n1597 & n3715 ;
  assign n3716 = ~x253 ;
  assign n3291 = x125 & n3716 ;
  assign n3717 = ~x252 ;
  assign n3293 = x124 & n3717 ;
  assign n1600 = n3291 | n3293 ;
  assign n1602 = n1599 | n1600 ;
  assign n3718 = ~n1601 ;
  assign n1603 = n3718 & n1602 ;
  assign n3719 = ~x127 ;
  assign n3299 = n3719 & x255 ;
  assign n3720 = ~x254 ;
  assign n3301 = x126 & n3720 ;
  assign n1604 = n3299 | n3301 ;
  assign n1605 = n1603 | n1604 ;
  assign n3721 = ~n1134 ;
  assign n1606 = n3721 & n1605 ;
  assign n1674 = x0 & n1606 ;
  assign n3722 = ~n1606 ;
  assign n2906 = x128 & n3722 ;
  assign n2907 = n1674 | n2906 ;
  assign n3129 = x127 & x255 ;
  assign n3131 = x383 & x511 ;
  assign n3723 = ~n3129 ;
  assign n3303 = n3723 & n3131 ;
  assign n3724 = ~x383 ;
  assign n3305 = n3724 & x511 ;
  assign n3725 = ~x510 ;
  assign n3217 = x382 & n3725 ;
  assign n3726 = ~x509 ;
  assign n3219 = x381 & n3726 ;
  assign n1060 = n3217 | n3219 ;
  assign n3727 = ~x379 ;
  assign n3307 = n3727 & x507 ;
  assign n3728 = ~x506 ;
  assign n1053 = x378 & n3728 ;
  assign n3729 = ~x503 ;
  assign n3309 = x375 & n3729 ;
  assign n3730 = ~x374 ;
  assign n3311 = n3730 & x502 ;
  assign n3731 = ~x372 ;
  assign n1037 = n3731 & x500 ;
  assign n3732 = ~x373 ;
  assign n1038 = n3732 & x501 ;
  assign n1039 = n1037 | n1038 ;
  assign n3733 = ~x371 ;
  assign n3313 = n3733 & x499 ;
  assign n3734 = ~x498 ;
  assign n3315 = x370 & n3734 ;
  assign n3735 = ~x369 ;
  assign n1027 = n3735 & x497 ;
  assign n3736 = ~x370 ;
  assign n1028 = n3736 & x498 ;
  assign n1029 = n1027 | n1028 ;
  assign n3737 = ~x368 ;
  assign n3317 = n3737 & x496 ;
  assign n3738 = ~x495 ;
  assign n3319 = x367 & n3738 ;
  assign n3739 = ~x366 ;
  assign n1017 = n3739 & x494 ;
  assign n3740 = ~x367 ;
  assign n1018 = n3740 & x495 ;
  assign n1019 = n1017 | n1018 ;
  assign n3741 = ~x494 ;
  assign n3321 = x366 & n3741 ;
  assign n3742 = ~x365 ;
  assign n3323 = n3742 & x493 ;
  assign n3743 = ~x364 ;
  assign n1007 = n3743 & x492 ;
  assign n3744 = ~x363 ;
  assign n1008 = n3744 & x491 ;
  assign n1009 = n1007 | n1008 ;
  assign n3745 = ~x491 ;
  assign n3325 = x363 & n3745 ;
  assign n3746 = ~x362 ;
  assign n3327 = n3746 & x490 ;
  assign n3747 = ~x361 ;
  assign n997 = n3747 & x489 ;
  assign n3748 = ~x360 ;
  assign n998 = n3748 & x488 ;
  assign n999 = n997 | n998 ;
  assign n3749 = ~x486 ;
  assign n3329 = x358 & n3749 ;
  assign n3750 = ~x357 ;
  assign n986 = n3750 & x485 ;
  assign n3751 = ~x483 ;
  assign n3331 = x355 & n3751 ;
  assign n3752 = ~x354 ;
  assign n976 = n3752 & x482 ;
  assign n3753 = ~x353 ;
  assign n3333 = n3753 & x481 ;
  assign n3754 = ~x480 ;
  assign n3335 = x352 & n3754 ;
  assign n3755 = ~x351 ;
  assign n967 = n3755 & x479 ;
  assign n3756 = ~x352 ;
  assign n968 = n3756 & x480 ;
  assign n969 = n967 | n968 ;
  assign n3757 = ~x348 ;
  assign n954 = n3757 & x476 ;
  assign n3758 = ~x475 ;
  assign n3337 = x347 & n3758 ;
  assign n3759 = ~x344 ;
  assign n941 = n3759 & x472 ;
  assign n3760 = ~x345 ;
  assign n942 = n3760 & x473 ;
  assign n943 = n941 | n942 ;
  assign n3761 = ~x340 ;
  assign n924 = n3761 & x468 ;
  assign n3762 = ~x467 ;
  assign n3339 = x339 & n3762 ;
  assign n3763 = ~x339 ;
  assign n3341 = n3763 & x467 ;
  assign n3764 = ~x466 ;
  assign n3343 = x338 & n3764 ;
  assign n3765 = ~x338 ;
  assign n3345 = n3765 & x466 ;
  assign n3766 = ~x465 ;
  assign n3347 = x337 & n3766 ;
  assign n3767 = ~x337 ;
  assign n3349 = n3767 & x465 ;
  assign n3768 = ~x464 ;
  assign n3351 = x336 & n3768 ;
  assign n3769 = ~x336 ;
  assign n3353 = n3769 & x464 ;
  assign n3770 = ~x463 ;
  assign n3355 = x335 & n3770 ;
  assign n3771 = ~x335 ;
  assign n3357 = n3771 & x463 ;
  assign n3772 = ~x462 ;
  assign n3359 = x334 & n3772 ;
  assign n3773 = ~x334 ;
  assign n3361 = n3773 & x462 ;
  assign n3774 = ~x461 ;
  assign n3363 = x333 & n3774 ;
  assign n3775 = ~x333 ;
  assign n3365 = n3775 & x461 ;
  assign n3776 = ~x460 ;
  assign n3367 = x332 & n3776 ;
  assign n3777 = ~x332 ;
  assign n905 = n3777 & x460 ;
  assign n3778 = ~x331 ;
  assign n906 = n3778 & x459 ;
  assign n907 = n905 | n906 ;
  assign n3779 = ~x457 ;
  assign n3369 = x329 & n3779 ;
  assign n3780 = ~x328 ;
  assign n894 = n3780 & x456 ;
  assign n3781 = ~x454 ;
  assign n3371 = x326 & n3781 ;
  assign n3782 = ~x325 ;
  assign n884 = n3782 & x453 ;
  assign n3783 = ~x451 ;
  assign n3373 = x323 & n3783 ;
  assign n3784 = ~x322 ;
  assign n874 = n3784 & x450 ;
  assign n3785 = ~x319 ;
  assign n862 = n3785 & x447 ;
  assign n3786 = ~x446 ;
  assign n3375 = x318 & n3786 ;
  assign n3787 = ~x316 ;
  assign n849 = n3787 & x444 ;
  assign n3788 = ~x315 ;
  assign n850 = n3788 & x443 ;
  assign n851 = n849 | n850 ;
  assign n3789 = ~x443 ;
  assign n3377 = x315 & n3789 ;
  assign n3790 = ~x314 ;
  assign n3379 = n3790 & x442 ;
  assign n3791 = ~x312 ;
  assign n839 = n3791 & x440 ;
  assign n3792 = ~x313 ;
  assign n840 = n3792 & x441 ;
  assign n841 = n839 | n840 ;
  assign n3793 = ~x440 ;
  assign n3381 = x312 & n3793 ;
  assign n3794 = ~x311 ;
  assign n3383 = n3794 & x439 ;
  assign n3795 = ~x310 ;
  assign n829 = n3795 & x438 ;
  assign n3796 = ~x309 ;
  assign n830 = n3796 & x437 ;
  assign n831 = n829 | n830 ;
  assign n3797 = ~x437 ;
  assign n4416 = x309 & n3797 ;
  assign n3798 = ~x308 ;
  assign n4418 = n3798 & x436 ;
  assign n3799 = ~x307 ;
  assign n819 = n3799 & x435 ;
  assign n3800 = ~x306 ;
  assign n820 = n3800 & x434 ;
  assign n821 = n819 | n820 ;
  assign n3801 = ~x302 ;
  assign n803 = n3801 & x430 ;
  assign n3802 = ~x303 ;
  assign n804 = n3802 & x431 ;
  assign n805 = n803 | n804 ;
  assign n3803 = ~x297 ;
  assign n783 = n3803 & x425 ;
  assign n3804 = ~x298 ;
  assign n784 = n3804 & x426 ;
  assign n785 = n783 | n784 ;
  assign n3805 = ~x423 ;
  assign n643 = x295 & n3805 ;
  assign n3806 = ~x294 ;
  assign n644 = n3806 & x422 ;
  assign n3807 = ~x422 ;
  assign n645 = x294 & n3807 ;
  assign n3808 = ~x293 ;
  assign n646 = n3808 & x421 ;
  assign n3809 = ~x291 ;
  assign n763 = n3809 & x419 ;
  assign n3810 = ~x292 ;
  assign n764 = n3810 & x420 ;
  assign n765 = n763 | n764 ;
  assign n3811 = ~x290 ;
  assign n647 = n3811 & x418 ;
  assign n3812 = ~x288 ;
  assign n752 = n3812 & x416 ;
  assign n3813 = ~x289 ;
  assign n753 = n3813 & x417 ;
  assign n754 = n752 | n753 ;
  assign n3814 = ~x416 ;
  assign n648 = x288 & n3814 ;
  assign n3815 = ~x286 ;
  assign n741 = n3815 & x414 ;
  assign n3816 = ~x285 ;
  assign n742 = n3816 & x413 ;
  assign n743 = n741 | n742 ;
  assign n3817 = ~x413 ;
  assign n649 = x285 & n3817 ;
  assign n3818 = ~x284 ;
  assign n650 = n3818 & x412 ;
  assign n3819 = ~x283 ;
  assign n734 = n3819 & x411 ;
  assign n3820 = ~x410 ;
  assign n651 = x282 & n3820 ;
  assign n3821 = ~x409 ;
  assign n652 = x281 & n3821 ;
  assign n3822 = ~x280 ;
  assign n726 = n3822 & x408 ;
  assign n3823 = ~x277 ;
  assign n714 = n3823 & x405 ;
  assign n3824 = ~x404 ;
  assign n653 = x276 & n3824 ;
  assign n3825 = ~x274 ;
  assign n704 = n3825 & x402 ;
  assign n3826 = ~x271 ;
  assign n693 = n3826 & x399 ;
  assign n3827 = ~x398 ;
  assign n654 = x270 & n3827 ;
  assign n3828 = ~x267 ;
  assign n3165 = n3828 & x395 ;
  assign n3829 = ~x268 ;
  assign n681 = n3829 & x396 ;
  assign n682 = n3165 | n681 ;
  assign n3830 = ~x395 ;
  assign n655 = x267 & n3830 ;
  assign n3831 = ~x266 ;
  assign n3163 = n3831 & x394 ;
  assign n3832 = ~x265 ;
  assign n3155 = n3832 & x393 ;
  assign n3833 = ~x264 ;
  assign n3157 = n3833 & x392 ;
  assign n675 = n3155 | n3157 ;
  assign n3834 = ~x392 ;
  assign n656 = x264 & n3834 ;
  assign n3835 = ~x263 ;
  assign n3153 = n3835 & x391 ;
  assign n3836 = ~x262 ;
  assign n3145 = n3836 & x390 ;
  assign n3837 = ~x261 ;
  assign n3147 = n3837 & x389 ;
  assign n669 = n3145 | n3147 ;
  assign n3838 = ~x389 ;
  assign n657 = x261 & n3838 ;
  assign n3839 = ~x260 ;
  assign n3143 = n3839 & x388 ;
  assign n3840 = ~x259 ;
  assign n3135 = n3840 & x387 ;
  assign n3841 = ~x258 ;
  assign n3137 = n3841 & x386 ;
  assign n663 = n3135 | n3137 ;
  assign n3842 = ~x257 ;
  assign n3133 = n3842 & x385 ;
  assign n3843 = ~x384 ;
  assign n658 = x256 & n3843 ;
  assign n3844 = ~n3133 ;
  assign n659 = n3844 & n658 ;
  assign n3845 = ~x386 ;
  assign n660 = x258 & n3845 ;
  assign n3846 = ~x385 ;
  assign n661 = x257 & n3846 ;
  assign n662 = n660 | n661 ;
  assign n664 = n659 | n662 ;
  assign n3847 = ~n663 ;
  assign n665 = n3847 & n664 ;
  assign n3848 = ~x388 ;
  assign n3139 = x260 & n3848 ;
  assign n3849 = ~x387 ;
  assign n3141 = x259 & n3849 ;
  assign n666 = n3139 | n3141 ;
  assign n667 = n665 | n666 ;
  assign n3850 = ~n3143 ;
  assign n668 = n3850 & n667 ;
  assign n670 = n657 | n668 ;
  assign n3851 = ~n669 ;
  assign n671 = n3851 & n670 ;
  assign n3852 = ~x391 ;
  assign n3149 = x263 & n3852 ;
  assign n3853 = ~x390 ;
  assign n3151 = x262 & n3853 ;
  assign n672 = n3149 | n3151 ;
  assign n673 = n671 | n672 ;
  assign n3854 = ~n3153 ;
  assign n674 = n3854 & n673 ;
  assign n676 = n656 | n674 ;
  assign n3855 = ~n675 ;
  assign n677 = n3855 & n676 ;
  assign n3856 = ~x393 ;
  assign n3159 = x265 & n3856 ;
  assign n3857 = ~x394 ;
  assign n3161 = x266 & n3857 ;
  assign n678 = n3159 | n3161 ;
  assign n679 = n677 | n678 ;
  assign n3858 = ~n3163 ;
  assign n680 = n3858 & n679 ;
  assign n683 = n655 | n680 ;
  assign n3859 = ~n682 ;
  assign n684 = n3859 & n683 ;
  assign n3860 = ~x396 ;
  assign n685 = x268 & n3860 ;
  assign n3861 = ~x397 ;
  assign n686 = x269 & n3861 ;
  assign n687 = n685 | n686 ;
  assign n688 = n684 | n687 ;
  assign n3862 = ~x270 ;
  assign n689 = n3862 & x398 ;
  assign n3863 = ~x269 ;
  assign n690 = n3863 & x397 ;
  assign n691 = n689 | n690 ;
  assign n3864 = ~n691 ;
  assign n692 = n688 & n3864 ;
  assign n694 = n654 | n692 ;
  assign n3865 = ~n693 ;
  assign n695 = n3865 & n694 ;
  assign n3866 = ~x399 ;
  assign n3167 = x271 & n3866 ;
  assign n3867 = ~x400 ;
  assign n696 = x272 & n3867 ;
  assign n697 = n3167 | n696 ;
  assign n698 = n695 | n697 ;
  assign n3868 = ~x273 ;
  assign n699 = n3868 & x401 ;
  assign n3869 = ~x272 ;
  assign n700 = n3869 & x400 ;
  assign n701 = n699 | n700 ;
  assign n3870 = ~n701 ;
  assign n702 = n698 & n3870 ;
  assign n3871 = ~x401 ;
  assign n703 = x273 & n3871 ;
  assign n705 = n702 | n703 ;
  assign n3872 = ~n704 ;
  assign n706 = n3872 & n705 ;
  assign n3873 = ~x402 ;
  assign n3169 = x274 & n3873 ;
  assign n3874 = ~x403 ;
  assign n707 = x275 & n3874 ;
  assign n708 = n3169 | n707 ;
  assign n709 = n706 | n708 ;
  assign n3875 = ~x275 ;
  assign n710 = n3875 & x403 ;
  assign n3876 = ~x276 ;
  assign n711 = n3876 & x404 ;
  assign n712 = n710 | n711 ;
  assign n3877 = ~n712 ;
  assign n713 = n709 & n3877 ;
  assign n715 = n653 | n713 ;
  assign n3878 = ~n714 ;
  assign n716 = n3878 & n715 ;
  assign n3879 = ~x405 ;
  assign n3171 = x277 & n3879 ;
  assign n3880 = ~x406 ;
  assign n717 = x278 & n3880 ;
  assign n718 = n3171 | n717 ;
  assign n719 = n716 | n718 ;
  assign n3881 = ~x278 ;
  assign n720 = n3881 & x406 ;
  assign n3882 = ~x279 ;
  assign n721 = n3882 & x407 ;
  assign n722 = n720 | n721 ;
  assign n3883 = ~n722 ;
  assign n723 = n719 & n3883 ;
  assign n3884 = ~x408 ;
  assign n3173 = x280 & n3884 ;
  assign n3885 = ~x407 ;
  assign n724 = x279 & n3885 ;
  assign n725 = n3173 | n724 ;
  assign n727 = n723 | n725 ;
  assign n3886 = ~n726 ;
  assign n728 = n3886 & n727 ;
  assign n729 = n652 | n728 ;
  assign n3887 = ~x281 ;
  assign n730 = n3887 & x409 ;
  assign n3888 = ~x282 ;
  assign n731 = n3888 & x410 ;
  assign n732 = n730 | n731 ;
  assign n3889 = ~n732 ;
  assign n733 = n729 & n3889 ;
  assign n735 = n651 | n733 ;
  assign n3890 = ~n734 ;
  assign n736 = n3890 & n735 ;
  assign n3891 = ~x411 ;
  assign n3175 = x283 & n3891 ;
  assign n3892 = ~x412 ;
  assign n737 = x284 & n3892 ;
  assign n738 = n3175 | n737 ;
  assign n739 = n736 | n738 ;
  assign n3893 = ~n650 ;
  assign n740 = n3893 & n739 ;
  assign n744 = n649 | n740 ;
  assign n3894 = ~n743 ;
  assign n745 = n3894 & n744 ;
  assign n3895 = ~x415 ;
  assign n746 = x287 & n3895 ;
  assign n3896 = ~x414 ;
  assign n747 = x286 & n3896 ;
  assign n748 = n746 | n747 ;
  assign n749 = n745 | n748 ;
  assign n3897 = ~x287 ;
  assign n750 = n3897 & x415 ;
  assign n3898 = ~n750 ;
  assign n751 = n749 & n3898 ;
  assign n755 = n648 | n751 ;
  assign n3899 = ~n754 ;
  assign n756 = n3899 & n755 ;
  assign n3900 = ~x417 ;
  assign n757 = x289 & n3900 ;
  assign n758 = n756 | n757 ;
  assign n3901 = ~n647 ;
  assign n759 = n3901 & n758 ;
  assign n3902 = ~x418 ;
  assign n760 = x290 & n3902 ;
  assign n3903 = ~x419 ;
  assign n761 = x291 & n3903 ;
  assign n762 = n760 | n761 ;
  assign n766 = n759 | n762 ;
  assign n3904 = ~n765 ;
  assign n767 = n3904 & n766 ;
  assign n3905 = ~x421 ;
  assign n768 = x293 & n3905 ;
  assign n3906 = ~x420 ;
  assign n769 = x292 & n3906 ;
  assign n770 = n768 | n769 ;
  assign n771 = n767 | n770 ;
  assign n3907 = ~n646 ;
  assign n772 = n3907 & n771 ;
  assign n773 = n645 | n772 ;
  assign n3908 = ~n644 ;
  assign n774 = n3908 & n773 ;
  assign n775 = n643 | n774 ;
  assign n3909 = ~x296 ;
  assign n776 = n3909 & x424 ;
  assign n3910 = ~x295 ;
  assign n777 = n3910 & x423 ;
  assign n778 = n776 | n777 ;
  assign n3911 = ~n778 ;
  assign n779 = n775 & n3911 ;
  assign n3912 = ~x425 ;
  assign n780 = x297 & n3912 ;
  assign n3913 = ~x424 ;
  assign n781 = x296 & n3913 ;
  assign n782 = n780 | n781 ;
  assign n786 = n779 | n782 ;
  assign n3914 = ~n785 ;
  assign n787 = n3914 & n786 ;
  assign n3915 = ~x427 ;
  assign n3177 = x299 & n3915 ;
  assign n3916 = ~x426 ;
  assign n788 = x298 & n3916 ;
  assign n789 = n3177 | n788 ;
  assign n790 = n787 | n789 ;
  assign n3917 = ~x300 ;
  assign n791 = n3917 & x428 ;
  assign n3918 = ~x301 ;
  assign n792 = n3918 & x429 ;
  assign n793 = n791 | n792 ;
  assign n3919 = ~x299 ;
  assign n794 = n3919 & x427 ;
  assign n795 = n793 | n794 ;
  assign n3920 = ~n795 ;
  assign n796 = n790 & n3920 ;
  assign n3921 = ~x428 ;
  assign n797 = x300 & n3921 ;
  assign n3922 = ~n792 ;
  assign n798 = n3922 & n797 ;
  assign n3923 = ~x429 ;
  assign n799 = x301 & n3923 ;
  assign n3924 = ~x430 ;
  assign n800 = x302 & n3924 ;
  assign n801 = n799 | n800 ;
  assign n802 = n798 | n801 ;
  assign n806 = n796 | n802 ;
  assign n3925 = ~n805 ;
  assign n807 = n3925 & n806 ;
  assign n3926 = ~x432 ;
  assign n808 = x304 & n3926 ;
  assign n3927 = ~x431 ;
  assign n809 = x303 & n3927 ;
  assign n810 = n808 | n809 ;
  assign n811 = n807 | n810 ;
  assign n3928 = ~x304 ;
  assign n812 = n3928 & x432 ;
  assign n3929 = ~x305 ;
  assign n813 = n3929 & x433 ;
  assign n814 = n812 | n813 ;
  assign n3930 = ~n814 ;
  assign n815 = n811 & n3930 ;
  assign n3931 = ~x433 ;
  assign n816 = x305 & n3931 ;
  assign n3932 = ~x434 ;
  assign n817 = x306 & n3932 ;
  assign n818 = n816 | n817 ;
  assign n822 = n815 | n818 ;
  assign n3933 = ~n821 ;
  assign n823 = n3933 & n822 ;
  assign n3934 = ~x435 ;
  assign n824 = x307 & n3934 ;
  assign n3935 = ~x436 ;
  assign n825 = x308 & n3935 ;
  assign n826 = n824 | n825 ;
  assign n827 = n823 | n826 ;
  assign n3936 = ~n4418 ;
  assign n828 = n3936 & n827 ;
  assign n832 = n4416 | n828 ;
  assign n3937 = ~n831 ;
  assign n833 = n3937 & n832 ;
  assign n3938 = ~x439 ;
  assign n834 = x311 & n3938 ;
  assign n3939 = ~x438 ;
  assign n835 = x310 & n3939 ;
  assign n836 = n834 | n835 ;
  assign n837 = n833 | n836 ;
  assign n3940 = ~n3383 ;
  assign n838 = n3940 & n837 ;
  assign n842 = n3381 | n838 ;
  assign n3941 = ~n841 ;
  assign n843 = n3941 & n842 ;
  assign n3942 = ~x441 ;
  assign n844 = x313 & n3942 ;
  assign n3943 = ~x442 ;
  assign n845 = x314 & n3943 ;
  assign n846 = n844 | n845 ;
  assign n847 = n843 | n846 ;
  assign n3944 = ~n3379 ;
  assign n848 = n3944 & n847 ;
  assign n852 = n3377 | n848 ;
  assign n3945 = ~n851 ;
  assign n853 = n3945 & n852 ;
  assign n3946 = ~x444 ;
  assign n854 = x316 & n3946 ;
  assign n3947 = ~x445 ;
  assign n855 = x317 & n3947 ;
  assign n856 = n854 | n855 ;
  assign n857 = n853 | n856 ;
  assign n3948 = ~x317 ;
  assign n858 = n3948 & x445 ;
  assign n3949 = ~x318 ;
  assign n859 = n3949 & x446 ;
  assign n860 = n858 | n859 ;
  assign n3950 = ~n860 ;
  assign n861 = n857 & n3950 ;
  assign n863 = n3375 | n861 ;
  assign n3951 = ~n862 ;
  assign n864 = n3951 & n863 ;
  assign n3952 = ~x447 ;
  assign n3179 = x319 & n3952 ;
  assign n3953 = ~x448 ;
  assign n865 = x320 & n3953 ;
  assign n866 = n3179 | n865 ;
  assign n867 = n864 | n866 ;
  assign n3954 = ~x320 ;
  assign n868 = n3954 & x448 ;
  assign n3955 = ~x321 ;
  assign n869 = n3955 & x449 ;
  assign n870 = n868 | n869 ;
  assign n3956 = ~n870 ;
  assign n871 = n867 & n3956 ;
  assign n3957 = ~x450 ;
  assign n3181 = x322 & n3957 ;
  assign n3958 = ~x449 ;
  assign n872 = x321 & n3958 ;
  assign n873 = n3181 | n872 ;
  assign n875 = n871 | n873 ;
  assign n3959 = ~n874 ;
  assign n876 = n3959 & n875 ;
  assign n877 = n3373 | n876 ;
  assign n3960 = ~x324 ;
  assign n878 = n3960 & x452 ;
  assign n3961 = ~x323 ;
  assign n879 = n3961 & x451 ;
  assign n880 = n878 | n879 ;
  assign n3962 = ~n880 ;
  assign n881 = n877 & n3962 ;
  assign n3963 = ~x453 ;
  assign n3183 = x325 & n3963 ;
  assign n3964 = ~x452 ;
  assign n882 = x324 & n3964 ;
  assign n883 = n3183 | n882 ;
  assign n885 = n881 | n883 ;
  assign n3965 = ~n884 ;
  assign n886 = n3965 & n885 ;
  assign n887 = n3371 | n886 ;
  assign n3966 = ~x327 ;
  assign n888 = n3966 & x455 ;
  assign n3967 = ~x326 ;
  assign n889 = n3967 & x454 ;
  assign n890 = n888 | n889 ;
  assign n3968 = ~n890 ;
  assign n891 = n887 & n3968 ;
  assign n3969 = ~x456 ;
  assign n3185 = x328 & n3969 ;
  assign n3970 = ~x455 ;
  assign n892 = x327 & n3970 ;
  assign n893 = n3185 | n892 ;
  assign n895 = n891 | n893 ;
  assign n3971 = ~n894 ;
  assign n896 = n3971 & n895 ;
  assign n897 = n3369 | n896 ;
  assign n3972 = ~x329 ;
  assign n898 = n3972 & x457 ;
  assign n3973 = ~x330 ;
  assign n899 = n3973 & x458 ;
  assign n900 = n898 | n899 ;
  assign n3974 = ~n900 ;
  assign n901 = n897 & n3974 ;
  assign n3975 = ~x458 ;
  assign n902 = x330 & n3975 ;
  assign n3976 = ~x459 ;
  assign n903 = x331 & n3976 ;
  assign n904 = n902 | n903 ;
  assign n908 = n901 | n904 ;
  assign n3977 = ~n907 ;
  assign n909 = n3977 & n908 ;
  assign n910 = n3367 | n909 ;
  assign n3978 = ~n3365 ;
  assign n911 = n3978 & n910 ;
  assign n912 = n3363 | n911 ;
  assign n3979 = ~n3361 ;
  assign n913 = n3979 & n912 ;
  assign n914 = n3359 | n913 ;
  assign n3980 = ~n3357 ;
  assign n915 = n3980 & n914 ;
  assign n916 = n3355 | n915 ;
  assign n3981 = ~n3353 ;
  assign n917 = n3981 & n916 ;
  assign n918 = n3351 | n917 ;
  assign n3982 = ~n3349 ;
  assign n919 = n3982 & n918 ;
  assign n920 = n3347 | n919 ;
  assign n3983 = ~n3345 ;
  assign n921 = n3983 & n920 ;
  assign n922 = n3343 | n921 ;
  assign n3984 = ~n3341 ;
  assign n923 = n3984 & n922 ;
  assign n925 = n3339 | n923 ;
  assign n3985 = ~n924 ;
  assign n926 = n3985 & n925 ;
  assign n3986 = ~x469 ;
  assign n3187 = x341 & n3986 ;
  assign n3987 = ~x468 ;
  assign n3189 = x340 & n3987 ;
  assign n927 = n3187 | n3189 ;
  assign n928 = n926 | n927 ;
  assign n3988 = ~x342 ;
  assign n929 = n3988 & x470 ;
  assign n3989 = ~x343 ;
  assign n930 = n3989 & x471 ;
  assign n931 = n929 | n930 ;
  assign n3990 = ~x341 ;
  assign n932 = n3990 & x469 ;
  assign n933 = n931 | n932 ;
  assign n3991 = ~n933 ;
  assign n934 = n928 & n3991 ;
  assign n3992 = ~x470 ;
  assign n935 = x342 & n3992 ;
  assign n3993 = ~n930 ;
  assign n936 = n3993 & n935 ;
  assign n3994 = ~x471 ;
  assign n937 = x343 & n3994 ;
  assign n3995 = ~x472 ;
  assign n938 = x344 & n3995 ;
  assign n939 = n937 | n938 ;
  assign n940 = n936 | n939 ;
  assign n944 = n934 | n940 ;
  assign n3996 = ~n943 ;
  assign n945 = n3996 & n944 ;
  assign n3997 = ~x474 ;
  assign n946 = x346 & n3997 ;
  assign n3998 = ~x473 ;
  assign n947 = x345 & n3998 ;
  assign n948 = n946 | n947 ;
  assign n949 = n945 | n948 ;
  assign n3999 = ~x346 ;
  assign n950 = n3999 & x474 ;
  assign n4000 = ~x347 ;
  assign n951 = n4000 & x475 ;
  assign n952 = n950 | n951 ;
  assign n4001 = ~n952 ;
  assign n953 = n949 & n4001 ;
  assign n955 = n3337 | n953 ;
  assign n4002 = ~n954 ;
  assign n956 = n4002 & n955 ;
  assign n4003 = ~x476 ;
  assign n3191 = x348 & n4003 ;
  assign n4004 = ~x477 ;
  assign n957 = x349 & n4004 ;
  assign n958 = n3191 | n957 ;
  assign n959 = n956 | n958 ;
  assign n4005 = ~x349 ;
  assign n960 = n4005 & x477 ;
  assign n4006 = ~x350 ;
  assign n961 = n4006 & x478 ;
  assign n962 = n960 | n961 ;
  assign n4007 = ~n962 ;
  assign n963 = n959 & n4007 ;
  assign n4008 = ~x479 ;
  assign n964 = x351 & n4008 ;
  assign n4009 = ~x478 ;
  assign n965 = x350 & n4009 ;
  assign n966 = n964 | n965 ;
  assign n970 = n963 | n966 ;
  assign n4010 = ~n969 ;
  assign n971 = n4010 & n970 ;
  assign n972 = n3335 | n971 ;
  assign n4011 = ~n3333 ;
  assign n973 = n4011 & n972 ;
  assign n4012 = ~x482 ;
  assign n3193 = x354 & n4012 ;
  assign n4013 = ~x481 ;
  assign n974 = x353 & n4013 ;
  assign n975 = n3193 | n974 ;
  assign n977 = n973 | n975 ;
  assign n4014 = ~n976 ;
  assign n978 = n4014 & n977 ;
  assign n979 = n3331 | n978 ;
  assign n4015 = ~x356 ;
  assign n980 = n4015 & x484 ;
  assign n4016 = ~x355 ;
  assign n981 = n4016 & x483 ;
  assign n982 = n980 | n981 ;
  assign n4017 = ~n982 ;
  assign n983 = n979 & n4017 ;
  assign n4018 = ~x485 ;
  assign n3195 = x357 & n4018 ;
  assign n4019 = ~x484 ;
  assign n984 = x356 & n4019 ;
  assign n985 = n3195 | n984 ;
  assign n987 = n983 | n985 ;
  assign n4020 = ~n986 ;
  assign n988 = n4020 & n987 ;
  assign n989 = n3329 | n988 ;
  assign n4021 = ~x358 ;
  assign n990 = n4021 & x486 ;
  assign n4022 = ~x359 ;
  assign n991 = n4022 & x487 ;
  assign n992 = n990 | n991 ;
  assign n4023 = ~n992 ;
  assign n993 = n989 & n4023 ;
  assign n4024 = ~x487 ;
  assign n994 = x359 & n4024 ;
  assign n4025 = ~x488 ;
  assign n995 = x360 & n4025 ;
  assign n996 = n994 | n995 ;
  assign n1000 = n993 | n996 ;
  assign n4026 = ~n999 ;
  assign n1001 = n4026 & n1000 ;
  assign n4027 = ~x489 ;
  assign n1002 = x361 & n4027 ;
  assign n4028 = ~x490 ;
  assign n1003 = x362 & n4028 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = n1001 | n1004 ;
  assign n4029 = ~n3327 ;
  assign n1006 = n4029 & n1005 ;
  assign n1010 = n3325 | n1006 ;
  assign n4030 = ~n1009 ;
  assign n1011 = n4030 & n1010 ;
  assign n4031 = ~x493 ;
  assign n1012 = x365 & n4031 ;
  assign n4032 = ~x492 ;
  assign n1013 = x364 & n4032 ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = n1011 | n1014 ;
  assign n4033 = ~n3323 ;
  assign n1016 = n4033 & n1015 ;
  assign n1020 = n3321 | n1016 ;
  assign n4034 = ~n1019 ;
  assign n1021 = n4034 & n1020 ;
  assign n1022 = n3319 | n1021 ;
  assign n4035 = ~n3317 ;
  assign n1023 = n4035 & n1022 ;
  assign n4036 = ~x496 ;
  assign n1024 = x368 & n4036 ;
  assign n4037 = ~x497 ;
  assign n1025 = x369 & n4037 ;
  assign n1026 = n1024 | n1025 ;
  assign n1030 = n1023 | n1026 ;
  assign n4038 = ~n1029 ;
  assign n1031 = n4038 & n1030 ;
  assign n1032 = n3315 | n1031 ;
  assign n4039 = ~n3313 ;
  assign n1033 = n4039 & n1032 ;
  assign n4040 = ~x500 ;
  assign n1034 = x372 & n4040 ;
  assign n4041 = ~x499 ;
  assign n1035 = x371 & n4041 ;
  assign n1036 = n1034 | n1035 ;
  assign n1040 = n1033 | n1036 ;
  assign n4042 = ~n1039 ;
  assign n1041 = n4042 & n1040 ;
  assign n4043 = ~x501 ;
  assign n1042 = x373 & n4043 ;
  assign n4044 = ~x502 ;
  assign n1043 = x374 & n4044 ;
  assign n1044 = n1042 | n1043 ;
  assign n1045 = n1041 | n1044 ;
  assign n4045 = ~n3311 ;
  assign n1046 = n4045 & n1045 ;
  assign n1047 = n3309 | n1046 ;
  assign n4046 = ~x376 ;
  assign n3197 = n4046 & x504 ;
  assign n4047 = ~x375 ;
  assign n3199 = n4047 & x503 ;
  assign n1048 = n3197 | n3199 ;
  assign n4048 = ~n1048 ;
  assign n1049 = n1047 & n4048 ;
  assign n4049 = ~x505 ;
  assign n3201 = x377 & n4049 ;
  assign n4050 = ~x504 ;
  assign n3203 = x376 & n4050 ;
  assign n1050 = n3201 | n3203 ;
  assign n1051 = n1049 | n1050 ;
  assign n4051 = ~x377 ;
  assign n3205 = n4051 & x505 ;
  assign n4052 = ~x378 ;
  assign n3207 = n4052 & x506 ;
  assign n1052 = n3205 | n3207 ;
  assign n4053 = ~n1052 ;
  assign n1054 = n1051 & n4053 ;
  assign n1055 = n1053 | n1054 ;
  assign n4054 = ~n3307 ;
  assign n1056 = n4054 & n1055 ;
  assign n4055 = ~x508 ;
  assign n3209 = x380 & n4055 ;
  assign n4056 = ~x507 ;
  assign n3211 = x379 & n4056 ;
  assign n1057 = n3209 | n3211 ;
  assign n1058 = n1056 | n1057 ;
  assign n4057 = ~x381 ;
  assign n3213 = n4057 & x509 ;
  assign n4058 = ~x380 ;
  assign n3215 = n4058 & x508 ;
  assign n1059 = n3213 | n3215 ;
  assign n4059 = ~n1059 ;
  assign n1061 = n1058 & n4059 ;
  assign n1062 = n1060 | n1061 ;
  assign n4060 = ~x382 ;
  assign n3221 = n4060 & x510 ;
  assign n4061 = ~x511 ;
  assign n3223 = x383 & n4061 ;
  assign n1063 = n3221 | n3223 ;
  assign n4062 = ~n1063 ;
  assign n1064 = n1062 & n4062 ;
  assign n1065 = n3305 | n1064 ;
  assign n4063 = ~n1065 ;
  assign n1130 = x510 & n4063 ;
  assign n2817 = x382 & n1065 ;
  assign n2818 = n1130 | n2817 ;
  assign n1662 = x126 & n1606 ;
  assign n2819 = x254 & n3722 ;
  assign n2820 = n1662 | n2819 ;
  assign n4064 = ~n2820 ;
  assign n2826 = n2818 & n4064 ;
  assign n4065 = ~n3131 ;
  assign n2827 = n3129 & n4065 ;
  assign n2828 = n2826 | n2827 ;
  assign n4066 = ~n2818 ;
  assign n2821 = n4066 & n2820 ;
  assign n1746 = x381 & n1065 ;
  assign n2811 = x509 & n4063 ;
  assign n2812 = n1746 | n2811 ;
  assign n1812 = x253 & n3722 ;
  assign n2813 = x125 & n1606 ;
  assign n2814 = n1812 | n2813 ;
  assign n4067 = ~n2812 ;
  assign n2822 = n4067 & n2814 ;
  assign n2823 = n2821 | n2822 ;
  assign n1673 = x124 & n1606 ;
  assign n2802 = x252 & n3722 ;
  assign n2803 = n1673 | n2802 ;
  assign n1129 = x508 & n4063 ;
  assign n2804 = x380 & n1065 ;
  assign n2805 = n1129 | n2804 ;
  assign n4068 = ~n2803 ;
  assign n2810 = n4068 & n2805 ;
  assign n4069 = ~n2814 ;
  assign n2815 = n2812 & n4069 ;
  assign n2816 = n2810 | n2815 ;
  assign n4070 = ~n2805 ;
  assign n2806 = n2803 & n4070 ;
  assign n1745 = x379 & n1065 ;
  assign n2795 = x507 & n4063 ;
  assign n2796 = n1745 | n2795 ;
  assign n1786 = x251 & n3722 ;
  assign n2797 = x123 & n1606 ;
  assign n2798 = n1786 | n2797 ;
  assign n4071 = ~n2796 ;
  assign n2807 = n4071 & n2798 ;
  assign n2808 = n2806 | n2807 ;
  assign n1672 = x122 & n1606 ;
  assign n2786 = x250 & n3722 ;
  assign n2787 = n1672 | n2786 ;
  assign n1128 = x506 & n4063 ;
  assign n2788 = x378 & n1065 ;
  assign n2789 = n1128 | n2788 ;
  assign n4072 = ~n2787 ;
  assign n2794 = n4072 & n2789 ;
  assign n4073 = ~n2798 ;
  assign n2799 = n2796 & n4073 ;
  assign n2800 = n2794 | n2799 ;
  assign n1127 = x505 & n4063 ;
  assign n2778 = x377 & n1065 ;
  assign n2779 = n1127 | n2778 ;
  assign n1671 = x121 & n1606 ;
  assign n2780 = x249 & n3722 ;
  assign n2781 = n1671 | n2780 ;
  assign n4074 = ~n2779 ;
  assign n2785 = n4074 & n2781 ;
  assign n4075 = ~n2789 ;
  assign n2790 = n2787 & n4075 ;
  assign n2791 = n2785 | n2790 ;
  assign n4076 = ~n2781 ;
  assign n2782 = n2779 & n4076 ;
  assign n1811 = x248 & n3722 ;
  assign n2770 = x120 & n1606 ;
  assign n2771 = n1811 | n2770 ;
  assign n1687 = x376 & n1065 ;
  assign n2772 = x504 & n4063 ;
  assign n2773 = n1687 | n2772 ;
  assign n4077 = ~n2771 ;
  assign n2783 = n4077 & n2773 ;
  assign n2784 = n2782 | n2783 ;
  assign n4078 = ~n2773 ;
  assign n2774 = n2771 & n4078 ;
  assign n1099 = x503 & n4063 ;
  assign n2762 = x375 & n1065 ;
  assign n2763 = n1099 | n2762 ;
  assign n1637 = x119 & n1606 ;
  assign n2764 = x247 & n3722 ;
  assign n2765 = n1637 | n2764 ;
  assign n4079 = ~n2763 ;
  assign n2775 = n4079 & n2765 ;
  assign n2776 = n2774 | n2775 ;
  assign n4080 = ~n2765 ;
  assign n2766 = n2763 & n4080 ;
  assign n1711 = x374 & n1065 ;
  assign n2753 = x502 & n4063 ;
  assign n2754 = n1711 | n2753 ;
  assign n1750 = x246 & n3722 ;
  assign n2755 = x118 & n1606 ;
  assign n2756 = n1750 | n2755 ;
  assign n4081 = ~n2756 ;
  assign n2767 = n2754 & n4081 ;
  assign n2768 = n2766 | n2767 ;
  assign n1693 = x373 & n1065 ;
  assign n2747 = x501 & n4063 ;
  assign n2748 = n1693 | n2747 ;
  assign n1770 = x245 & n3722 ;
  assign n2749 = x117 & n1606 ;
  assign n2750 = n1770 | n2749 ;
  assign n4082 = ~n2748 ;
  assign n2757 = n4082 & n2750 ;
  assign n4083 = ~n2754 ;
  assign n2758 = n4083 & n2756 ;
  assign n2759 = n2757 | n2758 ;
  assign n1088 = x500 & n4063 ;
  assign n1132 = x372 & n1065 ;
  assign n1133 = n1088 | n1132 ;
  assign n1666 = x116 & n1606 ;
  assign n1677 = x244 & n3722 ;
  assign n1678 = n1666 | n1677 ;
  assign n4084 = ~n1678 ;
  assign n1679 = n1133 & n4084 ;
  assign n4085 = ~n2750 ;
  assign n2751 = n2748 & n4085 ;
  assign n2752 = n1679 | n2751 ;
  assign n4086 = ~n1133 ;
  assign n1680 = n4086 & n1678 ;
  assign n1729 = x371 & n1065 ;
  assign n1748 = x499 & n4063 ;
  assign n1749 = n1729 | n1748 ;
  assign n1798 = x243 & n3722 ;
  assign n1813 = x115 & n1606 ;
  assign n1814 = n1798 | n1813 ;
  assign n4087 = ~n1814 ;
  assign n1815 = n1749 & n4087 ;
  assign n4088 = ~n1749 ;
  assign n2740 = n4088 & n1814 ;
  assign n1670 = x114 & n1606 ;
  assign n2734 = x242 & n3722 ;
  assign n2735 = n1670 | n2734 ;
  assign n1113 = x498 & n4063 ;
  assign n2736 = x370 & n1065 ;
  assign n2737 = n1113 | n2736 ;
  assign n4089 = ~n2737 ;
  assign n2741 = n2735 & n4089 ;
  assign n2742 = n2740 | n2741 ;
  assign n1669 = x113 & n1606 ;
  assign n2725 = x241 & n3722 ;
  assign n2726 = n1669 | n2725 ;
  assign n1066 = x497 & n4063 ;
  assign n2727 = x369 & n1065 ;
  assign n2728 = n1066 | n2727 ;
  assign n4090 = ~n2726 ;
  assign n2733 = n4090 & n2728 ;
  assign n4091 = ~n2735 ;
  assign n2738 = n4091 & n2737 ;
  assign n2739 = n2733 | n2738 ;
  assign n4092 = ~n2728 ;
  assign n2729 = n2726 & n4092 ;
  assign n1744 = x368 & n1065 ;
  assign n2718 = x496 & n4063 ;
  assign n2719 = n1744 | n2718 ;
  assign n1772 = x240 & n3722 ;
  assign n2720 = x112 & n1606 ;
  assign n2721 = n1772 | n2720 ;
  assign n4093 = ~n2719 ;
  assign n2730 = n4093 & n2721 ;
  assign n2731 = n2729 | n2730 ;
  assign n1090 = x495 & n4063 ;
  assign n2708 = x367 & n1065 ;
  assign n2709 = n1090 | n2708 ;
  assign n1668 = x111 & n1606 ;
  assign n2710 = x239 & n3722 ;
  assign n2711 = n1668 | n2710 ;
  assign n4094 = ~n2711 ;
  assign n2717 = n2709 & n4094 ;
  assign n4095 = ~n2721 ;
  assign n2722 = n2719 & n4095 ;
  assign n2723 = n2717 | n2722 ;
  assign n4096 = ~n2709 ;
  assign n2712 = n4096 & n2711 ;
  assign n1067 = x494 & n4063 ;
  assign n2701 = x366 & n1065 ;
  assign n2702 = n1067 | n2701 ;
  assign n1623 = x110 & n1606 ;
  assign n2703 = x238 & n3722 ;
  assign n2704 = n1623 | n2703 ;
  assign n4097 = ~n2702 ;
  assign n2713 = n4097 & n2704 ;
  assign n2714 = n2712 | n2713 ;
  assign n4098 = ~n2704 ;
  assign n2705 = n2702 & n4098 ;
  assign n1736 = x365 & n1065 ;
  assign n2694 = x493 & n4063 ;
  assign n2695 = n1736 | n2694 ;
  assign n1781 = x237 & n3722 ;
  assign n2696 = x109 & n1606 ;
  assign n2697 = n1781 | n2696 ;
  assign n4099 = ~n2697 ;
  assign n2706 = n2695 & n4099 ;
  assign n2707 = n2705 | n2706 ;
  assign n1721 = x364 & n1065 ;
  assign n2685 = x492 & n4063 ;
  assign n2686 = n1721 | n2685 ;
  assign n1752 = x236 & n3722 ;
  assign n2687 = x108 & n1606 ;
  assign n2688 = n1752 | n2687 ;
  assign n4100 = ~n2686 ;
  assign n2693 = n4100 & n2688 ;
  assign n4101 = ~n2695 ;
  assign n2698 = n4101 & n2697 ;
  assign n2699 = n2693 | n2698 ;
  assign n4102 = ~n2688 ;
  assign n2689 = n2686 & n4102 ;
  assign n1077 = x491 & n4063 ;
  assign n2676 = x363 & n1065 ;
  assign n2677 = n1077 | n2676 ;
  assign n1607 = x107 & n1606 ;
  assign n2678 = x235 & n3722 ;
  assign n2679 = n1607 | n2678 ;
  assign n4103 = ~n2679 ;
  assign n2690 = n2677 & n4103 ;
  assign n2691 = n2689 | n2690 ;
  assign n4104 = ~n2677 ;
  assign n2680 = n4104 & n2679 ;
  assign n1704 = x362 & n1065 ;
  assign n2669 = x490 & n4063 ;
  assign n2670 = n1704 | n2669 ;
  assign n1753 = x234 & n3722 ;
  assign n2671 = x106 & n1606 ;
  assign n2672 = n1753 | n2671 ;
  assign n4105 = ~n2670 ;
  assign n2681 = n4105 & n2672 ;
  assign n2682 = n2680 | n2681 ;
  assign n4106 = ~n2672 ;
  assign n2673 = n2670 & n4106 ;
  assign n1791 = x233 & n3722 ;
  assign n2661 = x105 & n1606 ;
  assign n2662 = n1791 | n2661 ;
  assign n1702 = x361 & n1065 ;
  assign n2663 = x489 & n4063 ;
  assign n2664 = n1702 | n2663 ;
  assign n4107 = ~n2662 ;
  assign n2674 = n4107 & n2664 ;
  assign n2675 = n2673 | n2674 ;
  assign n4108 = ~n2664 ;
  assign n2665 = n2662 & n4108 ;
  assign n1078 = x488 & n4063 ;
  assign n2654 = x360 & n1065 ;
  assign n2655 = n1078 | n2654 ;
  assign n1652 = x104 & n1606 ;
  assign n2656 = x232 & n3722 ;
  assign n2657 = n1652 | n2656 ;
  assign n4109 = ~n2655 ;
  assign n2666 = n4109 & n2657 ;
  assign n2667 = n2665 | n2666 ;
  assign n1755 = x231 & n3722 ;
  assign n2644 = x103 & n1606 ;
  assign n2645 = n1755 | n2644 ;
  assign n1681 = x359 & n1065 ;
  assign n2646 = x487 & n4063 ;
  assign n2647 = n1681 | n2646 ;
  assign n4110 = ~n2645 ;
  assign n2653 = n4110 & n2647 ;
  assign n4111 = ~n2657 ;
  assign n2658 = n2655 & n4111 ;
  assign n2659 = n2653 | n2658 ;
  assign n4112 = ~n2647 ;
  assign n2648 = n2645 & n4112 ;
  assign n1085 = x486 & n4063 ;
  assign n2638 = x358 & n1065 ;
  assign n2639 = n1085 | n2638 ;
  assign n1609 = x102 & n1606 ;
  assign n2640 = x230 & n3722 ;
  assign n2641 = n1609 | n2640 ;
  assign n4113 = ~n2639 ;
  assign n2649 = n4113 & n2641 ;
  assign n2650 = n2648 | n2649 ;
  assign n1714 = x357 & n1065 ;
  assign n2629 = x485 & n4063 ;
  assign n2630 = n1714 | n2629 ;
  assign n1766 = x229 & n3722 ;
  assign n2631 = x101 & n1606 ;
  assign n2632 = n1766 | n2631 ;
  assign n4114 = ~n2632 ;
  assign n2637 = n2630 & n4114 ;
  assign n4115 = ~n2641 ;
  assign n2642 = n2639 & n4115 ;
  assign n2643 = n2637 | n2642 ;
  assign n4116 = ~n2630 ;
  assign n2633 = n4116 & n2632 ;
  assign n1757 = x228 & n3722 ;
  assign n2621 = x100 & n1606 ;
  assign n2622 = n1757 | n2621 ;
  assign n1724 = x356 & n1065 ;
  assign n2623 = x484 & n4063 ;
  assign n2624 = n1724 | n2623 ;
  assign n4117 = ~n2624 ;
  assign n2634 = n2622 & n4117 ;
  assign n2635 = n2633 | n2634 ;
  assign n4118 = ~n2622 ;
  assign n2625 = n4118 & n2624 ;
  assign n1068 = x483 & n4063 ;
  assign n2612 = x355 & n1065 ;
  assign n2613 = n1068 | n2612 ;
  assign n1610 = x99 & n1606 ;
  assign n2614 = x227 & n3722 ;
  assign n2615 = n1610 | n2614 ;
  assign n4119 = ~n2615 ;
  assign n2626 = n2613 & n4119 ;
  assign n2627 = n2625 | n2626 ;
  assign n4120 = ~n2613 ;
  assign n2616 = n4120 & n2615 ;
  assign n1682 = x354 & n1065 ;
  assign n2605 = x482 & n4063 ;
  assign n2606 = n1682 | n2605 ;
  assign n1758 = x226 & n3722 ;
  assign n2607 = x98 & n1606 ;
  assign n2608 = n1758 | n2607 ;
  assign n4121 = ~n2606 ;
  assign n2617 = n4121 & n2608 ;
  assign n2618 = n2616 | n2617 ;
  assign n4122 = ~n2608 ;
  assign n2609 = n2606 & n4122 ;
  assign n1685 = x353 & n1065 ;
  assign n2597 = x481 & n4063 ;
  assign n2598 = n1685 | n2597 ;
  assign n1759 = x225 & n3722 ;
  assign n2599 = x97 & n1606 ;
  assign n2600 = n1759 | n2599 ;
  assign n4123 = ~n2600 ;
  assign n2610 = n2598 & n4123 ;
  assign n2611 = n2609 | n2610 ;
  assign n4124 = ~n2598 ;
  assign n2601 = n4124 & n2600 ;
  assign n1611 = x96 & n1606 ;
  assign n2590 = x224 & n3722 ;
  assign n2591 = n1611 | n2590 ;
  assign n1070 = x480 & n4063 ;
  assign n2592 = x352 & n1065 ;
  assign n2593 = n1070 | n2592 ;
  assign n4125 = ~n2593 ;
  assign n2602 = n2591 & n4125 ;
  assign n2603 = n2601 | n2602 ;
  assign n1613 = x95 & n1606 ;
  assign n2581 = x223 & n3722 ;
  assign n2582 = n1613 | n2581 ;
  assign n1072 = x479 & n4063 ;
  assign n2583 = x351 & n1065 ;
  assign n2584 = n1072 | n2583 ;
  assign n4126 = ~n2582 ;
  assign n2589 = n4126 & n2584 ;
  assign n4127 = ~n2591 ;
  assign n2594 = n4127 & n2593 ;
  assign n2595 = n2589 | n2594 ;
  assign n1797 = x222 & n3722 ;
  assign n2574 = x94 & n1606 ;
  assign n2575 = n1797 | n2574 ;
  assign n1686 = x350 & n1065 ;
  assign n2576 = x478 & n4063 ;
  assign n2577 = n1686 | n2576 ;
  assign n4128 = ~n2577 ;
  assign n2580 = n2575 & n4128 ;
  assign n4129 = ~n2584 ;
  assign n2585 = n2582 & n4129 ;
  assign n2586 = n2580 | n2585 ;
  assign n1073 = x477 & n4063 ;
  assign n2565 = x349 & n1065 ;
  assign n2566 = n1073 | n2565 ;
  assign n1648 = x93 & n1606 ;
  assign n2567 = x221 & n3722 ;
  assign n2568 = n1648 | n2567 ;
  assign n4130 = ~n2568 ;
  assign n2573 = n2566 & n4130 ;
  assign n4131 = ~n2575 ;
  assign n2578 = n4131 & n2577 ;
  assign n2579 = n2573 | n2578 ;
  assign n4132 = ~n2566 ;
  assign n2569 = n4132 & n2568 ;
  assign n1761 = x220 & n3722 ;
  assign n2557 = x92 & n1606 ;
  assign n2558 = n1761 | n2557 ;
  assign n1688 = x348 & n1065 ;
  assign n2559 = x476 & n4063 ;
  assign n2560 = n1688 | n2559 ;
  assign n4133 = ~n2560 ;
  assign n2570 = n2558 & n4133 ;
  assign n2571 = n2569 | n2570 ;
  assign n4134 = ~n2558 ;
  assign n2561 = n4134 & n2560 ;
  assign n1081 = x475 & n4063 ;
  assign n2548 = x347 & n1065 ;
  assign n2549 = n1081 | n2548 ;
  assign n1620 = x91 & n1606 ;
  assign n2550 = x219 & n3722 ;
  assign n2551 = n1620 | n2550 ;
  assign n4135 = ~n2551 ;
  assign n2562 = n2549 & n4135 ;
  assign n2563 = n2561 | n2562 ;
  assign n4136 = ~n2549 ;
  assign n2552 = n4136 & n2551 ;
  assign n1074 = x474 & n4063 ;
  assign n2542 = x346 & n1065 ;
  assign n2543 = n1074 | n2542 ;
  assign n1762 = x218 & n3722 ;
  assign n2544 = x90 & n1606 ;
  assign n2545 = n1762 | n2544 ;
  assign n4137 = ~n2543 ;
  assign n2553 = n4137 & n2545 ;
  assign n2554 = n2552 | n2553 ;
  assign n1763 = x217 & n3722 ;
  assign n2533 = x89 & n1606 ;
  assign n2534 = n1763 | n2533 ;
  assign n1733 = x345 & n1065 ;
  assign n2535 = x473 & n4063 ;
  assign n2536 = n1733 | n2535 ;
  assign n4138 = ~n2534 ;
  assign n2541 = n4138 & n2536 ;
  assign n4139 = ~n2545 ;
  assign n2546 = n2543 & n4139 ;
  assign n2547 = n2541 | n2546 ;
  assign n4140 = ~n2536 ;
  assign n2537 = n2534 & n4140 ;
  assign n1095 = x472 & n4063 ;
  assign n2526 = x344 & n1065 ;
  assign n2527 = n1095 | n2526 ;
  assign n1614 = x88 & n1606 ;
  assign n2528 = x216 & n3722 ;
  assign n2529 = n1614 | n2528 ;
  assign n4141 = ~n2527 ;
  assign n2538 = n4141 & n2529 ;
  assign n2539 = n2537 | n2538 ;
  assign n1765 = x215 & n3722 ;
  assign n2516 = x87 & n1606 ;
  assign n2517 = n1765 | n2516 ;
  assign n1689 = x343 & n1065 ;
  assign n2518 = x471 & n4063 ;
  assign n2519 = n1689 | n2518 ;
  assign n4142 = ~n2517 ;
  assign n2525 = n4142 & n2519 ;
  assign n4143 = ~n2529 ;
  assign n2530 = n2527 & n4143 ;
  assign n2531 = n2525 | n2530 ;
  assign n4144 = ~n2519 ;
  assign n2520 = n2517 & n4144 ;
  assign n1723 = x342 & n1065 ;
  assign n1816 = x470 & n4063 ;
  assign n1817 = n1723 | n1816 ;
  assign n1659 = x86 & n1606 ;
  assign n1818 = x214 & n3722 ;
  assign n1819 = n1659 | n1818 ;
  assign n4145 = ~n1817 ;
  assign n2521 = n4145 & n1819 ;
  assign n2522 = n2520 | n2521 ;
  assign n4146 = ~n1819 ;
  assign n1820 = n1817 & n4146 ;
  assign n1116 = x469 & n4063 ;
  assign n1821 = x341 & n1065 ;
  assign n1822 = n1116 | n1821 ;
  assign n1658 = x85 & n1606 ;
  assign n1823 = x213 & n3722 ;
  assign n1824 = n1658 | n1823 ;
  assign n4147 = ~n1822 ;
  assign n1825 = n4147 & n1824 ;
  assign n4148 = ~n1824 ;
  assign n2511 = n1822 & n4148 ;
  assign n1760 = x212 & n3722 ;
  assign n2503 = x84 & n1606 ;
  assign n2504 = n1760 | n2503 ;
  assign n1694 = x340 & n1065 ;
  assign n2505 = x468 & n4063 ;
  assign n2506 = n1694 | n2505 ;
  assign n4149 = ~n2504 ;
  assign n2512 = n4149 & n2506 ;
  assign n2513 = n2511 | n2512 ;
  assign n1612 = x83 & n1606 ;
  assign n1826 = x211 & n3722 ;
  assign n1827 = n1612 | n1826 ;
  assign n1106 = x467 & n4063 ;
  assign n1828 = x339 & n1065 ;
  assign n1829 = n1106 | n1828 ;
  assign n4150 = ~n1829 ;
  assign n2502 = n1827 & n4150 ;
  assign n4151 = ~n2506 ;
  assign n2507 = n2504 & n4151 ;
  assign n2508 = n2502 | n2507 ;
  assign n4152 = ~n1827 ;
  assign n1830 = n4152 & n1829 ;
  assign n1651 = x82 & n1606 ;
  assign n1831 = x210 & n3722 ;
  assign n1832 = n1651 | n1831 ;
  assign n1109 = x466 & n4063 ;
  assign n1833 = x338 & n1065 ;
  assign n1834 = n1109 | n1833 ;
  assign n4153 = ~n1834 ;
  assign n1835 = n1832 & n4153 ;
  assign n1789 = x209 & n3722 ;
  assign n2488 = x81 & n1606 ;
  assign n2489 = n1789 | n2488 ;
  assign n1076 = x465 & n4063 ;
  assign n2490 = x337 & n1065 ;
  assign n2491 = n1076 | n2490 ;
  assign n4154 = ~n2489 ;
  assign n2497 = n4154 & n2491 ;
  assign n4155 = ~n1832 ;
  assign n2498 = n4155 & n1834 ;
  assign n2499 = n2497 | n2498 ;
  assign n1616 = x80 & n1606 ;
  assign n2482 = x208 & n3722 ;
  assign n2483 = n1616 | n2482 ;
  assign n1071 = x464 & n4063 ;
  assign n2484 = x336 & n1065 ;
  assign n2485 = n1071 | n2484 ;
  assign n4156 = ~n2485 ;
  assign n2492 = n2483 & n4156 ;
  assign n4157 = ~n2491 ;
  assign n2493 = n2489 & n4157 ;
  assign n2494 = n2492 | n2493 ;
  assign n1101 = x463 & n4063 ;
  assign n1836 = x335 & n1065 ;
  assign n1837 = n1101 | n1836 ;
  assign n1639 = x79 & n1606 ;
  assign n1838 = x207 & n3722 ;
  assign n1839 = n1639 | n1838 ;
  assign n4158 = ~n1839 ;
  assign n1840 = n1837 & n4158 ;
  assign n4159 = ~n2483 ;
  assign n2486 = n4159 & n2485 ;
  assign n2487 = n1840 | n2486 ;
  assign n4160 = ~n1837 ;
  assign n1841 = n4160 & n1839 ;
  assign n1098 = x462 & n4063 ;
  assign n1842 = x334 & n1065 ;
  assign n1843 = n1098 | n1842 ;
  assign n1793 = x206 & n3722 ;
  assign n1844 = x78 & n1606 ;
  assign n1845 = n1793 | n1844 ;
  assign n4161 = ~n1845 ;
  assign n1846 = n1843 & n4161 ;
  assign n4162 = ~n1843 ;
  assign n2475 = n4162 & n1845 ;
  assign n1617 = x77 & n1606 ;
  assign n2469 = x205 & n3722 ;
  assign n2470 = n1617 | n2469 ;
  assign n1080 = x461 & n4063 ;
  assign n2471 = x333 & n1065 ;
  assign n2472 = n1080 | n2471 ;
  assign n4163 = ~n2472 ;
  assign n2476 = n2470 & n4163 ;
  assign n2477 = n2475 | n2476 ;
  assign n1618 = x76 & n1606 ;
  assign n2460 = x204 & n3722 ;
  assign n2461 = n1618 | n2460 ;
  assign n1107 = x460 & n4063 ;
  assign n2462 = x332 & n1065 ;
  assign n2463 = n1107 | n2462 ;
  assign n4164 = ~n2461 ;
  assign n2468 = n4164 & n2463 ;
  assign n4165 = ~n2470 ;
  assign n2473 = n4165 & n2472 ;
  assign n2474 = n2468 | n2473 ;
  assign n4166 = ~n2463 ;
  assign n2464 = n2461 & n4166 ;
  assign n1075 = x459 & n4063 ;
  assign n1847 = x331 & n1065 ;
  assign n1848 = n1075 | n1847 ;
  assign n1779 = x203 & n3722 ;
  assign n1849 = x75 & n1606 ;
  assign n1850 = n1779 | n1849 ;
  assign n4167 = ~n1848 ;
  assign n2465 = n4167 & n1850 ;
  assign n2466 = n2464 | n2465 ;
  assign n4168 = ~n1850 ;
  assign n1851 = n1848 & n4168 ;
  assign n1718 = x330 & n1065 ;
  assign n1852 = x458 & n4063 ;
  assign n1853 = n1718 | n1852 ;
  assign n1633 = x74 & n1606 ;
  assign n1854 = x202 & n3722 ;
  assign n1855 = n1633 | n1854 ;
  assign n4169 = ~n1853 ;
  assign n1856 = n4169 & n1855 ;
  assign n4170 = ~n1855 ;
  assign n2454 = n1853 & n4170 ;
  assign n1656 = x73 & n1606 ;
  assign n2447 = x201 & n3722 ;
  assign n2448 = n1656 | n2447 ;
  assign n1083 = x457 & n4063 ;
  assign n2449 = x329 & n1065 ;
  assign n2450 = n1083 | n2449 ;
  assign n4171 = ~n2448 ;
  assign n2455 = n4171 & n2450 ;
  assign n2456 = n2454 | n2455 ;
  assign n1806 = x200 & n3722 ;
  assign n2438 = x72 & n1606 ;
  assign n2439 = n1806 | n2438 ;
  assign n1737 = x328 & n1065 ;
  assign n2440 = x456 & n4063 ;
  assign n2441 = n1737 | n2440 ;
  assign n4172 = ~n2441 ;
  assign n2446 = n2439 & n4172 ;
  assign n4173 = ~n2450 ;
  assign n2451 = n2448 & n4173 ;
  assign n2452 = n2446 | n2451 ;
  assign n4174 = ~n2439 ;
  assign n2442 = n4174 & n2441 ;
  assign n1642 = x71 & n1606 ;
  assign n2429 = x199 & n3722 ;
  assign n2430 = n1642 | n2429 ;
  assign n1691 = x327 & n1065 ;
  assign n2431 = x455 & n4063 ;
  assign n2432 = n1691 | n2431 ;
  assign n4175 = ~n2430 ;
  assign n2443 = n4175 & n2432 ;
  assign n2444 = n2442 | n2443 ;
  assign n4176 = ~n2432 ;
  assign n2433 = n2430 & n4176 ;
  assign n1091 = x454 & n4063 ;
  assign n2422 = x326 & n1065 ;
  assign n2423 = n1091 | n2422 ;
  assign n1767 = x198 & n3722 ;
  assign n2424 = x70 & n1606 ;
  assign n2425 = n1767 | n2424 ;
  assign n4177 = ~n2423 ;
  assign n2434 = n4177 & n2425 ;
  assign n2435 = n2433 | n2434 ;
  assign n4178 = ~n2425 ;
  assign n2426 = n2423 & n4178 ;
  assign n1692 = x325 & n1065 ;
  assign n2414 = x453 & n4063 ;
  assign n2415 = n1692 | n2414 ;
  assign n1638 = x69 & n1606 ;
  assign n2416 = x197 & n3722 ;
  assign n2417 = n1638 | n2416 ;
  assign n4179 = ~n2417 ;
  assign n2427 = n2415 & n4179 ;
  assign n2428 = n2426 | n2427 ;
  assign n1619 = x68 & n1606 ;
  assign n2407 = x196 & n3722 ;
  assign n2408 = n1619 | n2407 ;
  assign n1695 = x324 & n1065 ;
  assign n2409 = x452 & n4063 ;
  assign n2410 = n1695 | n2409 ;
  assign n4180 = ~n2410 ;
  assign n2418 = n2408 & n4180 ;
  assign n4181 = ~n2415 ;
  assign n2419 = n4181 & n2417 ;
  assign n2420 = n2418 | n2419 ;
  assign n1751 = x195 & n3722 ;
  assign n1857 = x67 & n1606 ;
  assign n1858 = n1751 | n1857 ;
  assign n1097 = x451 & n4063 ;
  assign n1859 = x323 & n1065 ;
  assign n1860 = n1097 | n1859 ;
  assign n4182 = ~n1858 ;
  assign n1861 = n4182 & n1860 ;
  assign n4183 = ~n2408 ;
  assign n2411 = n4183 & n2410 ;
  assign n2412 = n1861 | n2411 ;
  assign n4184 = ~n1860 ;
  assign n2404 = n1858 & n4184 ;
  assign n1635 = x66 & n1606 ;
  assign n1862 = x194 & n3722 ;
  assign n1863 = n1635 | n1862 ;
  assign n1712 = x322 & n1065 ;
  assign n1864 = x450 & n4063 ;
  assign n1865 = n1712 | n1864 ;
  assign n4185 = ~n1863 ;
  assign n1866 = n4185 & n1865 ;
  assign n1754 = x193 & n3722 ;
  assign n2393 = x65 & n1606 ;
  assign n2394 = n1754 | n2393 ;
  assign n1717 = x321 & n1065 ;
  assign n2395 = x449 & n4063 ;
  assign n2396 = n1717 | n2395 ;
  assign n4186 = ~n2396 ;
  assign n2400 = n2394 & n4186 ;
  assign n4187 = ~n1865 ;
  assign n2401 = n1863 & n4187 ;
  assign n2402 = n2400 | n2401 ;
  assign n1636 = x64 & n1606 ;
  assign n1867 = x192 & n3722 ;
  assign n1868 = n1636 | n1867 ;
  assign n1102 = x448 & n4063 ;
  assign n1869 = x320 & n1065 ;
  assign n1870 = n1102 | n1869 ;
  assign n4188 = ~n1868 ;
  assign n1871 = n4188 & n1870 ;
  assign n4189 = ~n2394 ;
  assign n2397 = n4189 & n2396 ;
  assign n2398 = n1871 | n2397 ;
  assign n4190 = ~n1870 ;
  assign n2390 = n1868 & n4190 ;
  assign n1768 = x191 & n3722 ;
  assign n1872 = x63 & n1606 ;
  assign n1873 = n1768 | n1872 ;
  assign n1716 = x319 & n1065 ;
  assign n1874 = x447 & n4063 ;
  assign n1875 = n1716 | n1874 ;
  assign n4191 = ~n1873 ;
  assign n1876 = n4191 & n1875 ;
  assign n1621 = x62 & n1606 ;
  assign n2379 = x190 & n3722 ;
  assign n2380 = n1621 | n2379 ;
  assign n1079 = x446 & n4063 ;
  assign n2381 = x318 & n1065 ;
  assign n2382 = n1079 | n2381 ;
  assign n4192 = ~n2382 ;
  assign n2386 = n2380 & n4192 ;
  assign n4193 = ~n1875 ;
  assign n2387 = n1873 & n4193 ;
  assign n2388 = n2386 | n2387 ;
  assign n1608 = x61 & n1606 ;
  assign n2369 = x189 & n3722 ;
  assign n2370 = n1608 | n2369 ;
  assign n1084 = x445 & n4063 ;
  assign n2371 = x317 & n1065 ;
  assign n2372 = n1084 | n2371 ;
  assign n4194 = ~n2370 ;
  assign n2378 = n4194 & n2372 ;
  assign n4195 = ~n2380 ;
  assign n2383 = n4195 & n2382 ;
  assign n2384 = n2378 | n2383 ;
  assign n4196 = ~n2372 ;
  assign n2373 = n2370 & n4196 ;
  assign n1715 = x316 & n1065 ;
  assign n1877 = x444 & n4063 ;
  assign n1878 = n1715 | n1877 ;
  assign n1645 = x60 & n1606 ;
  assign n1879 = x188 & n3722 ;
  assign n1880 = n1645 | n1879 ;
  assign n4197 = ~n1878 ;
  assign n2374 = n4197 & n1880 ;
  assign n2375 = n2373 | n2374 ;
  assign n4198 = ~n1880 ;
  assign n1881 = n1878 & n4198 ;
  assign n1120 = x443 & n4063 ;
  assign n1882 = x315 & n1065 ;
  assign n1883 = n1120 | n1882 ;
  assign n1787 = x187 & n3722 ;
  assign n1884 = x59 & n1606 ;
  assign n1885 = n1787 | n1884 ;
  assign n4199 = ~n1883 ;
  assign n1886 = n4199 & n1885 ;
  assign n4200 = ~n1885 ;
  assign n2364 = n1883 & n4200 ;
  assign n1622 = x58 & n1606 ;
  assign n2356 = x186 & n3722 ;
  assign n2357 = n1622 | n2356 ;
  assign n1697 = x314 & n1065 ;
  assign n2358 = x442 & n4063 ;
  assign n2359 = n1697 | n2358 ;
  assign n4201 = ~n2357 ;
  assign n2365 = n4201 & n2359 ;
  assign n2366 = n2364 | n2365 ;
  assign n1782 = x185 & n3722 ;
  assign n2349 = x57 & n1606 ;
  assign n2350 = n1782 | n2349 ;
  assign n1698 = x313 & n1065 ;
  assign n2351 = x441 & n4063 ;
  assign n2352 = n1698 | n2351 ;
  assign n4202 = ~n2352 ;
  assign n2355 = n2350 & n4202 ;
  assign n4203 = ~n2359 ;
  assign n2360 = n2357 & n4203 ;
  assign n2361 = n2355 | n2360 ;
  assign n1114 = x440 & n4063 ;
  assign n2340 = x312 & n1065 ;
  assign n2341 = n1114 | n2340 ;
  assign n1769 = x184 & n3722 ;
  assign n2342 = x56 & n1606 ;
  assign n2343 = n1769 | n2342 ;
  assign n4204 = ~n2343 ;
  assign n2348 = n2341 & n4204 ;
  assign n4205 = ~n2350 ;
  assign n2353 = n4205 & n2352 ;
  assign n2354 = n2348 | n2353 ;
  assign n4206 = ~n2341 ;
  assign n2344 = n4206 & n2343 ;
  assign n1624 = x55 & n1606 ;
  assign n2333 = x183 & n3722 ;
  assign n2334 = n1624 | n2333 ;
  assign n1696 = x311 & n1065 ;
  assign n2335 = x439 & n4063 ;
  assign n2336 = n1696 | n2335 ;
  assign n4207 = ~n2336 ;
  assign n2345 = n2334 & n4207 ;
  assign n2346 = n2344 | n2345 ;
  assign n1731 = x310 & n1065 ;
  assign n2323 = x438 & n4063 ;
  assign n2324 = n1731 | n2323 ;
  assign n1632 = x54 & n1606 ;
  assign n2325 = x182 & n3722 ;
  assign n2326 = n1632 | n2325 ;
  assign n4208 = ~n2326 ;
  assign n2332 = n2324 & n4208 ;
  assign n4209 = ~n2334 ;
  assign n2337 = n4209 & n2336 ;
  assign n2338 = n2332 | n2337 ;
  assign n4210 = ~n2324 ;
  assign n2327 = n4210 & n2326 ;
  assign n1086 = x437 & n4063 ;
  assign n2316 = x309 & n1065 ;
  assign n2317 = n1086 | n2316 ;
  assign n1771 = x181 & n3722 ;
  assign n2318 = x53 & n1606 ;
  assign n2319 = n1771 | n2318 ;
  assign n4211 = ~n2317 ;
  assign n2328 = n4211 & n2319 ;
  assign n2329 = n2327 | n2328 ;
  assign n4212 = ~n2319 ;
  assign n2320 = n2317 & n4212 ;
  assign n1699 = x308 & n1065 ;
  assign n2309 = x436 & n4063 ;
  assign n2310 = n1699 | n2309 ;
  assign n1625 = x52 & n1606 ;
  assign n2311 = x180 & n3722 ;
  assign n2312 = n1625 | n2311 ;
  assign n4213 = ~n2312 ;
  assign n2321 = n2310 & n4213 ;
  assign n2322 = n2320 | n2321 ;
  assign n1626 = x51 & n1606 ;
  assign n2300 = x179 & n3722 ;
  assign n2301 = n1626 | n2300 ;
  assign n1740 = x307 & n1065 ;
  assign n2302 = x435 & n4063 ;
  assign n2303 = n1740 | n2302 ;
  assign n4214 = ~n2303 ;
  assign n2308 = n2301 & n4214 ;
  assign n4215 = ~n2310 ;
  assign n2313 = n4215 & n2312 ;
  assign n2314 = n2308 | n2313 ;
  assign n4216 = ~n2301 ;
  assign n2304 = n4216 & n2303 ;
  assign n1069 = x434 & n4063 ;
  assign n2292 = x306 & n1065 ;
  assign n2293 = n1069 | n2292 ;
  assign n1776 = x178 & n3722 ;
  assign n2294 = x50 & n1606 ;
  assign n2295 = n1776 | n2294 ;
  assign n4217 = ~n2295 ;
  assign n2305 = n2293 & n4217 ;
  assign n2306 = n2304 | n2305 ;
  assign n1773 = x177 & n3722 ;
  assign n2284 = x49 & n1606 ;
  assign n2285 = n1773 | n2284 ;
  assign n1727 = x305 & n1065 ;
  assign n2286 = x433 & n4063 ;
  assign n2287 = n1727 | n2286 ;
  assign n4218 = ~n2287 ;
  assign n2291 = n2285 & n4218 ;
  assign n4219 = ~n2293 ;
  assign n2296 = n4219 & n2295 ;
  assign n2297 = n2291 | n2296 ;
  assign n4220 = ~n2285 ;
  assign n2288 = n4220 & n2287 ;
  assign n1087 = x432 & n4063 ;
  assign n2276 = x304 & n1065 ;
  assign n2277 = n1087 | n2276 ;
  assign n1650 = x48 & n1606 ;
  assign n2278 = x176 & n3722 ;
  assign n2279 = n1650 | n2278 ;
  assign n4221 = ~n2279 ;
  assign n2289 = n2277 & n4221 ;
  assign n2290 = n2288 | n2289 ;
  assign n1701 = x303 & n1065 ;
  assign n2269 = x431 & n4063 ;
  assign n2270 = n1701 | n2269 ;
  assign n1660 = x47 & n1606 ;
  assign n2271 = x175 & n3722 ;
  assign n2272 = n1660 | n2271 ;
  assign n4222 = ~n2270 ;
  assign n2280 = n4222 & n2272 ;
  assign n4223 = ~n2277 ;
  assign n2281 = n4223 & n2279 ;
  assign n2282 = n2280 | n2281 ;
  assign n1094 = x430 & n4063 ;
  assign n1887 = x302 & n1065 ;
  assign n1888 = n1094 | n1887 ;
  assign n1785 = x174 & n3722 ;
  assign n1889 = x46 & n1606 ;
  assign n1890 = n1785 | n1889 ;
  assign n4224 = ~n1890 ;
  assign n1891 = n1888 & n4224 ;
  assign n4225 = ~n2272 ;
  assign n2273 = n2270 & n4225 ;
  assign n2274 = n1891 | n2273 ;
  assign n4226 = ~n1888 ;
  assign n2266 = n4226 & n1890 ;
  assign n1700 = x301 & n1065 ;
  assign n1892 = x429 & n4063 ;
  assign n1893 = n1700 | n1892 ;
  assign n1792 = x173 & n3722 ;
  assign n1894 = x45 & n1606 ;
  assign n1895 = n1792 | n1894 ;
  assign n4227 = ~n1895 ;
  assign n1896 = n1893 & n4227 ;
  assign n1630 = x44 & n1606 ;
  assign n2254 = x172 & n3722 ;
  assign n2255 = n1630 | n2254 ;
  assign n1703 = x300 & n1065 ;
  assign n2256 = x428 & n4063 ;
  assign n2257 = n1703 | n2256 ;
  assign n4228 = ~n2257 ;
  assign n2262 = n2255 & n4228 ;
  assign n4229 = ~n1893 ;
  assign n2263 = n4229 & n1895 ;
  assign n2264 = n2262 | n2263 ;
  assign n4230 = ~n2255 ;
  assign n2258 = n4230 & n2257 ;
  assign n1104 = x427 & n4063 ;
  assign n2246 = x299 & n1065 ;
  assign n2247 = n1104 | n2246 ;
  assign n1800 = x171 & n3722 ;
  assign n2248 = x43 & n1606 ;
  assign n2249 = n1800 | n2248 ;
  assign n4231 = ~n2249 ;
  assign n2259 = n2247 & n4231 ;
  assign n2260 = n2258 | n2259 ;
  assign n1705 = x298 & n1065 ;
  assign n2239 = x426 & n4063 ;
  assign n2240 = n1705 | n2239 ;
  assign n1774 = x170 & n3722 ;
  assign n2241 = x42 & n1606 ;
  assign n2242 = n1774 | n2241 ;
  assign n4232 = ~n2240 ;
  assign n2245 = n4232 & n2242 ;
  assign n4233 = ~n2247 ;
  assign n2250 = n4233 & n2249 ;
  assign n2251 = n2245 | n2250 ;
  assign n1105 = x425 & n4063 ;
  assign n2230 = x297 & n1065 ;
  assign n2231 = n1105 | n2230 ;
  assign n1627 = x41 & n1606 ;
  assign n2232 = x169 & n3722 ;
  assign n2233 = n1627 | n2232 ;
  assign n4234 = ~n2233 ;
  assign n2238 = n2231 & n4234 ;
  assign n4235 = ~n2242 ;
  assign n2243 = n2240 & n4235 ;
  assign n2244 = n2238 | n2243 ;
  assign n4236 = ~n2231 ;
  assign n2234 = n4236 & n2233 ;
  assign n1710 = x296 & n1065 ;
  assign n1897 = x424 & n4063 ;
  assign n1898 = n1710 | n1897 ;
  assign n1644 = x40 & n1606 ;
  assign n1899 = x168 & n3722 ;
  assign n1900 = n1644 | n1899 ;
  assign n4237 = ~n1898 ;
  assign n2235 = n4237 & n1900 ;
  assign n2236 = n2234 | n2235 ;
  assign n4238 = ~n1900 ;
  assign n1901 = n1898 & n4238 ;
  assign n1103 = x423 & n4063 ;
  assign n1902 = x295 & n1065 ;
  assign n1903 = n1103 | n1902 ;
  assign n1780 = x167 & n3722 ;
  assign n1904 = x39 & n1606 ;
  assign n1905 = n1780 | n1904 ;
  assign n4239 = ~n1903 ;
  assign n1906 = n4239 & n1905 ;
  assign n1628 = x38 & n1606 ;
  assign n2216 = x166 & n3722 ;
  assign n2217 = n1628 | n2216 ;
  assign n1706 = x294 & n1065 ;
  assign n2218 = x422 & n4063 ;
  assign n2219 = n1706 | n2218 ;
  assign n4240 = ~n2217 ;
  assign n2224 = n4240 & n2219 ;
  assign n4241 = ~n1905 ;
  assign n2225 = n1903 & n4241 ;
  assign n2226 = n2224 | n2225 ;
  assign n1743 = x293 & n1065 ;
  assign n2209 = x421 & n4063 ;
  assign n2210 = n1743 | n2209 ;
  assign n1775 = x165 & n3722 ;
  assign n2211 = x37 & n1606 ;
  assign n2212 = n1775 | n2211 ;
  assign n4242 = ~n2210 ;
  assign n2220 = n4242 & n2212 ;
  assign n4243 = ~n2219 ;
  assign n2221 = n2217 & n4243 ;
  assign n2222 = n2220 | n2221 ;
  assign n1640 = x36 & n1606 ;
  assign n1907 = x164 & n3722 ;
  assign n1908 = n1640 | n1907 ;
  assign n1708 = x292 & n1065 ;
  assign n1909 = x420 & n4063 ;
  assign n1910 = n1708 | n1909 ;
  assign n4244 = ~n1908 ;
  assign n1911 = n4244 & n1910 ;
  assign n4245 = ~n2212 ;
  assign n2213 = n2210 & n4245 ;
  assign n2214 = n1911 | n2213 ;
  assign n4246 = ~n1910 ;
  assign n2206 = n1908 & n4246 ;
  assign n1778 = x163 & n3722 ;
  assign n1912 = x35 & n1606 ;
  assign n1913 = n1778 | n1912 ;
  assign n1108 = x419 & n4063 ;
  assign n1914 = x291 & n1065 ;
  assign n1915 = n1108 | n1914 ;
  assign n4247 = ~n1913 ;
  assign n1916 = n4247 & n1915 ;
  assign n1720 = x290 & n1065 ;
  assign n2195 = x418 & n4063 ;
  assign n2196 = n1720 | n2195 ;
  assign n1643 = x34 & n1606 ;
  assign n2197 = x162 & n3722 ;
  assign n2198 = n1643 | n2197 ;
  assign n4248 = ~n2196 ;
  assign n2202 = n4248 & n2198 ;
  assign n4249 = ~n1915 ;
  assign n2203 = n1913 & n4249 ;
  assign n2204 = n2202 | n2203 ;
  assign n1667 = x33 & n1606 ;
  assign n2185 = x161 & n3722 ;
  assign n2186 = n1667 | n2185 ;
  assign n1722 = x289 & n1065 ;
  assign n2187 = x417 & n4063 ;
  assign n2188 = n1722 | n2187 ;
  assign n4250 = ~n2186 ;
  assign n2194 = n4250 & n2188 ;
  assign n4251 = ~n2198 ;
  assign n2199 = n2196 & n4251 ;
  assign n2200 = n2194 | n2199 ;
  assign n4252 = ~n2188 ;
  assign n2189 = n2186 & n4252 ;
  assign n1092 = x416 & n4063 ;
  assign n2178 = x288 & n1065 ;
  assign n2179 = n1092 | n2178 ;
  assign n1634 = x32 & n1606 ;
  assign n2180 = x160 & n3722 ;
  assign n2181 = n1634 | n2180 ;
  assign n4253 = ~n2179 ;
  assign n2190 = n4253 & n2181 ;
  assign n2191 = n2189 | n2190 ;
  assign n4254 = ~n2181 ;
  assign n2182 = n2179 & n4254 ;
  assign n1093 = x415 & n4063 ;
  assign n2170 = x287 & n1065 ;
  assign n2171 = n1093 | n2170 ;
  assign n1810 = x159 & n3722 ;
  assign n2172 = x31 & n1606 ;
  assign n2173 = n1810 | n2172 ;
  assign n4255 = ~n2173 ;
  assign n2183 = n2171 & n4255 ;
  assign n2184 = n2182 | n2183 ;
  assign n4256 = ~n2171 ;
  assign n2174 = n4256 & n2173 ;
  assign n1713 = x286 & n1065 ;
  assign n2163 = x414 & n4063 ;
  assign n2164 = n1713 | n2163 ;
  assign n1629 = x30 & n1606 ;
  assign n2165 = x158 & n3722 ;
  assign n2166 = n1629 | n2165 ;
  assign n4257 = ~n2164 ;
  assign n2175 = n4257 & n2166 ;
  assign n2176 = n2174 | n2175 ;
  assign n1783 = x157 & n3722 ;
  assign n2153 = x29 & n1606 ;
  assign n2154 = n1783 | n2153 ;
  assign n1082 = x413 & n4063 ;
  assign n2155 = x285 & n1065 ;
  assign n2156 = n1082 | n2155 ;
  assign n4258 = ~n2154 ;
  assign n2162 = n4258 & n2156 ;
  assign n4259 = ~n2166 ;
  assign n2167 = n2164 & n4259 ;
  assign n2168 = n2162 | n2167 ;
  assign n4260 = ~n2156 ;
  assign n2157 = n2154 & n4260 ;
  assign n1684 = x284 & n1065 ;
  assign n2147 = x412 & n4063 ;
  assign n2148 = n1684 | n2147 ;
  assign n1809 = x156 & n3722 ;
  assign n2149 = x28 & n1606 ;
  assign n2150 = n1809 | n2149 ;
  assign n4261 = ~n2148 ;
  assign n2158 = n4261 & n2150 ;
  assign n2159 = n2157 | n2158 ;
  assign n1615 = x27 & n1606 ;
  assign n2139 = x155 & n3722 ;
  assign n2140 = n1615 | n2139 ;
  assign n1741 = x283 & n1065 ;
  assign n2141 = x411 & n4063 ;
  assign n2142 = n1741 | n2141 ;
  assign n4262 = ~n2140 ;
  assign n2146 = n4262 & n2142 ;
  assign n4263 = ~n2150 ;
  assign n2151 = n2148 & n4263 ;
  assign n2152 = n2146 | n2151 ;
  assign n1121 = x410 & n4063 ;
  assign n2130 = x282 & n1065 ;
  assign n2131 = n1121 | n2130 ;
  assign n1808 = x154 & n3722 ;
  assign n2132 = x26 & n1606 ;
  assign n2133 = n1808 | n2132 ;
  assign n4264 = ~n2131 ;
  assign n2138 = n4264 & n2133 ;
  assign n4265 = ~n2142 ;
  assign n2143 = n2140 & n4265 ;
  assign n2144 = n2138 | n2143 ;
  assign n4266 = ~n2133 ;
  assign n2134 = n2131 & n4266 ;
  assign n1126 = x409 & n4063 ;
  assign n2122 = x281 & n1065 ;
  assign n2123 = n1126 | n2122 ;
  assign n1665 = x25 & n1606 ;
  assign n2124 = x153 & n3722 ;
  assign n2125 = n1665 | n2124 ;
  assign n4267 = ~n2125 ;
  assign n2135 = n2123 & n4267 ;
  assign n2136 = n2134 | n2135 ;
  assign n1739 = x280 & n1065 ;
  assign n2114 = x408 & n4063 ;
  assign n2115 = n1739 | n2114 ;
  assign n1653 = x24 & n1606 ;
  assign n2116 = x152 & n3722 ;
  assign n2117 = n1653 | n2116 ;
  assign n4268 = ~n2115 ;
  assign n2121 = n4268 & n2117 ;
  assign n4269 = ~n2123 ;
  assign n2126 = n4269 & n2125 ;
  assign n2127 = n2121 | n2126 ;
  assign n4270 = ~n2117 ;
  assign n2118 = n2115 & n4270 ;
  assign n1683 = x279 & n1065 ;
  assign n2106 = x407 & n4063 ;
  assign n2107 = n1683 | n2106 ;
  assign n1764 = x151 & n3722 ;
  assign n2108 = x23 & n1606 ;
  assign n2109 = n1764 | n2108 ;
  assign n4271 = ~n2109 ;
  assign n2119 = n2107 & n4271 ;
  assign n2120 = n2118 | n2119 ;
  assign n4272 = ~n2107 ;
  assign n2110 = n4272 & n2109 ;
  assign n1112 = x406 & n4063 ;
  assign n2099 = x278 & n1065 ;
  assign n2100 = n1112 | n2099 ;
  assign n1664 = x22 & n1606 ;
  assign n2101 = x150 & n3722 ;
  assign n2102 = n1664 | n2101 ;
  assign n4273 = ~n2100 ;
  assign n2111 = n4273 & n2102 ;
  assign n2112 = n2110 | n2111 ;
  assign n1805 = x149 & n3722 ;
  assign n2089 = x21 & n1606 ;
  assign n2090 = n1805 | n2089 ;
  assign n1690 = x277 & n1065 ;
  assign n2091 = x405 & n4063 ;
  assign n2092 = n1690 | n2091 ;
  assign n4274 = ~n2090 ;
  assign n2098 = n4274 & n2092 ;
  assign n4275 = ~n2102 ;
  assign n2103 = n2100 & n4275 ;
  assign n2104 = n2098 | n2103 ;
  assign n4276 = ~n2092 ;
  assign n2093 = n2090 & n4276 ;
  assign n1089 = x404 & n4063 ;
  assign n2083 = x276 & n1065 ;
  assign n2084 = n1089 | n2083 ;
  assign n1756 = x148 & n3722 ;
  assign n2085 = x20 & n1606 ;
  assign n2086 = n1756 | n2085 ;
  assign n4277 = ~n2084 ;
  assign n2094 = n4277 & n2086 ;
  assign n2095 = n2093 | n2094 ;
  assign n1655 = x19 & n1606 ;
  assign n2074 = x147 & n3722 ;
  assign n2075 = n1655 | n2074 ;
  assign n1124 = x403 & n4063 ;
  assign n2076 = x275 & n1065 ;
  assign n2077 = n1124 | n2076 ;
  assign n4278 = ~n2075 ;
  assign n2082 = n4278 & n2077 ;
  assign n4279 = ~n2086 ;
  assign n2087 = n2084 & n4279 ;
  assign n2088 = n2082 | n2087 ;
  assign n4280 = ~n2077 ;
  assign n2078 = n2075 & n4280 ;
  assign n1735 = x274 & n1065 ;
  assign n2066 = x402 & n4063 ;
  assign n2067 = n1735 | n2066 ;
  assign n1804 = x146 & n3722 ;
  assign n2068 = x18 & n1606 ;
  assign n2069 = n1804 | n2068 ;
  assign n4281 = ~n2067 ;
  assign n2079 = n4281 & n2069 ;
  assign n2080 = n2078 | n2079 ;
  assign n4282 = ~n2069 ;
  assign n2070 = n2067 & n4282 ;
  assign n1732 = x273 & n1065 ;
  assign n2057 = x401 & n4063 ;
  assign n2058 = n1732 | n2057 ;
  assign n1654 = x17 & n1606 ;
  assign n2059 = x145 & n3722 ;
  assign n2060 = n1654 | n2059 ;
  assign n4283 = ~n2060 ;
  assign n2071 = n2058 & n4283 ;
  assign n2072 = n2070 | n2071 ;
  assign n4284 = ~n2058 ;
  assign n2061 = n4284 & n2060 ;
  assign n1796 = x144 & n3722 ;
  assign n2051 = x16 & n1606 ;
  assign n2052 = n1796 | n2051 ;
  assign n1110 = x400 & n4063 ;
  assign n2053 = x272 & n1065 ;
  assign n2054 = n1110 | n2053 ;
  assign n4285 = ~n2054 ;
  assign n2062 = n2052 & n4285 ;
  assign n2063 = n2061 | n2062 ;
  assign n1709 = x271 & n1065 ;
  assign n2042 = x399 & n4063 ;
  assign n2043 = n1709 | n2042 ;
  assign n1795 = x143 & n3722 ;
  assign n2044 = x15 & n1606 ;
  assign n2045 = n1795 | n2044 ;
  assign n4286 = ~n2045 ;
  assign n2050 = n2043 & n4286 ;
  assign n4287 = ~n2052 ;
  assign n2055 = n4287 & n2054 ;
  assign n2056 = n2050 | n2055 ;
  assign n1122 = x398 & n4063 ;
  assign n2035 = x270 & n1065 ;
  assign n2036 = n1122 | n2035 ;
  assign n1649 = x14 & n1606 ;
  assign n2037 = x142 & n3722 ;
  assign n2038 = n1649 | n2037 ;
  assign n4288 = ~n2036 ;
  assign n2046 = n4288 & n2038 ;
  assign n4289 = ~n2043 ;
  assign n2047 = n4289 & n2045 ;
  assign n2048 = n2046 | n2047 ;
  assign n1123 = x397 & n4063 ;
  assign n2025 = x269 & n1065 ;
  assign n2026 = n1123 | n2025 ;
  assign n1661 = x13 & n1606 ;
  assign n2027 = x141 & n3722 ;
  assign n2028 = n1661 | n2027 ;
  assign n4290 = ~n2028 ;
  assign n2029 = n2026 & n4290 ;
  assign n4291 = ~n2038 ;
  assign n2039 = n2036 & n4291 ;
  assign n2040 = n2029 | n2039 ;
  assign n4292 = ~n2026 ;
  assign n2030 = n4292 & n2028 ;
  assign n1719 = x268 & n1065 ;
  assign n2018 = x396 & n4063 ;
  assign n2019 = n1719 | n2018 ;
  assign n1803 = x140 & n3722 ;
  assign n2020 = x12 & n1606 ;
  assign n2021 = n1803 | n2020 ;
  assign n4293 = ~n2019 ;
  assign n2031 = n4293 & n2021 ;
  assign n2032 = n2030 | n2031 ;
  assign n4294 = ~n2021 ;
  assign n2022 = n2019 & n4294 ;
  assign n1119 = x395 & n4063 ;
  assign n2011 = x267 & n1065 ;
  assign n2012 = n1119 | n2011 ;
  assign n1801 = x139 & n3722 ;
  assign n2013 = x11 & n1606 ;
  assign n2014 = n1801 | n2013 ;
  assign n4295 = ~n2014 ;
  assign n2023 = n2012 & n4295 ;
  assign n2024 = n2022 | n2023 ;
  assign n1730 = x266 & n1065 ;
  assign n2002 = x394 & n4063 ;
  assign n2003 = n1730 | n2002 ;
  assign n1646 = x10 & n1606 ;
  assign n2004 = x138 & n3722 ;
  assign n2005 = n1646 | n2004 ;
  assign n4296 = ~n2003 ;
  assign n2010 = n4296 & n2005 ;
  assign n4297 = ~n2012 ;
  assign n2015 = n4297 & n2014 ;
  assign n2016 = n2010 | n2015 ;
  assign n4298 = ~n2005 ;
  assign n2006 = n2003 & n4298 ;
  assign n1728 = x265 & n1065 ;
  assign n1993 = x393 & n4063 ;
  assign n1994 = n1728 | n1993 ;
  assign n1794 = x137 & n3722 ;
  assign n1995 = x9 & n1606 ;
  assign n1996 = n1794 | n1995 ;
  assign n4299 = ~n1996 ;
  assign n2007 = n1994 & n4299 ;
  assign n2008 = n2006 | n2007 ;
  assign n1802 = x136 & n3722 ;
  assign n1987 = x8 & n1606 ;
  assign n1988 = n1802 | n1987 ;
  assign n1118 = x392 & n4063 ;
  assign n1989 = x264 & n1065 ;
  assign n1990 = n1118 | n1989 ;
  assign n4300 = ~n1990 ;
  assign n1997 = n1988 & n4300 ;
  assign n4301 = ~n1994 ;
  assign n1998 = n4301 & n1996 ;
  assign n1999 = n1997 | n1998 ;
  assign n1663 = x7 & n1606 ;
  assign n1979 = x135 & n3722 ;
  assign n1980 = n1663 | n1979 ;
  assign n1096 = x391 & n4063 ;
  assign n1981 = x263 & n1065 ;
  assign n1982 = n1096 | n1981 ;
  assign n4302 = ~n1980 ;
  assign n1984 = n4302 & n1982 ;
  assign n4303 = ~n1988 ;
  assign n1991 = n4303 & n1990 ;
  assign n1992 = n1984 | n1991 ;
  assign n1726 = x262 & n1065 ;
  assign n1971 = x390 & n4063 ;
  assign n1972 = n1726 | n1971 ;
  assign n1647 = x6 & n1606 ;
  assign n1973 = x134 & n3722 ;
  assign n1974 = n1647 | n1973 ;
  assign n4304 = ~n1972 ;
  assign n1976 = n4304 & n1974 ;
  assign n4305 = ~n1982 ;
  assign n1983 = n1980 & n4305 ;
  assign n1985 = n1976 | n1983 ;
  assign n1790 = x131 & n3722 ;
  assign n1945 = x3 & n1606 ;
  assign n1946 = n1790 | n1945 ;
  assign n1742 = n3840 & n1065 ;
  assign n1947 = x387 | n1065 ;
  assign n4306 = ~n1742 ;
  assign n1948 = n4306 & n1947 ;
  assign n4307 = ~n1948 ;
  assign n1949 = n1946 & n4307 ;
  assign n1131 = x386 | n1065 ;
  assign n2917 = n3841 & n1065 ;
  assign n4308 = ~n2917 ;
  assign n2918 = n1131 & n4308 ;
  assign n1675 = x2 & n1606 ;
  assign n2919 = x130 & n3722 ;
  assign n2920 = n1675 | n2919 ;
  assign n4309 = ~n2918 ;
  assign n2921 = n4309 & n2920 ;
  assign n2925 = n1949 | n2921 ;
  assign n4310 = ~x256 ;
  assign n1747 = n4310 & n1065 ;
  assign n2908 = x384 | n1065 ;
  assign n4311 = ~n1747 ;
  assign n2909 = n4311 & n2908 ;
  assign n4312 = ~n2909 ;
  assign n2910 = n2907 & n4312 ;
  assign n1725 = n3842 & n1065 ;
  assign n2911 = x385 | n1065 ;
  assign n4313 = ~n1725 ;
  assign n2912 = n4313 & n2911 ;
  assign n1784 = x129 & n3722 ;
  assign n2913 = x1 & n1606 ;
  assign n2914 = n1784 | n2913 ;
  assign n4314 = ~n2912 ;
  assign n2915 = n4314 & n2914 ;
  assign n2916 = n2910 | n2915 ;
  assign n4315 = ~n2914 ;
  assign n2922 = n2912 & n4315 ;
  assign n4316 = ~n2920 ;
  assign n2923 = n2918 & n4316 ;
  assign n2924 = n2922 | n2923 ;
  assign n4317 = ~n2924 ;
  assign n2926 = n2916 & n4317 ;
  assign n2927 = n2925 | n2926 ;
  assign n1788 = x131 | n1606 ;
  assign n1936 = n3520 & n1606 ;
  assign n4318 = ~n1936 ;
  assign n1937 = n1788 & n4318 ;
  assign n1738 = x259 & n1065 ;
  assign n1938 = x387 & n4063 ;
  assign n1939 = n1738 | n1938 ;
  assign n4319 = ~n1937 ;
  assign n1940 = n4319 & n1939 ;
  assign n1100 = x388 & n4063 ;
  assign n2928 = x260 & n1065 ;
  assign n2929 = n1100 | n2928 ;
  assign n1676 = n3519 & n1606 ;
  assign n2931 = x132 | n1606 ;
  assign n4320 = ~n1676 ;
  assign n2932 = n4320 & n2931 ;
  assign n4321 = ~n2932 ;
  assign n2933 = n2929 & n4321 ;
  assign n2934 = n1940 | n2933 ;
  assign n4322 = ~n2934 ;
  assign n2935 = n2927 & n4322 ;
  assign n4323 = ~n2929 ;
  assign n2936 = n4323 & n2932 ;
  assign n1807 = x133 | n1606 ;
  assign n1966 = n3525 & n1606 ;
  assign n4324 = ~n1966 ;
  assign n1967 = n1807 & n4324 ;
  assign n1125 = x389 & n4063 ;
  assign n1968 = x261 & n1065 ;
  assign n1969 = n1125 | n1968 ;
  assign n4325 = ~n1969 ;
  assign n2937 = n1967 & n4325 ;
  assign n2938 = n2936 | n2937 ;
  assign n2939 = n2935 | n2938 ;
  assign n4326 = ~n1974 ;
  assign n1975 = n1972 & n4326 ;
  assign n1799 = x133 & n3722 ;
  assign n1958 = x5 & n1606 ;
  assign n1959 = n1799 | n1958 ;
  assign n1117 = x389 | n1065 ;
  assign n1960 = n3837 & n1065 ;
  assign n4327 = ~n1960 ;
  assign n1961 = n1117 & n4327 ;
  assign n4328 = ~n1959 ;
  assign n2940 = n4328 & n1961 ;
  assign n2941 = n1975 | n2940 ;
  assign n4329 = ~n2941 ;
  assign n2942 = n2939 & n4329 ;
  assign n2943 = n1985 | n2942 ;
  assign n4330 = ~n1992 ;
  assign n2944 = n4330 & n2943 ;
  assign n2945 = n1999 | n2944 ;
  assign n4331 = ~n2008 ;
  assign n2946 = n4331 & n2945 ;
  assign n2947 = n2016 | n2946 ;
  assign n4332 = ~n2024 ;
  assign n2948 = n4332 & n2947 ;
  assign n2949 = n2032 | n2948 ;
  assign n4333 = ~n2040 ;
  assign n2950 = n4333 & n2949 ;
  assign n2951 = n2048 | n2950 ;
  assign n4334 = ~n2056 ;
  assign n2952 = n4334 & n2951 ;
  assign n2953 = n2063 | n2952 ;
  assign n4335 = ~n2072 ;
  assign n2954 = n4335 & n2953 ;
  assign n2955 = n2080 | n2954 ;
  assign n4336 = ~n2088 ;
  assign n2956 = n4336 & n2955 ;
  assign n2957 = n2095 | n2956 ;
  assign n4337 = ~n2104 ;
  assign n2958 = n4337 & n2957 ;
  assign n2959 = n2112 | n2958 ;
  assign n4338 = ~n2120 ;
  assign n2960 = n4338 & n2959 ;
  assign n2961 = n2127 | n2960 ;
  assign n4339 = ~n2136 ;
  assign n2962 = n4339 & n2961 ;
  assign n2963 = n2144 | n2962 ;
  assign n4340 = ~n2152 ;
  assign n2964 = n4340 & n2963 ;
  assign n2965 = n2159 | n2964 ;
  assign n4341 = ~n2168 ;
  assign n2966 = n4341 & n2965 ;
  assign n2967 = n2176 | n2966 ;
  assign n4342 = ~n2184 ;
  assign n2968 = n4342 & n2967 ;
  assign n2969 = n2191 | n2968 ;
  assign n4343 = ~n2200 ;
  assign n2970 = n4343 & n2969 ;
  assign n2971 = n2204 | n2970 ;
  assign n4344 = ~n1916 ;
  assign n2972 = n4344 & n2971 ;
  assign n2973 = n2206 | n2972 ;
  assign n4345 = ~n2214 ;
  assign n2974 = n4345 & n2973 ;
  assign n2975 = n2222 | n2974 ;
  assign n4346 = ~n2226 ;
  assign n2976 = n4346 & n2975 ;
  assign n2977 = n1906 | n2976 ;
  assign n4347 = ~n1901 ;
  assign n2978 = n4347 & n2977 ;
  assign n2979 = n2236 | n2978 ;
  assign n4348 = ~n2244 ;
  assign n2980 = n4348 & n2979 ;
  assign n2981 = n2251 | n2980 ;
  assign n4349 = ~n2260 ;
  assign n2982 = n4349 & n2981 ;
  assign n2983 = n2264 | n2982 ;
  assign n4350 = ~n1896 ;
  assign n2984 = n4350 & n2983 ;
  assign n2985 = n2266 | n2984 ;
  assign n4351 = ~n2274 ;
  assign n2986 = n4351 & n2985 ;
  assign n2987 = n2282 | n2986 ;
  assign n4352 = ~n2290 ;
  assign n2988 = n4352 & n2987 ;
  assign n2989 = n2297 | n2988 ;
  assign n4353 = ~n2306 ;
  assign n2990 = n4353 & n2989 ;
  assign n2991 = n2314 | n2990 ;
  assign n4354 = ~n2322 ;
  assign n2992 = n4354 & n2991 ;
  assign n2993 = n2329 | n2992 ;
  assign n4355 = ~n2338 ;
  assign n2994 = n4355 & n2993 ;
  assign n2995 = n2346 | n2994 ;
  assign n4356 = ~n2354 ;
  assign n2996 = n4356 & n2995 ;
  assign n2997 = n2361 | n2996 ;
  assign n4357 = ~n2366 ;
  assign n2998 = n4357 & n2997 ;
  assign n2999 = n1886 | n2998 ;
  assign n4358 = ~n1881 ;
  assign n3000 = n4358 & n2999 ;
  assign n3001 = n2375 | n3000 ;
  assign n4359 = ~n2384 ;
  assign n3002 = n4359 & n3001 ;
  assign n3003 = n2388 | n3002 ;
  assign n4360 = ~n1876 ;
  assign n3004 = n4360 & n3003 ;
  assign n3005 = n2390 | n3004 ;
  assign n4361 = ~n2398 ;
  assign n3006 = n4361 & n3005 ;
  assign n3007 = n2402 | n3006 ;
  assign n4362 = ~n1866 ;
  assign n3008 = n4362 & n3007 ;
  assign n3009 = n2404 | n3008 ;
  assign n4363 = ~n2412 ;
  assign n3010 = n4363 & n3009 ;
  assign n3011 = n2420 | n3010 ;
  assign n4364 = ~n2428 ;
  assign n3012 = n4364 & n3011 ;
  assign n3013 = n2435 | n3012 ;
  assign n4365 = ~n2444 ;
  assign n3014 = n4365 & n3013 ;
  assign n3015 = n2452 | n3014 ;
  assign n4366 = ~n2456 ;
  assign n3016 = n4366 & n3015 ;
  assign n3017 = n1856 | n3016 ;
  assign n4367 = ~n1851 ;
  assign n3018 = n4367 & n3017 ;
  assign n3019 = n2466 | n3018 ;
  assign n4368 = ~n2474 ;
  assign n3020 = n4368 & n3019 ;
  assign n3021 = n2477 | n3020 ;
  assign n4369 = ~n1846 ;
  assign n3022 = n4369 & n3021 ;
  assign n3023 = n1841 | n3022 ;
  assign n4370 = ~n2487 ;
  assign n3024 = n4370 & n3023 ;
  assign n3025 = n2494 | n3024 ;
  assign n4371 = ~n2499 ;
  assign n3026 = n4371 & n3025 ;
  assign n3027 = n1835 | n3026 ;
  assign n4372 = ~n1830 ;
  assign n3028 = n4372 & n3027 ;
  assign n3029 = n2508 | n3028 ;
  assign n4373 = ~n2513 ;
  assign n3030 = n4373 & n3029 ;
  assign n3031 = n1825 | n3030 ;
  assign n4374 = ~n1820 ;
  assign n3032 = n4374 & n3031 ;
  assign n3033 = n2522 | n3032 ;
  assign n4375 = ~n2531 ;
  assign n3034 = n4375 & n3033 ;
  assign n3035 = n2539 | n3034 ;
  assign n4376 = ~n2547 ;
  assign n3036 = n4376 & n3035 ;
  assign n3037 = n2554 | n3036 ;
  assign n4377 = ~n2563 ;
  assign n3038 = n4377 & n3037 ;
  assign n3039 = n2571 | n3038 ;
  assign n4378 = ~n2579 ;
  assign n3040 = n4378 & n3039 ;
  assign n3041 = n2586 | n3040 ;
  assign n4379 = ~n2595 ;
  assign n3042 = n4379 & n3041 ;
  assign n3043 = n2603 | n3042 ;
  assign n4380 = ~n2611 ;
  assign n3044 = n4380 & n3043 ;
  assign n3045 = n2618 | n3044 ;
  assign n4381 = ~n2627 ;
  assign n3046 = n4381 & n3045 ;
  assign n3047 = n2635 | n3046 ;
  assign n4382 = ~n2643 ;
  assign n3048 = n4382 & n3047 ;
  assign n3049 = n2650 | n3048 ;
  assign n4383 = ~n2659 ;
  assign n3050 = n4383 & n3049 ;
  assign n3051 = n2667 | n3050 ;
  assign n4384 = ~n2675 ;
  assign n3052 = n4384 & n3051 ;
  assign n3053 = n2682 | n3052 ;
  assign n4385 = ~n2691 ;
  assign n3054 = n4385 & n3053 ;
  assign n3055 = n2699 | n3054 ;
  assign n4386 = ~n2707 ;
  assign n3056 = n4386 & n3055 ;
  assign n3057 = n2714 | n3056 ;
  assign n4387 = ~n2723 ;
  assign n3058 = n4387 & n3057 ;
  assign n3059 = n2731 | n3058 ;
  assign n4388 = ~n2739 ;
  assign n3060 = n4388 & n3059 ;
  assign n3061 = n2742 | n3060 ;
  assign n4389 = ~n1815 ;
  assign n3062 = n4389 & n3061 ;
  assign n3063 = n1680 | n3062 ;
  assign n4390 = ~n2752 ;
  assign n3064 = n4390 & n3063 ;
  assign n3065 = n2759 | n3064 ;
  assign n4391 = ~n2768 ;
  assign n3066 = n4391 & n3065 ;
  assign n3067 = n2776 | n3066 ;
  assign n4392 = ~n2784 ;
  assign n3068 = n4392 & n3067 ;
  assign n3069 = n2791 | n3068 ;
  assign n4393 = ~n2800 ;
  assign n3070 = n4393 & n3069 ;
  assign n3071 = n2808 | n3070 ;
  assign n4394 = ~n2816 ;
  assign n3072 = n4394 & n3071 ;
  assign n3073 = n2823 | n3072 ;
  assign n4395 = ~n2828 ;
  assign n3074 = n4395 & n3073 ;
  assign n3075 = n3303 | n3074 ;
  assign n3126 = n2907 & n3075 ;
  assign n1734 = x256 & n1065 ;
  assign n1919 = x384 & n4063 ;
  assign n1920 = n1734 | n1919 ;
  assign n4396 = ~n3075 ;
  assign n3382 = n1920 & n4396 ;
  assign n513 = n3126 | n3382 ;
  assign n1707 = x257 & n1065 ;
  assign n1921 = x385 & n4063 ;
  assign n1922 = n1707 | n1921 ;
  assign n1115 = x388 | n1065 ;
  assign n1950 = n3839 & n1065 ;
  assign n4397 = ~n1950 ;
  assign n1951 = n1115 & n4397 ;
  assign n1641 = x4 & n1606 ;
  assign n1952 = x132 & n3722 ;
  assign n1953 = n1641 | n1952 ;
  assign n4398 = ~n1951 ;
  assign n1954 = n4398 & n1953 ;
  assign n4399 = ~n1961 ;
  assign n1962 = n1959 & n4399 ;
  assign n1963 = n1954 | n1962 ;
  assign n4400 = ~x0 ;
  assign n1631 = n4400 & n1606 ;
  assign n1917 = x128 | n1606 ;
  assign n4401 = ~n1631 ;
  assign n1918 = n4401 & n1917 ;
  assign n4402 = ~n1920 ;
  assign n1926 = n1918 & n4402 ;
  assign n1777 = x129 | n1606 ;
  assign n1923 = n3515 & n1606 ;
  assign n4403 = ~n1923 ;
  assign n1924 = n1777 & n4403 ;
  assign n4404 = ~n1922 ;
  assign n1927 = n4404 & n1924 ;
  assign n1928 = n1926 | n1927 ;
  assign n4405 = ~n1924 ;
  assign n1925 = n1922 & n4405 ;
  assign n1111 = x386 & n4063 ;
  assign n1929 = x258 & n1065 ;
  assign n1930 = n1111 | n1929 ;
  assign n1657 = n3513 & n1606 ;
  assign n1931 = x130 | n1606 ;
  assign n4406 = ~n1657 ;
  assign n1932 = n4406 & n1931 ;
  assign n4407 = ~n1932 ;
  assign n1933 = n1930 & n4407 ;
  assign n1934 = n1925 | n1933 ;
  assign n4408 = ~n1934 ;
  assign n1935 = n1928 & n4408 ;
  assign n4409 = ~n1930 ;
  assign n1941 = n4409 & n1932 ;
  assign n4410 = ~n1939 ;
  assign n1942 = n1937 & n4410 ;
  assign n1943 = n1941 | n1942 ;
  assign n1944 = n1935 | n1943 ;
  assign n4411 = ~n1946 ;
  assign n1955 = n4411 & n1948 ;
  assign n4412 = ~n1953 ;
  assign n1956 = n1951 & n4412 ;
  assign n1957 = n1955 | n1956 ;
  assign n4413 = ~n1957 ;
  assign n1964 = n1944 & n4413 ;
  assign n1965 = n1963 | n1964 ;
  assign n4414 = ~n1967 ;
  assign n1970 = n4414 & n1969 ;
  assign n1977 = n1970 | n1975 ;
  assign n4415 = ~n1977 ;
  assign n1978 = n1965 & n4415 ;
  assign n1986 = n1978 | n1985 ;
  assign n2000 = n1986 & n4330 ;
  assign n2001 = n1999 | n2000 ;
  assign n2009 = n2001 & n4331 ;
  assign n2017 = n2009 | n2016 ;
  assign n2033 = n2017 & n4332 ;
  assign n2034 = n2032 | n2033 ;
  assign n2041 = n2034 & n4333 ;
  assign n2049 = n2041 | n2048 ;
  assign n2064 = n2049 & n4334 ;
  assign n2065 = n2063 | n2064 ;
  assign n2073 = n2065 & n4335 ;
  assign n2081 = n2073 | n2080 ;
  assign n2096 = n2081 & n4336 ;
  assign n2097 = n2095 | n2096 ;
  assign n2105 = n2097 & n4337 ;
  assign n2113 = n2105 | n2112 ;
  assign n2128 = n2113 & n4338 ;
  assign n2129 = n2127 | n2128 ;
  assign n2137 = n2129 & n4339 ;
  assign n2145 = n2137 | n2144 ;
  assign n2160 = n2145 & n4340 ;
  assign n2161 = n2159 | n2160 ;
  assign n2169 = n2161 & n4341 ;
  assign n2177 = n2169 | n2176 ;
  assign n2192 = n2177 & n4342 ;
  assign n2193 = n2191 | n2192 ;
  assign n2201 = n2193 & n4343 ;
  assign n2205 = n2201 | n2204 ;
  assign n2207 = n4344 & n2205 ;
  assign n2208 = n2206 | n2207 ;
  assign n2215 = n2208 & n4345 ;
  assign n2223 = n2215 | n2222 ;
  assign n2227 = n2223 & n4346 ;
  assign n2228 = n1906 | n2227 ;
  assign n2229 = n4347 & n2228 ;
  assign n2237 = n2229 | n2236 ;
  assign n2252 = n2237 & n4348 ;
  assign n2253 = n2251 | n2252 ;
  assign n2261 = n2253 & n4349 ;
  assign n2265 = n2261 | n2264 ;
  assign n2267 = n4350 & n2265 ;
  assign n2268 = n2266 | n2267 ;
  assign n2275 = n2268 & n4351 ;
  assign n2283 = n2275 | n2282 ;
  assign n2298 = n2283 & n4352 ;
  assign n2299 = n2297 | n2298 ;
  assign n2307 = n2299 & n4353 ;
  assign n2315 = n2307 | n2314 ;
  assign n2330 = n2315 & n4354 ;
  assign n2331 = n2329 | n2330 ;
  assign n2339 = n2331 & n4355 ;
  assign n2347 = n2339 | n2346 ;
  assign n2362 = n2347 & n4356 ;
  assign n2363 = n2361 | n2362 ;
  assign n2367 = n2363 & n4357 ;
  assign n2368 = n1886 | n2367 ;
  assign n2376 = n4358 & n2368 ;
  assign n2377 = n2375 | n2376 ;
  assign n2385 = n2377 & n4359 ;
  assign n2389 = n2385 | n2388 ;
  assign n2391 = n4360 & n2389 ;
  assign n2392 = n2390 | n2391 ;
  assign n2399 = n2392 & n4361 ;
  assign n2403 = n2399 | n2402 ;
  assign n2405 = n4362 & n2403 ;
  assign n2406 = n2404 | n2405 ;
  assign n2413 = n2406 & n4363 ;
  assign n2421 = n2413 | n2420 ;
  assign n2436 = n2421 & n4364 ;
  assign n2437 = n2435 | n2436 ;
  assign n2445 = n2437 & n4365 ;
  assign n2453 = n2445 | n2452 ;
  assign n2457 = n2453 & n4366 ;
  assign n2458 = n1856 | n2457 ;
  assign n2459 = n4367 & n2458 ;
  assign n2467 = n2459 | n2466 ;
  assign n2478 = n2467 & n4368 ;
  assign n2479 = n2477 | n2478 ;
  assign n2480 = n4369 & n2479 ;
  assign n2481 = n1841 | n2480 ;
  assign n2495 = n2481 & n4370 ;
  assign n2496 = n2494 | n2495 ;
  assign n2500 = n2496 & n4371 ;
  assign n2501 = n1835 | n2500 ;
  assign n2509 = n4372 & n2501 ;
  assign n2510 = n2508 | n2509 ;
  assign n2514 = n2510 & n4373 ;
  assign n2515 = n1825 | n2514 ;
  assign n2523 = n4374 & n2515 ;
  assign n2524 = n2522 | n2523 ;
  assign n2532 = n2524 & n4375 ;
  assign n2540 = n2532 | n2539 ;
  assign n2555 = n2540 & n4376 ;
  assign n2556 = n2554 | n2555 ;
  assign n2564 = n2556 & n4377 ;
  assign n2572 = n2564 | n2571 ;
  assign n2587 = n2572 & n4378 ;
  assign n2588 = n2586 | n2587 ;
  assign n2596 = n2588 & n4379 ;
  assign n2604 = n2596 | n2603 ;
  assign n2619 = n2604 & n4380 ;
  assign n2620 = n2618 | n2619 ;
  assign n2628 = n2620 & n4381 ;
  assign n2636 = n2628 | n2635 ;
  assign n2651 = n2636 & n4382 ;
  assign n2652 = n2650 | n2651 ;
  assign n2660 = n2652 & n4383 ;
  assign n2668 = n2660 | n2667 ;
  assign n2683 = n2668 & n4384 ;
  assign n2684 = n2682 | n2683 ;
  assign n2692 = n2684 & n4385 ;
  assign n2700 = n2692 | n2699 ;
  assign n2715 = n2700 & n4386 ;
  assign n2716 = n2714 | n2715 ;
  assign n2724 = n2716 & n4387 ;
  assign n2732 = n2724 | n2731 ;
  assign n2743 = n2732 & n4388 ;
  assign n2744 = n2742 | n2743 ;
  assign n2745 = n4389 & n2744 ;
  assign n2746 = n1680 | n2745 ;
  assign n2760 = n2746 & n4390 ;
  assign n2761 = n2759 | n2760 ;
  assign n2769 = n2761 & n4391 ;
  assign n2777 = n2769 | n2776 ;
  assign n2792 = n2777 & n4392 ;
  assign n2793 = n2791 | n2792 ;
  assign n2801 = n2793 & n4393 ;
  assign n2809 = n2801 | n2808 ;
  assign n2824 = n2809 & n4394 ;
  assign n2825 = n2823 | n2824 ;
  assign n2829 = n2825 & n4395 ;
  assign n2830 = n3303 | n2829 ;
  assign n642 = ~n2830 ;
  assign n2905 = n1922 & n642 ;
  assign n3380 = n2830 & n2914 ;
  assign n514 = n2905 | n3380 ;
  assign n2863 = n1930 & n642 ;
  assign n3378 = n2830 & n2920 ;
  assign n515 = n2863 | n3378 ;
  assign n3127 = n1946 & n3075 ;
  assign n3228 = n1939 & n4396 ;
  assign n516 = n3127 | n3228 ;
  assign n2930 = n642 & n2929 ;
  assign n3376 = n1953 & n2830 ;
  assign n517 = n2930 | n3376 ;
  assign n3125 = n1959 & n3075 ;
  assign n3226 = n1969 & n4396 ;
  assign n518 = n3125 | n3226 ;
  assign n2904 = n1972 & n642 ;
  assign n3374 = n1974 & n2830 ;
  assign n519 = n2904 | n3374 ;
  assign n3124 = n1980 & n3075 ;
  assign n3224 = n1982 & n4396 ;
  assign n520 = n3124 | n3224 ;
  assign n3123 = n1988 & n3075 ;
  assign n3222 = n1990 & n4396 ;
  assign n521 = n3123 | n3222 ;
  assign n2903 = n1994 & n642 ;
  assign n3372 = n1996 & n2830 ;
  assign n522 = n2903 | n3372 ;
  assign n2902 = n2003 & n642 ;
  assign n3370 = n2005 & n2830 ;
  assign n523 = n2902 | n3370 ;
  assign n2901 = n2012 & n642 ;
  assign n3368 = n2014 & n2830 ;
  assign n524 = n2901 | n3368 ;
  assign n2900 = n2019 & n642 ;
  assign n3366 = n2021 & n2830 ;
  assign n525 = n2900 | n3366 ;
  assign n2899 = n2026 & n642 ;
  assign n3364 = n2028 & n2830 ;
  assign n526 = n2899 | n3364 ;
  assign n2898 = n2036 & n642 ;
  assign n3362 = n2038 & n2830 ;
  assign n527 = n2898 | n3362 ;
  assign n2849 = n2043 & n642 ;
  assign n3360 = n2045 & n2830 ;
  assign n528 = n2849 | n3360 ;
  assign n3122 = n2052 & n3075 ;
  assign n3220 = n2054 & n4396 ;
  assign n529 = n3122 | n3220 ;
  assign n2896 = n2058 & n642 ;
  assign n3358 = n2060 & n2830 ;
  assign n530 = n2896 | n3358 ;
  assign n2897 = n2067 & n642 ;
  assign n3356 = n2069 & n2830 ;
  assign n531 = n2897 | n3356 ;
  assign n3105 = n2075 & n3075 ;
  assign n3218 = n2077 & n4396 ;
  assign n532 = n3105 | n3218 ;
  assign n2893 = n2084 & n642 ;
  assign n3354 = n2086 & n2830 ;
  assign n533 = n2893 | n3354 ;
  assign n3117 = n2090 & n3075 ;
  assign n3216 = n2092 & n4396 ;
  assign n534 = n3117 | n3216 ;
  assign n2853 = n2100 & n642 ;
  assign n3352 = n2102 & n2830 ;
  assign n535 = n2853 | n3352 ;
  assign n2895 = n2107 & n642 ;
  assign n3350 = n2109 & n2830 ;
  assign n536 = n2895 | n3350 ;
  assign n2894 = n2115 & n642 ;
  assign n3348 = n2117 & n2830 ;
  assign n537 = n2894 | n3348 ;
  assign n2848 = n2123 & n642 ;
  assign n3346 = n2125 & n2830 ;
  assign n538 = n2848 | n3346 ;
  assign n2841 = n2131 & n642 ;
  assign n3344 = n2133 & n2830 ;
  assign n539 = n2841 | n3344 ;
  assign n3121 = n2140 & n3075 ;
  assign n3214 = n2142 & n4396 ;
  assign n540 = n3121 | n3214 ;
  assign n2858 = n2148 & n642 ;
  assign n3342 = n2150 & n2830 ;
  assign n541 = n2858 | n3342 ;
  assign n3108 = n2154 & n3075 ;
  assign n3212 = n2156 & n4396 ;
  assign n542 = n3108 | n3212 ;
  assign n2881 = n2164 & n642 ;
  assign n3340 = n2166 & n2830 ;
  assign n543 = n2881 | n3340 ;
  assign n2834 = n2171 & n642 ;
  assign n3338 = n2173 & n2830 ;
  assign n544 = n2834 | n3338 ;
  assign n2831 = n2179 & n642 ;
  assign n3336 = n2181 & n2830 ;
  assign n545 = n2831 | n3336 ;
  assign n3087 = n2186 & n3075 ;
  assign n3210 = n2188 & n4396 ;
  assign n546 = n3087 | n3210 ;
  assign n2872 = n2196 & n642 ;
  assign n3334 = n2198 & n2830 ;
  assign n547 = n2872 | n3334 ;
  assign n3093 = n1913 & n3075 ;
  assign n3208 = n1915 & n4396 ;
  assign n548 = n3093 | n3208 ;
  assign n3120 = n1908 & n3075 ;
  assign n3206 = n1910 & n4396 ;
  assign n549 = n3120 | n3206 ;
  assign n2832 = n2210 & n642 ;
  assign n3332 = n2212 & n2830 ;
  assign n550 = n2832 | n3332 ;
  assign n3083 = n2217 & n3075 ;
  assign n3204 = n2219 & n4396 ;
  assign n551 = n3083 | n3204 ;
  assign n2889 = n1903 & n642 ;
  assign n3330 = n1905 & n2830 ;
  assign n552 = n2889 | n3330 ;
  assign n2833 = n1898 & n642 ;
  assign n3328 = n1900 & n2830 ;
  assign n553 = n2833 | n3328 ;
  assign n2837 = n2231 & n642 ;
  assign n3326 = n2233 & n2830 ;
  assign n554 = n2837 | n3326 ;
  assign n2838 = n2240 & n642 ;
  assign n3324 = n2242 & n2830 ;
  assign n555 = n2838 | n3324 ;
  assign n2891 = n2247 & n642 ;
  assign n3322 = n2249 & n2830 ;
  assign n556 = n2891 | n3322 ;
  assign n3119 = n2255 & n3075 ;
  assign n3202 = n2257 & n4396 ;
  assign n557 = n3119 | n3202 ;
  assign n2864 = n1893 & n642 ;
  assign n3320 = n1895 & n2830 ;
  assign n558 = n2864 | n3320 ;
  assign n2843 = n1888 & n642 ;
  assign n3318 = n1890 & n2830 ;
  assign n559 = n2843 | n3318 ;
  assign n2839 = n2270 & n642 ;
  assign n3316 = n2272 & n2830 ;
  assign n560 = n2839 | n3316 ;
  assign n2845 = n2277 & n642 ;
  assign n3314 = n2279 & n2830 ;
  assign n561 = n2845 | n3314 ;
  assign n3118 = n2285 & n3075 ;
  assign n3200 = n2287 & n4396 ;
  assign n562 = n3118 | n3200 ;
  assign n2846 = n2293 & n642 ;
  assign n3312 = n2295 & n2830 ;
  assign n563 = n2846 | n3312 ;
  assign n3101 = n2301 & n3075 ;
  assign n3198 = n2303 & n4396 ;
  assign n564 = n3101 | n3198 ;
  assign n2852 = n2310 & n642 ;
  assign n3310 = n2312 & n2830 ;
  assign n565 = n2852 | n3310 ;
  assign n2847 = n2317 & n642 ;
  assign n3308 = n2319 & n2830 ;
  assign n566 = n2847 | n3308 ;
  assign n2835 = n2324 & n642 ;
  assign n3306 = n2326 & n2830 ;
  assign n567 = n2835 | n3306 ;
  assign n3116 = n2334 & n3075 ;
  assign n3196 = n2336 & n4396 ;
  assign n568 = n3116 | n3196 ;
  assign n2850 = n2341 & n642 ;
  assign n3304 = n2343 & n2830 ;
  assign n569 = n2850 | n3304 ;
  assign n3082 = n2350 & n3075 ;
  assign n3194 = n2352 & n4396 ;
  assign n570 = n3082 | n3194 ;
  assign n3115 = n2357 & n3075 ;
  assign n3192 = n2359 & n4396 ;
  assign n571 = n3115 | n3192 ;
  assign n2842 = n1883 & n642 ;
  assign n3302 = n1885 & n2830 ;
  assign n572 = n2842 | n3302 ;
  assign n2869 = n1878 & n642 ;
  assign n3300 = n1880 & n2830 ;
  assign n573 = n2869 | n3300 ;
  assign n3114 = n2370 & n3075 ;
  assign n3190 = n2372 & n4396 ;
  assign n574 = n3114 | n3190 ;
  assign n3085 = n2380 & n3075 ;
  assign n3188 = n2382 & n4396 ;
  assign n575 = n3085 | n3188 ;
  assign n3113 = n1873 & n3075 ;
  assign n3186 = n1875 & n4396 ;
  assign n576 = n3113 | n3186 ;
  assign n3089 = n1868 & n3075 ;
  assign n3184 = n1870 & n4396 ;
  assign n577 = n3089 | n3184 ;
  assign n3079 = n2394 & n3075 ;
  assign n3182 = n2396 & n4396 ;
  assign n578 = n3079 | n3182 ;
  assign n3076 = n1863 & n3075 ;
  assign n3180 = n1865 & n4396 ;
  assign n579 = n3076 | n3180 ;
  assign n3077 = n1858 & n3075 ;
  assign n3178 = n1860 & n4396 ;
  assign n580 = n3077 | n3178 ;
  assign n3084 = n2408 & n3075 ;
  assign n3176 = n2410 & n4396 ;
  assign n581 = n3084 | n3176 ;
  assign n2873 = n2415 & n642 ;
  assign n3298 = n2417 & n2830 ;
  assign n582 = n2873 | n3298 ;
  assign n2854 = n2423 & n642 ;
  assign n3296 = n2425 & n2830 ;
  assign n583 = n2854 | n3296 ;
  assign n3098 = n2430 & n3075 ;
  assign n3174 = n2432 & n4396 ;
  assign n584 = n3098 | n3174 ;
  assign n3094 = n2439 & n3075 ;
  assign n3172 = n2441 & n4396 ;
  assign n585 = n3094 | n3172 ;
  assign n3081 = n2448 & n3075 ;
  assign n3170 = n2450 & n4396 ;
  assign n586 = n3081 | n3170 ;
  assign n2851 = n1853 & n642 ;
  assign n3294 = n1855 & n2830 ;
  assign n587 = n2851 | n3294 ;
  assign n2879 = n1848 & n642 ;
  assign n3292 = n1850 & n2830 ;
  assign n588 = n2879 | n3292 ;
  assign n3080 = n2461 & n3075 ;
  assign n3168 = n2463 & n4396 ;
  assign n589 = n3080 | n3168 ;
  assign n3086 = n2470 & n3075 ;
  assign n3166 = n2472 & n4396 ;
  assign n590 = n3086 | n3166 ;
  assign n2860 = n1843 & n642 ;
  assign n3290 = n1845 & n2830 ;
  assign n591 = n2860 | n3290 ;
  assign n2866 = n1837 & n642 ;
  assign n3288 = n1839 & n2830 ;
  assign n592 = n2866 | n3288 ;
  assign n3088 = n2483 & n3075 ;
  assign n3164 = n2485 & n4396 ;
  assign n593 = n3088 | n3164 ;
  assign n3078 = n2489 & n3075 ;
  assign n3162 = n2491 & n4396 ;
  assign n594 = n3078 | n3162 ;
  assign n3090 = n1832 & n3075 ;
  assign n3160 = n1834 & n4396 ;
  assign n595 = n3090 | n3160 ;
  assign n3091 = n1827 & n3075 ;
  assign n3158 = n1829 & n4396 ;
  assign n596 = n3091 | n3158 ;
  assign n3092 = n2504 & n3075 ;
  assign n3156 = n2506 & n4396 ;
  assign n597 = n3092 | n3156 ;
  assign n2844 = n1822 & n642 ;
  assign n3286 = n1824 & n2830 ;
  assign n598 = n2844 | n3286 ;
  assign n2890 = n1817 & n642 ;
  assign n3284 = n1819 & n2830 ;
  assign n599 = n2890 | n3284 ;
  assign n3095 = n2517 & n3075 ;
  assign n3154 = n2519 & n4396 ;
  assign n600 = n3095 | n3154 ;
  assign n2856 = n2527 & n642 ;
  assign n3282 = n2529 & n2830 ;
  assign n601 = n2856 | n3282 ;
  assign n3110 = n2534 & n3075 ;
  assign n3152 = n2536 & n4396 ;
  assign n602 = n3110 | n3152 ;
  assign n2880 = n2543 & n642 ;
  assign n3280 = n2545 & n2830 ;
  assign n603 = n2880 | n3280 ;
  assign n2888 = n2549 & n642 ;
  assign n3278 = n2551 & n2830 ;
  assign n604 = n2888 | n3278 ;
  assign n3102 = n2558 & n3075 ;
  assign n3150 = n2560 & n4396 ;
  assign n605 = n3102 | n3150 ;
  assign n2892 = n2566 & n642 ;
  assign n3276 = n2568 & n2830 ;
  assign n606 = n2892 | n3276 ;
  assign n3112 = n2575 & n3075 ;
  assign n3148 = n2577 & n4396 ;
  assign n607 = n3112 | n3148 ;
  assign n3109 = n2582 & n3075 ;
  assign n3146 = n2584 & n4396 ;
  assign n608 = n3109 | n3146 ;
  assign n3099 = n2591 & n3075 ;
  assign n3144 = n2593 & n4396 ;
  assign n609 = n3099 | n3144 ;
  assign n2871 = n2598 & n642 ;
  assign n3274 = n2600 & n2830 ;
  assign n610 = n2871 | n3274 ;
  assign n2884 = n2606 & n642 ;
  assign n3272 = n2608 & n2830 ;
  assign n611 = n2884 | n3272 ;
  assign n2887 = n2613 & n642 ;
  assign n3270 = n2615 & n2830 ;
  assign n612 = n2887 | n3270 ;
  assign n3096 = n2622 & n3075 ;
  assign n3142 = n2624 & n4396 ;
  assign n613 = n3096 | n3142 ;
  assign n2885 = n2630 & n642 ;
  assign n3268 = n2632 & n2830 ;
  assign n614 = n2885 | n3268 ;
  assign n2886 = n2639 & n642 ;
  assign n3266 = n2641 & n2830 ;
  assign n615 = n2886 | n3266 ;
  assign n3106 = n2645 & n3075 ;
  assign n3140 = n2647 & n4396 ;
  assign n616 = n3106 | n3140 ;
  assign n2861 = n2655 & n642 ;
  assign n3264 = n2657 & n2830 ;
  assign n617 = n2861 | n3264 ;
  assign n3104 = n2662 & n3075 ;
  assign n3138 = n2664 & n4396 ;
  assign n618 = n3104 | n3138 ;
  assign n2883 = n2670 & n642 ;
  assign n3262 = n2672 & n2830 ;
  assign n619 = n2883 | n3262 ;
  assign n2878 = n2677 & n642 ;
  assign n3260 = n2679 & n2830 ;
  assign n620 = n2878 | n3260 ;
  assign n2882 = n2686 & n642 ;
  assign n3258 = n2688 & n2830 ;
  assign n621 = n2882 | n3258 ;
  assign n2877 = n2695 & n642 ;
  assign n3256 = n2697 & n2830 ;
  assign n622 = n2877 | n3256 ;
  assign n2862 = n2702 & n642 ;
  assign n3254 = n2704 & n2830 ;
  assign n623 = n2862 | n3254 ;
  assign n2855 = n2709 & n642 ;
  assign n3252 = n2711 & n2830 ;
  assign n624 = n2855 | n3252 ;
  assign n2868 = n2719 & n642 ;
  assign n3250 = n2721 & n2830 ;
  assign n625 = n2868 | n3250 ;
  assign n3103 = n2726 & n3075 ;
  assign n3136 = n2728 & n4396 ;
  assign n626 = n3103 | n3136 ;
  assign n3100 = n2735 & n3075 ;
  assign n3134 = n2737 & n4396 ;
  assign n627 = n3100 | n3134 ;
  assign n2836 = n1749 & n642 ;
  assign n3248 = n1814 & n2830 ;
  assign n628 = n2836 | n3248 ;
  assign n2857 = n1133 & n642 ;
  assign n3246 = n1678 & n2830 ;
  assign n629 = n2857 | n3246 ;
  assign n2840 = n2748 & n642 ;
  assign n3244 = n2750 & n2830 ;
  assign n630 = n2840 | n3244 ;
  assign n2874 = n2754 & n642 ;
  assign n3242 = n2756 & n2830 ;
  assign n631 = n2874 | n3242 ;
  assign n2859 = n2763 & n642 ;
  assign n3240 = n2765 & n2830 ;
  assign n632 = n2859 | n3240 ;
  assign n3111 = n2771 & n3075 ;
  assign n3132 = n2773 & n4396 ;
  assign n633 = n3111 | n3132 ;
  assign n2865 = n2779 & n642 ;
  assign n3238 = n2781 & n2830 ;
  assign n634 = n2865 | n3238 ;
  assign n3097 = n2787 & n3075 ;
  assign n3130 = n2789 & n4396 ;
  assign n635 = n3097 | n3130 ;
  assign n2867 = n2796 & n642 ;
  assign n3236 = n2798 & n2830 ;
  assign n636 = n2867 | n3236 ;
  assign n3107 = n2803 & n3075 ;
  assign n3128 = n2805 & n4396 ;
  assign n637 = n3107 | n3128 ;
  assign n2870 = n2812 & n642 ;
  assign n3234 = n2814 & n2830 ;
  assign n638 = n2870 | n3234 ;
  assign n2875 = n2818 & n642 ;
  assign n3232 = n2820 & n2830 ;
  assign n639 = n2875 | n3232 ;
  assign n640 = n3129 & n3131 ;
  assign n2876 = n1065 | n2830 ;
  assign n3230 = n3722 & n2830 ;
  assign n4417 = ~n3230 ;
  assign n3231 = n2876 & n4417 ;
  assign n641 = ~n3231 ;
  assign y0 = n513 ;
  assign y1 = n514 ;
  assign y2 = n515 ;
  assign y3 = n516 ;
  assign y4 = n517 ;
  assign y5 = n518 ;
  assign y6 = n519 ;
  assign y7 = n520 ;
  assign y8 = n521 ;
  assign y9 = n522 ;
  assign y10 = n523 ;
  assign y11 = n524 ;
  assign y12 = n525 ;
  assign y13 = n526 ;
  assign y14 = n527 ;
  assign y15 = n528 ;
  assign y16 = n529 ;
  assign y17 = n530 ;
  assign y18 = n531 ;
  assign y19 = n532 ;
  assign y20 = n533 ;
  assign y21 = n534 ;
  assign y22 = n535 ;
  assign y23 = n536 ;
  assign y24 = n537 ;
  assign y25 = n538 ;
  assign y26 = n539 ;
  assign y27 = n540 ;
  assign y28 = n541 ;
  assign y29 = n542 ;
  assign y30 = n543 ;
  assign y31 = n544 ;
  assign y32 = n545 ;
  assign y33 = n546 ;
  assign y34 = n547 ;
  assign y35 = n548 ;
  assign y36 = n549 ;
  assign y37 = n550 ;
  assign y38 = n551 ;
  assign y39 = n552 ;
  assign y40 = n553 ;
  assign y41 = n554 ;
  assign y42 = n555 ;
  assign y43 = n556 ;
  assign y44 = n557 ;
  assign y45 = n558 ;
  assign y46 = n559 ;
  assign y47 = n560 ;
  assign y48 = n561 ;
  assign y49 = n562 ;
  assign y50 = n563 ;
  assign y51 = n564 ;
  assign y52 = n565 ;
  assign y53 = n566 ;
  assign y54 = n567 ;
  assign y55 = n568 ;
  assign y56 = n569 ;
  assign y57 = n570 ;
  assign y58 = n571 ;
  assign y59 = n572 ;
  assign y60 = n573 ;
  assign y61 = n574 ;
  assign y62 = n575 ;
  assign y63 = n576 ;
  assign y64 = n577 ;
  assign y65 = n578 ;
  assign y66 = n579 ;
  assign y67 = n580 ;
  assign y68 = n581 ;
  assign y69 = n582 ;
  assign y70 = n583 ;
  assign y71 = n584 ;
  assign y72 = n585 ;
  assign y73 = n586 ;
  assign y74 = n587 ;
  assign y75 = n588 ;
  assign y76 = n589 ;
  assign y77 = n590 ;
  assign y78 = n591 ;
  assign y79 = n592 ;
  assign y80 = n593 ;
  assign y81 = n594 ;
  assign y82 = n595 ;
  assign y83 = n596 ;
  assign y84 = n597 ;
  assign y85 = n598 ;
  assign y86 = n599 ;
  assign y87 = n600 ;
  assign y88 = n601 ;
  assign y89 = n602 ;
  assign y90 = n603 ;
  assign y91 = n604 ;
  assign y92 = n605 ;
  assign y93 = n606 ;
  assign y94 = n607 ;
  assign y95 = n608 ;
  assign y96 = n609 ;
  assign y97 = n610 ;
  assign y98 = n611 ;
  assign y99 = n612 ;
  assign y100 = n613 ;
  assign y101 = n614 ;
  assign y102 = n615 ;
  assign y103 = n616 ;
  assign y104 = n617 ;
  assign y105 = n618 ;
  assign y106 = n619 ;
  assign y107 = n620 ;
  assign y108 = n621 ;
  assign y109 = n622 ;
  assign y110 = n623 ;
  assign y111 = n624 ;
  assign y112 = n625 ;
  assign y113 = n626 ;
  assign y114 = n627 ;
  assign y115 = n628 ;
  assign y116 = n629 ;
  assign y117 = n630 ;
  assign y118 = n631 ;
  assign y119 = n632 ;
  assign y120 = n633 ;
  assign y121 = n634 ;
  assign y122 = n635 ;
  assign y123 = n636 ;
  assign y124 = n637 ;
  assign y125 = n638 ;
  assign y126 = n639 ;
  assign y127 = n640 ;
  assign y128 = n641 ;
  assign y129 = n642 ;
endmodule
