module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 ;
  assign n56 = x30 | x31 ;
  assign n57 = x29 | n56 ;
  assign n58 = x28 | n57 ;
  assign n59 = x27 | n58 ;
  assign n60 = x26 | n59 ;
  assign n61 = x25 | n60 ;
  assign n62 = x24 | n61 ;
  assign n63 = x23 | n62 ;
  assign n64 = x22 | n63 ;
  assign n65 = x21 | n64 ;
  assign n66 = x20 | n65 ;
  assign n67 = x19 | n66 ;
  assign n68 = x18 | n67 ;
  assign n69 = x17 | n68 ;
  assign n1113 = ~n69 ;
  assign n72 = x16 & n1113 ;
  assign n1114 = ~x14 ;
  assign n73 = n1114 & x16 ;
  assign n74 = n68 | n73 ;
  assign n1115 = ~n74 ;
  assign n75 = x17 & n1115 ;
  assign n1116 = ~n75 ;
  assign n76 = x15 & n1116 ;
  assign n1117 = ~n72 ;
  assign n77 = n1117 & n76 ;
  assign n1118 = ~x13 ;
  assign n78 = n1118 & x16 ;
  assign n79 = x17 | n78 ;
  assign n1119 = ~x15 ;
  assign n80 = n1119 & x17 ;
  assign n81 = n74 | n80 ;
  assign n47 = ~n81 ;
  assign n82 = x16 & n47 ;
  assign n1121 = ~n82 ;
  assign n83 = x14 & n1121 ;
  assign n84 = x17 & n78 ;
  assign n1122 = ~n84 ;
  assign n85 = n83 & n1122 ;
  assign n1123 = ~n85 ;
  assign n86 = n79 & n1123 ;
  assign n87 = x18 & n86 ;
  assign n88 = n67 | n87 ;
  assign n89 = x18 | n86 ;
  assign n1124 = ~n88 ;
  assign n90 = n1124 & n89 ;
  assign n1125 = ~n90 ;
  assign n91 = n77 & n1125 ;
  assign n1126 = ~x12 ;
  assign n92 = n1126 & x16 ;
  assign n94 = x17 | n92 ;
  assign n93 = x17 & n92 ;
  assign n1127 = ~n77 ;
  assign n95 = n1127 & n89 ;
  assign n96 = n88 | n95 ;
  assign n46 = ~n96 ;
  assign n97 = x16 & n46 ;
  assign n1129 = ~n97 ;
  assign n98 = x13 & n1129 ;
  assign n99 = n78 & n46 ;
  assign n100 = n98 | n99 ;
  assign n1130 = ~n93 ;
  assign n101 = n1130 & n100 ;
  assign n1131 = ~n101 ;
  assign n102 = n94 & n1131 ;
  assign n103 = x18 | n102 ;
  assign n104 = n79 & n1122 ;
  assign n105 = n46 & n104 ;
  assign n106 = n83 & n105 ;
  assign n107 = n83 | n105 ;
  assign n1132 = ~n106 ;
  assign n108 = n1132 & n107 ;
  assign n109 = x18 & n102 ;
  assign n1133 = ~n109 ;
  assign n110 = n108 & n1133 ;
  assign n1134 = ~n110 ;
  assign n111 = n103 & n1134 ;
  assign n112 = x19 | n111 ;
  assign n113 = x19 & n111 ;
  assign n114 = n66 | n113 ;
  assign n1135 = ~n114 ;
  assign n115 = n112 & n1135 ;
  assign n1136 = ~n115 ;
  assign n116 = n91 & n1136 ;
  assign n1137 = ~x11 ;
  assign n117 = n1137 & x16 ;
  assign n119 = x17 | n117 ;
  assign n118 = x17 & n117 ;
  assign n1138 = ~n91 ;
  assign n120 = n1138 & n112 ;
  assign n121 = n114 | n120 ;
  assign n45 = ~n121 ;
  assign n122 = x16 & n45 ;
  assign n123 = x12 & n122 ;
  assign n124 = x12 | n122 ;
  assign n1140 = ~n123 ;
  assign n125 = n1140 & n124 ;
  assign n1141 = ~n118 ;
  assign n126 = n1141 & n125 ;
  assign n1142 = ~n126 ;
  assign n127 = n119 & n1142 ;
  assign n128 = x18 | n127 ;
  assign n129 = x18 & n127 ;
  assign n130 = n1130 & n94 ;
  assign n131 = n45 & n130 ;
  assign n132 = n100 & n131 ;
  assign n133 = n100 | n131 ;
  assign n1143 = ~n132 ;
  assign n134 = n1143 & n133 ;
  assign n1144 = ~n129 ;
  assign n135 = n1144 & n134 ;
  assign n1145 = ~n135 ;
  assign n136 = n128 & n1145 ;
  assign n137 = x19 | n136 ;
  assign n138 = n103 & n1133 ;
  assign n139 = n45 & n138 ;
  assign n1146 = ~n108 ;
  assign n140 = n1146 & n139 ;
  assign n1147 = ~n139 ;
  assign n141 = n108 & n1147 ;
  assign n142 = n140 | n141 ;
  assign n143 = x19 & n136 ;
  assign n1148 = ~n143 ;
  assign n144 = n142 & n1148 ;
  assign n1149 = ~n144 ;
  assign n145 = n137 & n1149 ;
  assign n146 = x20 | n145 ;
  assign n147 = x20 & n145 ;
  assign n148 = n65 | n147 ;
  assign n1150 = ~n148 ;
  assign n149 = n146 & n1150 ;
  assign n1151 = ~n149 ;
  assign n150 = n116 & n1151 ;
  assign n1152 = ~x10 ;
  assign n151 = n1152 & x16 ;
  assign n153 = x17 | n151 ;
  assign n152 = x17 & n151 ;
  assign n1153 = ~n116 ;
  assign n154 = n1153 & n146 ;
  assign n155 = n148 | n154 ;
  assign n44 = ~n155 ;
  assign n156 = x16 & n44 ;
  assign n157 = x11 & n156 ;
  assign n158 = x11 | n156 ;
  assign n1155 = ~n157 ;
  assign n159 = n1155 & n158 ;
  assign n1156 = ~n152 ;
  assign n160 = n1156 & n159 ;
  assign n1157 = ~n160 ;
  assign n161 = n153 & n1157 ;
  assign n162 = x18 | n161 ;
  assign n163 = x18 & n161 ;
  assign n164 = n1141 & n119 ;
  assign n165 = n44 & n164 ;
  assign n166 = n125 & n165 ;
  assign n167 = n125 | n165 ;
  assign n1158 = ~n166 ;
  assign n168 = n1158 & n167 ;
  assign n1159 = ~n163 ;
  assign n169 = n1159 & n168 ;
  assign n1160 = ~n169 ;
  assign n170 = n162 & n1160 ;
  assign n171 = x19 | n170 ;
  assign n172 = x19 & n170 ;
  assign n173 = n128 & n1144 ;
  assign n174 = n44 & n173 ;
  assign n1161 = ~n134 ;
  assign n175 = n1161 & n174 ;
  assign n1162 = ~n174 ;
  assign n176 = n134 & n1162 ;
  assign n177 = n175 | n176 ;
  assign n1163 = ~n172 ;
  assign n178 = n1163 & n177 ;
  assign n1164 = ~n178 ;
  assign n179 = n171 & n1164 ;
  assign n180 = x20 | n179 ;
  assign n181 = n137 & n1148 ;
  assign n182 = n44 & n181 ;
  assign n1165 = ~n142 ;
  assign n183 = n1165 & n182 ;
  assign n1166 = ~n182 ;
  assign n184 = n142 & n1166 ;
  assign n185 = n183 | n184 ;
  assign n186 = x20 & n179 ;
  assign n1167 = ~n186 ;
  assign n187 = n185 & n1167 ;
  assign n1168 = ~n187 ;
  assign n188 = n180 & n1168 ;
  assign n189 = x21 | n188 ;
  assign n190 = x21 & n188 ;
  assign n191 = n64 | n190 ;
  assign n1169 = ~n191 ;
  assign n192 = n189 & n1169 ;
  assign n1170 = ~n192 ;
  assign n193 = n150 & n1170 ;
  assign n1171 = ~x9 ;
  assign n194 = n1171 & x16 ;
  assign n196 = x17 | n194 ;
  assign n195 = x17 & n194 ;
  assign n1172 = ~n150 ;
  assign n197 = n1172 & n189 ;
  assign n198 = n191 | n197 ;
  assign n43 = ~n198 ;
  assign n199 = x16 & n43 ;
  assign n200 = x10 & n199 ;
  assign n201 = x10 | n199 ;
  assign n1174 = ~n200 ;
  assign n202 = n1174 & n201 ;
  assign n1175 = ~n195 ;
  assign n203 = n1175 & n202 ;
  assign n1176 = ~n203 ;
  assign n204 = n196 & n1176 ;
  assign n205 = x18 & n204 ;
  assign n206 = n1156 & n153 ;
  assign n207 = n43 & n206 ;
  assign n208 = n159 & n207 ;
  assign n209 = n159 | n207 ;
  assign n1177 = ~n208 ;
  assign n210 = n1177 & n209 ;
  assign n211 = x18 | n204 ;
  assign n1178 = ~n210 ;
  assign n212 = n1178 & n211 ;
  assign n213 = n205 | n212 ;
  assign n216 = x19 | n213 ;
  assign n214 = x19 & n213 ;
  assign n217 = n162 & n1159 ;
  assign n218 = n43 & n217 ;
  assign n1179 = ~n168 ;
  assign n219 = n1179 & n218 ;
  assign n1180 = ~n218 ;
  assign n220 = n168 & n1180 ;
  assign n221 = n219 | n220 ;
  assign n1181 = ~n214 ;
  assign n222 = n1181 & n221 ;
  assign n1182 = ~n222 ;
  assign n223 = n216 & n1182 ;
  assign n224 = x20 | n223 ;
  assign n225 = x20 & n223 ;
  assign n226 = n171 & n1163 ;
  assign n227 = n43 & n226 ;
  assign n1183 = ~n177 ;
  assign n228 = n1183 & n227 ;
  assign n1184 = ~n227 ;
  assign n229 = n177 & n1184 ;
  assign n230 = n228 | n229 ;
  assign n1185 = ~n225 ;
  assign n231 = n1185 & n230 ;
  assign n1186 = ~n231 ;
  assign n232 = n224 & n1186 ;
  assign n233 = x21 | n232 ;
  assign n234 = n180 & n1167 ;
  assign n235 = n43 & n234 ;
  assign n1187 = ~n185 ;
  assign n236 = n1187 & n235 ;
  assign n1188 = ~n235 ;
  assign n237 = n185 & n1188 ;
  assign n238 = n236 | n237 ;
  assign n239 = x21 & n232 ;
  assign n1189 = ~n239 ;
  assign n240 = n238 & n1189 ;
  assign n1190 = ~n240 ;
  assign n241 = n233 & n1190 ;
  assign n242 = x22 | n241 ;
  assign n243 = x22 & n241 ;
  assign n244 = n63 | n243 ;
  assign n1191 = ~n244 ;
  assign n245 = n242 & n1191 ;
  assign n1192 = ~n245 ;
  assign n246 = n193 & n1192 ;
  assign n1193 = ~x8 ;
  assign n247 = n1193 & x16 ;
  assign n249 = x17 | n247 ;
  assign n248 = x17 & n247 ;
  assign n1194 = ~n193 ;
  assign n250 = n1194 & n242 ;
  assign n251 = n244 | n250 ;
  assign n42 = ~n251 ;
  assign n252 = x16 & n42 ;
  assign n253 = x9 & n252 ;
  assign n254 = x9 | n252 ;
  assign n1196 = ~n253 ;
  assign n255 = n1196 & n254 ;
  assign n1197 = ~n248 ;
  assign n256 = n1197 & n255 ;
  assign n1198 = ~n256 ;
  assign n257 = n249 & n1198 ;
  assign n258 = x18 | n257 ;
  assign n259 = x18 & n257 ;
  assign n260 = n1175 & n196 ;
  assign n261 = n42 & n260 ;
  assign n1199 = ~n261 ;
  assign n262 = n202 & n1199 ;
  assign n1200 = ~n202 ;
  assign n263 = n1200 & n261 ;
  assign n264 = n262 | n263 ;
  assign n1201 = ~n259 ;
  assign n265 = n1201 & n264 ;
  assign n1202 = ~n265 ;
  assign n266 = n258 & n1202 ;
  assign n267 = x19 | n266 ;
  assign n1203 = ~n205 ;
  assign n268 = n1203 & n211 ;
  assign n269 = n42 & n268 ;
  assign n270 = n210 & n269 ;
  assign n271 = n210 | n269 ;
  assign n1204 = ~n270 ;
  assign n272 = n1204 & n271 ;
  assign n273 = x19 & n266 ;
  assign n1205 = ~n273 ;
  assign n274 = n272 & n1205 ;
  assign n1206 = ~n274 ;
  assign n275 = n267 & n1206 ;
  assign n276 = x20 | n275 ;
  assign n277 = x20 & n275 ;
  assign n1207 = ~x19 ;
  assign n215 = n1207 & n213 ;
  assign n1208 = ~n213 ;
  assign n278 = x19 & n1208 ;
  assign n279 = n215 | n278 ;
  assign n280 = n42 & n279 ;
  assign n1209 = ~n221 ;
  assign n281 = n1209 & n280 ;
  assign n1210 = ~n280 ;
  assign n282 = n221 & n1210 ;
  assign n283 = n281 | n282 ;
  assign n1211 = ~n277 ;
  assign n284 = n1211 & n283 ;
  assign n1212 = ~n284 ;
  assign n285 = n276 & n1212 ;
  assign n286 = x21 | n285 ;
  assign n287 = x21 & n285 ;
  assign n288 = n224 & n1185 ;
  assign n289 = n42 & n288 ;
  assign n1213 = ~n230 ;
  assign n290 = n1213 & n289 ;
  assign n1214 = ~n289 ;
  assign n291 = n230 & n1214 ;
  assign n292 = n290 | n291 ;
  assign n1215 = ~n287 ;
  assign n293 = n1215 & n292 ;
  assign n1216 = ~n293 ;
  assign n294 = n286 & n1216 ;
  assign n295 = x22 | n294 ;
  assign n296 = n233 & n1189 ;
  assign n297 = n42 & n296 ;
  assign n1217 = ~n238 ;
  assign n298 = n1217 & n297 ;
  assign n1218 = ~n297 ;
  assign n299 = n238 & n1218 ;
  assign n300 = n298 | n299 ;
  assign n301 = x22 & n294 ;
  assign n1219 = ~n301 ;
  assign n302 = n300 & n1219 ;
  assign n1220 = ~n302 ;
  assign n303 = n295 & n1220 ;
  assign n304 = x23 | n303 ;
  assign n305 = x23 & n303 ;
  assign n306 = n62 | n305 ;
  assign n1221 = ~n306 ;
  assign n307 = n304 & n1221 ;
  assign n1222 = ~n307 ;
  assign n308 = n246 & n1222 ;
  assign n1223 = ~n246 ;
  assign n309 = n1223 & n304 ;
  assign n310 = n306 | n309 ;
  assign n313 = n258 & n1201 ;
  assign n41 = ~n310 ;
  assign n314 = n41 & n313 ;
  assign n1225 = ~n264 ;
  assign n315 = n1225 & n314 ;
  assign n1226 = ~n314 ;
  assign n316 = n264 & n1226 ;
  assign n317 = n315 | n316 ;
  assign n318 = n1207 & n317 ;
  assign n1227 = ~n317 ;
  assign n319 = x19 & n1227 ;
  assign n1228 = ~x7 ;
  assign n320 = n1228 & x16 ;
  assign n322 = x17 | n320 ;
  assign n321 = x17 & n320 ;
  assign n311 = n247 & n41 ;
  assign n312 = x16 & n41 ;
  assign n1229 = ~n312 ;
  assign n323 = x8 & n1229 ;
  assign n324 = n311 | n323 ;
  assign n1230 = ~n321 ;
  assign n325 = n1230 & n324 ;
  assign n1231 = ~n325 ;
  assign n326 = n322 & n1231 ;
  assign n329 = x18 | n326 ;
  assign n327 = x18 & n326 ;
  assign n330 = n1197 & n249 ;
  assign n331 = n41 & n330 ;
  assign n332 = n255 & n331 ;
  assign n333 = n255 | n331 ;
  assign n1232 = ~n332 ;
  assign n334 = n1232 & n333 ;
  assign n1233 = ~n327 ;
  assign n335 = n1233 & n334 ;
  assign n1234 = ~n335 ;
  assign n336 = n329 & n1234 ;
  assign n337 = n319 | n336 ;
  assign n1235 = ~n318 ;
  assign n338 = n1235 & n337 ;
  assign n339 = x20 | n338 ;
  assign n341 = n267 & n1205 ;
  assign n342 = n41 & n341 ;
  assign n1236 = ~n272 ;
  assign n343 = n1236 & n342 ;
  assign n1237 = ~n342 ;
  assign n344 = n272 & n1237 ;
  assign n345 = n343 | n344 ;
  assign n346 = x20 & n338 ;
  assign n1238 = ~n346 ;
  assign n347 = n345 & n1238 ;
  assign n1239 = ~n347 ;
  assign n348 = n339 & n1239 ;
  assign n349 = x21 | n348 ;
  assign n350 = x21 & n348 ;
  assign n352 = n276 & n1211 ;
  assign n353 = n41 & n352 ;
  assign n1240 = ~n283 ;
  assign n354 = n1240 & n353 ;
  assign n1241 = ~n353 ;
  assign n355 = n283 & n1241 ;
  assign n356 = n354 | n355 ;
  assign n1242 = ~n350 ;
  assign n357 = n1242 & n356 ;
  assign n1243 = ~n357 ;
  assign n358 = n349 & n1243 ;
  assign n359 = x22 | n358 ;
  assign n360 = x22 & n358 ;
  assign n362 = n286 & n1215 ;
  assign n363 = n41 & n362 ;
  assign n1244 = ~n292 ;
  assign n364 = n1244 & n363 ;
  assign n1245 = ~n363 ;
  assign n365 = n292 & n1245 ;
  assign n366 = n364 | n365 ;
  assign n1246 = ~n360 ;
  assign n367 = n1246 & n366 ;
  assign n1247 = ~n367 ;
  assign n368 = n359 & n1247 ;
  assign n369 = x23 | n368 ;
  assign n370 = n295 & n1219 ;
  assign n371 = n41 & n370 ;
  assign n1248 = ~n300 ;
  assign n372 = n1248 & n371 ;
  assign n1249 = ~n371 ;
  assign n373 = n300 & n1249 ;
  assign n374 = n372 | n373 ;
  assign n375 = x23 & n368 ;
  assign n1250 = ~n375 ;
  assign n377 = n374 & n1250 ;
  assign n1251 = ~n377 ;
  assign n378 = n369 & n1251 ;
  assign n379 = x24 | n378 ;
  assign n380 = x24 & n378 ;
  assign n381 = n61 | n380 ;
  assign n1252 = ~n381 ;
  assign n382 = n379 & n1252 ;
  assign n1253 = ~n382 ;
  assign n383 = n308 & n1253 ;
  assign n1254 = ~x6 ;
  assign n384 = n1254 & x16 ;
  assign n386 = x17 | n384 ;
  assign n385 = x17 & n384 ;
  assign n1255 = ~n308 ;
  assign n388 = n1255 & n379 ;
  assign n389 = n381 | n388 ;
  assign n40 = ~n389 ;
  assign n403 = x16 & n40 ;
  assign n404 = x7 & n403 ;
  assign n405 = x7 | n403 ;
  assign n1257 = ~n404 ;
  assign n406 = n1257 & n405 ;
  assign n1258 = ~n385 ;
  assign n407 = n1258 & n406 ;
  assign n1259 = ~n407 ;
  assign n408 = n386 & n1259 ;
  assign n409 = x18 & n408 ;
  assign n410 = n1230 & n322 ;
  assign n411 = n40 & n410 ;
  assign n412 = n324 & n411 ;
  assign n413 = n324 | n411 ;
  assign n1260 = ~n412 ;
  assign n414 = n1260 & n413 ;
  assign n415 = x18 | n408 ;
  assign n1261 = ~n414 ;
  assign n417 = n1261 & n415 ;
  assign n418 = n409 | n417 ;
  assign n423 = x19 | n418 ;
  assign n420 = x19 & n418 ;
  assign n1262 = ~x18 ;
  assign n328 = n1262 & n326 ;
  assign n1263 = ~n326 ;
  assign n424 = x18 & n1263 ;
  assign n425 = n328 | n424 ;
  assign n426 = n40 & n425 ;
  assign n1264 = ~n334 ;
  assign n427 = n1264 & n426 ;
  assign n1265 = ~n426 ;
  assign n428 = n334 & n1265 ;
  assign n429 = n427 | n428 ;
  assign n1266 = ~n420 ;
  assign n430 = n1266 & n429 ;
  assign n1267 = ~n430 ;
  assign n431 = n423 & n1267 ;
  assign n432 = x20 | n431 ;
  assign n433 = x20 & n431 ;
  assign n435 = n318 | n319 ;
  assign n402 = n336 & n40 ;
  assign n436 = x19 & n389 ;
  assign n437 = n402 | n436 ;
  assign n1268 = ~n435 ;
  assign n438 = n1268 & n437 ;
  assign n1269 = ~n437 ;
  assign n439 = n435 & n1269 ;
  assign n440 = n438 | n439 ;
  assign n1270 = ~n433 ;
  assign n441 = n1270 & n440 ;
  assign n1271 = ~n441 ;
  assign n442 = n432 & n1271 ;
  assign n443 = x21 | n442 ;
  assign n444 = x21 & n442 ;
  assign n1272 = ~n338 ;
  assign n340 = x20 & n1272 ;
  assign n1273 = ~x20 ;
  assign n446 = n1273 & n338 ;
  assign n447 = n340 | n446 ;
  assign n448 = n40 & n447 ;
  assign n449 = n345 & n448 ;
  assign n450 = n345 | n448 ;
  assign n1274 = ~n449 ;
  assign n451 = n1274 & n450 ;
  assign n1275 = ~n444 ;
  assign n452 = n1275 & n451 ;
  assign n1276 = ~n452 ;
  assign n453 = n443 & n1276 ;
  assign n454 = x22 | n453 ;
  assign n351 = n349 & n1242 ;
  assign n390 = n351 & n40 ;
  assign n1277 = ~n356 ;
  assign n391 = n1277 & n390 ;
  assign n1278 = ~n390 ;
  assign n392 = n356 & n1278 ;
  assign n393 = n391 | n392 ;
  assign n455 = x22 & n453 ;
  assign n1279 = ~n455 ;
  assign n456 = n393 & n1279 ;
  assign n1280 = ~n456 ;
  assign n457 = n454 & n1280 ;
  assign n458 = x23 | n457 ;
  assign n361 = n359 & n1246 ;
  assign n394 = n361 & n40 ;
  assign n1281 = ~n366 ;
  assign n395 = n1281 & n394 ;
  assign n1282 = ~n394 ;
  assign n396 = n366 & n1282 ;
  assign n397 = n395 | n396 ;
  assign n459 = x23 & n457 ;
  assign n1283 = ~n459 ;
  assign n460 = n397 & n1283 ;
  assign n1284 = ~n460 ;
  assign n461 = n458 & n1284 ;
  assign n462 = x24 | n461 ;
  assign n376 = n369 & n1250 ;
  assign n398 = n376 & n40 ;
  assign n1285 = ~n374 ;
  assign n399 = n1285 & n398 ;
  assign n1286 = ~n398 ;
  assign n400 = n374 & n1286 ;
  assign n401 = n399 | n400 ;
  assign n463 = x24 & n461 ;
  assign n1287 = ~n463 ;
  assign n464 = n401 & n1287 ;
  assign n1288 = ~n464 ;
  assign n465 = n462 & n1288 ;
  assign n466 = x25 | n465 ;
  assign n468 = x25 & n465 ;
  assign n469 = n60 | n468 ;
  assign n1289 = ~n469 ;
  assign n470 = n466 & n1289 ;
  assign n1290 = ~n470 ;
  assign n471 = n383 & n1290 ;
  assign n1291 = ~n409 ;
  assign n416 = n1291 & n415 ;
  assign n1292 = ~n383 ;
  assign n467 = n1292 & n466 ;
  assign n472 = n467 | n469 ;
  assign n39 = ~n472 ;
  assign n473 = n416 & n39 ;
  assign n474 = n414 & n473 ;
  assign n475 = n414 | n473 ;
  assign n1294 = ~n474 ;
  assign n476 = n1294 & n475 ;
  assign n477 = n1207 & n476 ;
  assign n1295 = ~n476 ;
  assign n478 = x19 & n1295 ;
  assign n1296 = ~x5 ;
  assign n1120 = n1296 & x16 ;
  assign n1139 = x17 | n1120 ;
  assign n1128 = x17 & n1120 ;
  assign n480 = x16 & n39 ;
  assign n481 = x6 & n480 ;
  assign n482 = x6 | n480 ;
  assign n1297 = ~n481 ;
  assign n483 = n1297 & n482 ;
  assign n1298 = ~n1128 ;
  assign n484 = n1298 & n483 ;
  assign n1299 = ~n484 ;
  assign n485 = n1139 & n1299 ;
  assign n487 = x18 | n485 ;
  assign n486 = x18 & n485 ;
  assign n387 = n1258 & n386 ;
  assign n493 = n387 & n39 ;
  assign n494 = n406 & n493 ;
  assign n495 = n406 | n493 ;
  assign n1300 = ~n494 ;
  assign n496 = n1300 & n495 ;
  assign n1301 = ~n486 ;
  assign n497 = n1301 & n496 ;
  assign n1302 = ~n497 ;
  assign n498 = n487 & n1302 ;
  assign n499 = n478 | n498 ;
  assign n1303 = ~n477 ;
  assign n500 = n1303 & n499 ;
  assign n501 = x20 | n500 ;
  assign n419 = n1207 & n418 ;
  assign n1304 = ~n418 ;
  assign n421 = x19 & n1304 ;
  assign n422 = n419 | n421 ;
  assign n489 = n422 & n39 ;
  assign n1305 = ~n429 ;
  assign n490 = n1305 & n489 ;
  assign n1306 = ~n489 ;
  assign n491 = n429 & n1306 ;
  assign n492 = n490 | n491 ;
  assign n502 = x20 & n500 ;
  assign n1307 = ~n502 ;
  assign n503 = n492 & n1307 ;
  assign n1308 = ~n503 ;
  assign n504 = n501 & n1308 ;
  assign n505 = x21 | n504 ;
  assign n506 = x21 & n504 ;
  assign n434 = n432 & n1270 ;
  assign n509 = n434 & n39 ;
  assign n510 = n440 & n509 ;
  assign n511 = n440 | n509 ;
  assign n1309 = ~n510 ;
  assign n512 = n1309 & n511 ;
  assign n1310 = ~n506 ;
  assign n513 = n1310 & n512 ;
  assign n1311 = ~n513 ;
  assign n514 = n505 & n1311 ;
  assign n515 = x22 | n514 ;
  assign n516 = x22 & n514 ;
  assign n445 = n443 & n1275 ;
  assign n518 = n445 & n39 ;
  assign n1312 = ~n451 ;
  assign n519 = n1312 & n518 ;
  assign n1313 = ~n518 ;
  assign n520 = n451 & n1313 ;
  assign n521 = n519 | n520 ;
  assign n1314 = ~n516 ;
  assign n522 = n1314 & n521 ;
  assign n1315 = ~n522 ;
  assign n523 = n515 & n1315 ;
  assign n524 = x23 | n523 ;
  assign n525 = x23 & n523 ;
  assign n537 = n454 & n1279 ;
  assign n538 = n39 & n537 ;
  assign n1316 = ~n393 ;
  assign n539 = n1316 & n538 ;
  assign n1317 = ~n538 ;
  assign n540 = n393 & n1317 ;
  assign n541 = n539 | n540 ;
  assign n1318 = ~n525 ;
  assign n542 = n1318 & n541 ;
  assign n1319 = ~n542 ;
  assign n543 = n524 & n1319 ;
  assign n544 = x24 | n543 ;
  assign n532 = n458 & n1283 ;
  assign n533 = n39 & n532 ;
  assign n1320 = ~n397 ;
  assign n534 = n1320 & n533 ;
  assign n1321 = ~n533 ;
  assign n535 = n397 & n1321 ;
  assign n536 = n534 | n535 ;
  assign n545 = x24 & n543 ;
  assign n1322 = ~n545 ;
  assign n546 = n536 & n1322 ;
  assign n1323 = ~n546 ;
  assign n547 = n544 & n1323 ;
  assign n548 = x25 | n547 ;
  assign n527 = n462 & n1287 ;
  assign n528 = n39 & n527 ;
  assign n1324 = ~n401 ;
  assign n529 = n1324 & n528 ;
  assign n1325 = ~n528 ;
  assign n530 = n401 & n1325 ;
  assign n531 = n529 | n530 ;
  assign n549 = x25 & n547 ;
  assign n1326 = ~n549 ;
  assign n550 = n531 & n1326 ;
  assign n1327 = ~n550 ;
  assign n551 = n548 & n1327 ;
  assign n552 = x26 | n551 ;
  assign n554 = x26 & n551 ;
  assign n555 = n59 | n554 ;
  assign n1328 = ~n555 ;
  assign n556 = n552 & n1328 ;
  assign n1329 = ~n556 ;
  assign n557 = n471 & n1329 ;
  assign n488 = n1301 & n487 ;
  assign n1330 = ~n471 ;
  assign n553 = n1330 & n552 ;
  assign n558 = n553 | n555 ;
  assign n38 = ~n558 ;
  assign n559 = n488 & n38 ;
  assign n1332 = ~n559 ;
  assign n560 = n496 & n1332 ;
  assign n1333 = ~n496 ;
  assign n561 = n1333 & n559 ;
  assign n562 = n560 | n561 ;
  assign n564 = n1207 & n562 ;
  assign n1334 = ~n562 ;
  assign n563 = x19 & n1334 ;
  assign n1335 = ~x4 ;
  assign n1154 = n1335 & x16 ;
  assign n1195 = x17 | n1154 ;
  assign n1173 = x17 & n1154 ;
  assign n566 = x16 & n38 ;
  assign n567 = x5 & n566 ;
  assign n568 = x5 | n566 ;
  assign n1336 = ~n567 ;
  assign n569 = n1336 & n568 ;
  assign n1337 = ~n1173 ;
  assign n570 = n1337 & n569 ;
  assign n1338 = ~n570 ;
  assign n571 = n1195 & n1338 ;
  assign n573 = x18 | n571 ;
  assign n572 = x18 & n571 ;
  assign n1224 = n1298 & n1139 ;
  assign n576 = n1224 & n38 ;
  assign n577 = n483 & n576 ;
  assign n578 = n483 | n576 ;
  assign n1339 = ~n577 ;
  assign n579 = n1339 & n578 ;
  assign n1340 = ~n572 ;
  assign n580 = n1340 & n579 ;
  assign n1341 = ~n580 ;
  assign n581 = n573 & n1341 ;
  assign n582 = n563 | n581 ;
  assign n1342 = ~n564 ;
  assign n583 = n1342 & n582 ;
  assign n584 = x20 | n583 ;
  assign n585 = x20 & n583 ;
  assign n479 = n477 | n478 ;
  assign n575 = x19 & n558 ;
  assign n591 = n498 & n38 ;
  assign n592 = n575 | n591 ;
  assign n1343 = ~n479 ;
  assign n593 = n1343 & n592 ;
  assign n1344 = ~n592 ;
  assign n594 = n479 & n1344 ;
  assign n595 = n593 | n594 ;
  assign n1345 = ~n585 ;
  assign n596 = n1345 & n595 ;
  assign n1346 = ~n596 ;
  assign n597 = n584 & n1346 ;
  assign n598 = x21 | n597 ;
  assign n599 = x21 & n597 ;
  assign n508 = n501 & n1307 ;
  assign n601 = n508 & n38 ;
  assign n1347 = ~n492 ;
  assign n602 = n1347 & n601 ;
  assign n1348 = ~n601 ;
  assign n603 = n492 & n1348 ;
  assign n604 = n602 | n603 ;
  assign n1349 = ~n599 ;
  assign n605 = n1349 & n604 ;
  assign n1350 = ~n605 ;
  assign n606 = n598 & n1350 ;
  assign n607 = x22 | n606 ;
  assign n507 = n505 & n1310 ;
  assign n587 = n507 & n38 ;
  assign n588 = n512 & n587 ;
  assign n589 = n512 | n587 ;
  assign n1351 = ~n588 ;
  assign n590 = n1351 & n589 ;
  assign n608 = x22 & n606 ;
  assign n1352 = ~n608 ;
  assign n609 = n590 & n1352 ;
  assign n1353 = ~n609 ;
  assign n610 = n607 & n1353 ;
  assign n611 = x23 | n610 ;
  assign n612 = x23 & n610 ;
  assign n517 = n515 & n1314 ;
  assign n615 = n517 & n38 ;
  assign n1354 = ~n521 ;
  assign n616 = n1354 & n615 ;
  assign n1355 = ~n615 ;
  assign n617 = n521 & n1355 ;
  assign n618 = n616 | n617 ;
  assign n1356 = ~n612 ;
  assign n619 = n1356 & n618 ;
  assign n1357 = ~n619 ;
  assign n620 = n611 & n1357 ;
  assign n621 = x24 | n620 ;
  assign n622 = x24 & n620 ;
  assign n526 = n524 & n1318 ;
  assign n624 = n526 & n38 ;
  assign n1358 = ~n541 ;
  assign n625 = n1358 & n624 ;
  assign n1359 = ~n624 ;
  assign n636 = n541 & n1359 ;
  assign n637 = n625 | n636 ;
  assign n1360 = ~n622 ;
  assign n638 = n1360 & n637 ;
  assign n1361 = ~n638 ;
  assign n639 = n621 & n1361 ;
  assign n640 = x25 | n639 ;
  assign n631 = n544 & n1322 ;
  assign n632 = n38 & n631 ;
  assign n1362 = ~n536 ;
  assign n633 = n1362 & n632 ;
  assign n1363 = ~n632 ;
  assign n634 = n536 & n1363 ;
  assign n635 = n633 | n634 ;
  assign n641 = x25 & n639 ;
  assign n1364 = ~n641 ;
  assign n642 = n635 & n1364 ;
  assign n1365 = ~n642 ;
  assign n643 = n640 & n1365 ;
  assign n644 = x26 | n643 ;
  assign n626 = n548 & n1326 ;
  assign n627 = n38 & n626 ;
  assign n1366 = ~n531 ;
  assign n628 = n1366 & n627 ;
  assign n1367 = ~n627 ;
  assign n629 = n531 & n1367 ;
  assign n630 = n628 | n629 ;
  assign n645 = x26 & n643 ;
  assign n1368 = ~n645 ;
  assign n646 = n630 & n1368 ;
  assign n1369 = ~n646 ;
  assign n647 = n644 & n1369 ;
  assign n648 = x27 | n647 ;
  assign n650 = x27 & n647 ;
  assign n651 = n58 | n650 ;
  assign n1370 = ~n651 ;
  assign n652 = n648 & n1370 ;
  assign n1371 = ~n652 ;
  assign n653 = n557 & n1371 ;
  assign n574 = n1340 & n573 ;
  assign n1372 = ~n557 ;
  assign n649 = n1372 & n648 ;
  assign n654 = n649 | n651 ;
  assign n37 = ~n654 ;
  assign n664 = n574 & n37 ;
  assign n1374 = ~n664 ;
  assign n665 = n579 & n1374 ;
  assign n1375 = ~n579 ;
  assign n666 = n1375 & n664 ;
  assign n667 = n665 | n666 ;
  assign n1376 = ~x3 ;
  assign n1256 = n1376 & x16 ;
  assign n1331 = x17 | n1256 ;
  assign n1293 = x17 & n1256 ;
  assign n655 = x16 & n37 ;
  assign n656 = x4 & n655 ;
  assign n657 = x4 | n655 ;
  assign n1377 = ~n656 ;
  assign n658 = n1377 & n657 ;
  assign n1378 = ~n1293 ;
  assign n659 = n1378 & n658 ;
  assign n1379 = ~n659 ;
  assign n660 = n1331 & n1379 ;
  assign n661 = x18 & n660 ;
  assign n662 = x18 | n660 ;
  assign n1373 = n1337 & n1195 ;
  assign n668 = n1373 & n37 ;
  assign n669 = n569 & n668 ;
  assign n670 = n569 | n668 ;
  assign n1380 = ~n669 ;
  assign n671 = n1380 & n670 ;
  assign n1381 = ~n671 ;
  assign n672 = n662 & n1381 ;
  assign n673 = n661 | n672 ;
  assign n674 = x19 & n673 ;
  assign n1382 = ~n674 ;
  assign n675 = n667 & n1382 ;
  assign n677 = x19 | n673 ;
  assign n1383 = ~n675 ;
  assign n678 = n1383 & n677 ;
  assign n679 = x20 | n678 ;
  assign n680 = x20 & n678 ;
  assign n565 = n563 | n564 ;
  assign n692 = n581 & n37 ;
  assign n701 = x19 & n654 ;
  assign n702 = n692 | n701 ;
  assign n1384 = ~n565 ;
  assign n703 = n1384 & n702 ;
  assign n1385 = ~n702 ;
  assign n704 = n565 & n1385 ;
  assign n705 = n703 | n704 ;
  assign n1386 = ~n680 ;
  assign n706 = n1386 & n705 ;
  assign n1387 = ~n706 ;
  assign n707 = n679 & n1387 ;
  assign n708 = x21 | n707 ;
  assign n586 = n584 & n1345 ;
  assign n693 = n586 & n37 ;
  assign n694 = n595 & n693 ;
  assign n695 = n595 | n693 ;
  assign n1388 = ~n694 ;
  assign n696 = n1388 & n695 ;
  assign n709 = x21 & n707 ;
  assign n1389 = ~n709 ;
  assign n710 = n696 & n1389 ;
  assign n1390 = ~n710 ;
  assign n711 = n708 & n1390 ;
  assign n712 = x22 | n711 ;
  assign n600 = n598 & n1349 ;
  assign n697 = n600 & n37 ;
  assign n1391 = ~n604 ;
  assign n698 = n1391 & n697 ;
  assign n1392 = ~n697 ;
  assign n699 = n604 & n1392 ;
  assign n700 = n698 | n699 ;
  assign n713 = x22 & n711 ;
  assign n1393 = ~n713 ;
  assign n714 = n700 & n1393 ;
  assign n1394 = ~n714 ;
  assign n715 = n712 & n1394 ;
  assign n716 = x23 | n715 ;
  assign n614 = n607 & n1352 ;
  assign n684 = n614 & n37 ;
  assign n1395 = ~n590 ;
  assign n685 = n1395 & n684 ;
  assign n1396 = ~n684 ;
  assign n686 = n590 & n1396 ;
  assign n687 = n685 | n686 ;
  assign n717 = x23 & n715 ;
  assign n1397 = ~n717 ;
  assign n718 = n687 & n1397 ;
  assign n1398 = ~n718 ;
  assign n719 = n716 & n1398 ;
  assign n720 = x24 | n719 ;
  assign n613 = n611 & n1356 ;
  assign n688 = n613 & n37 ;
  assign n1399 = ~n618 ;
  assign n689 = n1399 & n688 ;
  assign n1400 = ~n688 ;
  assign n690 = n618 & n1400 ;
  assign n691 = n689 | n690 ;
  assign n721 = x24 & n719 ;
  assign n1401 = ~n721 ;
  assign n722 = n691 & n1401 ;
  assign n1402 = ~n722 ;
  assign n723 = n720 & n1402 ;
  assign n724 = x25 | n723 ;
  assign n725 = x25 & n723 ;
  assign n623 = n621 & n1360 ;
  assign n731 = n623 & n37 ;
  assign n1403 = ~n637 ;
  assign n732 = n1403 & n731 ;
  assign n1404 = ~n731 ;
  assign n743 = n637 & n1404 ;
  assign n744 = n732 | n743 ;
  assign n1405 = ~n725 ;
  assign n745 = n1405 & n744 ;
  assign n1406 = ~n745 ;
  assign n746 = n724 & n1406 ;
  assign n747 = x26 | n746 ;
  assign n738 = n640 & n1364 ;
  assign n739 = n37 & n738 ;
  assign n1407 = ~n635 ;
  assign n740 = n1407 & n739 ;
  assign n1408 = ~n739 ;
  assign n741 = n635 & n1408 ;
  assign n742 = n740 | n741 ;
  assign n748 = x26 & n746 ;
  assign n1409 = ~n748 ;
  assign n749 = n742 & n1409 ;
  assign n1410 = ~n749 ;
  assign n750 = n747 & n1410 ;
  assign n751 = x27 | n750 ;
  assign n733 = n644 & n1368 ;
  assign n734 = n37 & n733 ;
  assign n1411 = ~n630 ;
  assign n735 = n1411 & n734 ;
  assign n1412 = ~n734 ;
  assign n736 = n630 & n1412 ;
  assign n737 = n735 | n736 ;
  assign n752 = x27 & n750 ;
  assign n1413 = ~n752 ;
  assign n753 = n737 & n1413 ;
  assign n1414 = ~n753 ;
  assign n754 = n751 & n1414 ;
  assign n755 = x28 | n754 ;
  assign n757 = x28 & n754 ;
  assign n758 = n57 | n757 ;
  assign n1415 = ~n758 ;
  assign n759 = n755 & n1415 ;
  assign n1416 = ~n759 ;
  assign n760 = n653 & n1416 ;
  assign n1417 = ~x2 ;
  assign n1419 = n1417 & x16 ;
  assign n1523 = x17 | n1419 ;
  assign n1469 = x17 & n1419 ;
  assign n1418 = ~n653 ;
  assign n756 = n1418 & n755 ;
  assign n761 = n756 | n758 ;
  assign n36 = ~n761 ;
  assign n762 = x16 & n36 ;
  assign n763 = x3 & n762 ;
  assign n764 = x3 | n762 ;
  assign n1420 = ~n763 ;
  assign n765 = n1420 & n764 ;
  assign n1421 = ~n1469 ;
  assign n766 = n1421 & n765 ;
  assign n1422 = ~n766 ;
  assign n767 = n1523 & n1422 ;
  assign n769 = x18 | n767 ;
  assign n768 = x18 & n767 ;
  assign n1582 = n1378 & n1331 ;
  assign n775 = n1582 & n36 ;
  assign n776 = n658 & n775 ;
  assign n777 = n658 | n775 ;
  assign n1423 = ~n776 ;
  assign n778 = n1423 & n777 ;
  assign n1424 = ~n768 ;
  assign n779 = n1424 & n778 ;
  assign n1425 = ~n779 ;
  assign n780 = n769 & n1425 ;
  assign n781 = x19 | n780 ;
  assign n1426 = ~n661 ;
  assign n663 = n1426 & n662 ;
  assign n771 = n663 & n36 ;
  assign n1427 = ~n771 ;
  assign n772 = n671 & n1427 ;
  assign n773 = n1381 & n771 ;
  assign n774 = n772 | n773 ;
  assign n782 = x19 & n780 ;
  assign n1428 = ~n782 ;
  assign n783 = n774 & n1428 ;
  assign n1429 = ~n783 ;
  assign n784 = n781 & n1429 ;
  assign n785 = x20 | n784 ;
  assign n786 = x20 & n784 ;
  assign n676 = n1207 & n673 ;
  assign n1430 = ~n673 ;
  assign n682 = x19 & n1430 ;
  assign n683 = n676 | n682 ;
  assign n789 = n683 & n36 ;
  assign n1431 = ~n667 ;
  assign n790 = n1431 & n789 ;
  assign n1432 = ~n789 ;
  assign n791 = n667 & n1432 ;
  assign n792 = n790 | n791 ;
  assign n1433 = ~n786 ;
  assign n793 = n1433 & n792 ;
  assign n1434 = ~n793 ;
  assign n794 = n785 & n1434 ;
  assign n795 = x21 | n794 ;
  assign n796 = x21 & n794 ;
  assign n681 = n679 & n1386 ;
  assign n798 = n681 & n36 ;
  assign n799 = n705 & n798 ;
  assign n800 = n705 | n798 ;
  assign n1435 = ~n799 ;
  assign n801 = n1435 & n800 ;
  assign n1436 = ~n796 ;
  assign n802 = n1436 & n801 ;
  assign n1437 = ~n802 ;
  assign n803 = n795 & n1437 ;
  assign n804 = x22 | n803 ;
  assign n805 = x22 & n803 ;
  assign n730 = n708 & n1389 ;
  assign n811 = n730 & n36 ;
  assign n812 = n696 & n811 ;
  assign n813 = n696 | n811 ;
  assign n1438 = ~n812 ;
  assign n814 = n1438 & n813 ;
  assign n1439 = ~n805 ;
  assign n815 = n1439 & n814 ;
  assign n1440 = ~n815 ;
  assign n816 = n804 & n1440 ;
  assign n817 = x23 | n816 ;
  assign n729 = n712 & n1393 ;
  assign n807 = n729 & n36 ;
  assign n1441 = ~n700 ;
  assign n808 = n1441 & n807 ;
  assign n1442 = ~n807 ;
  assign n809 = n700 & n1442 ;
  assign n810 = n808 | n809 ;
  assign n818 = x23 & n816 ;
  assign n1443 = ~n818 ;
  assign n819 = n810 & n1443 ;
  assign n1444 = ~n819 ;
  assign n820 = n817 & n1444 ;
  assign n821 = x24 | n820 ;
  assign n822 = x24 & n820 ;
  assign n728 = n716 & n1397 ;
  assign n829 = n728 & n36 ;
  assign n1445 = ~n687 ;
  assign n830 = n1445 & n829 ;
  assign n1446 = ~n829 ;
  assign n831 = n687 & n1446 ;
  assign n832 = n830 | n831 ;
  assign n1447 = ~n822 ;
  assign n833 = n1447 & n832 ;
  assign n1448 = ~n833 ;
  assign n834 = n821 & n1448 ;
  assign n835 = x25 | n834 ;
  assign n727 = n720 & n1401 ;
  assign n825 = n727 & n36 ;
  assign n1449 = ~n691 ;
  assign n826 = n1449 & n825 ;
  assign n1450 = ~n825 ;
  assign n827 = n691 & n1450 ;
  assign n828 = n826 | n827 ;
  assign n836 = x25 & n834 ;
  assign n1451 = ~n836 ;
  assign n837 = n828 & n1451 ;
  assign n1452 = ~n837 ;
  assign n838 = n835 & n1452 ;
  assign n839 = x26 | n838 ;
  assign n840 = x26 & n838 ;
  assign n726 = n724 & n1405 ;
  assign n843 = n726 & n36 ;
  assign n1453 = ~n744 ;
  assign n844 = n1453 & n843 ;
  assign n1454 = ~n843 ;
  assign n845 = n744 & n1454 ;
  assign n846 = n844 | n845 ;
  assign n1455 = ~n840 ;
  assign n847 = n1455 & n846 ;
  assign n1456 = ~n847 ;
  assign n848 = n839 & n1456 ;
  assign n849 = x27 | n848 ;
  assign n850 = x27 & n848 ;
  assign n857 = n747 & n1409 ;
  assign n858 = n36 & n857 ;
  assign n1457 = ~n742 ;
  assign n859 = n1457 & n858 ;
  assign n1458 = ~n858 ;
  assign n860 = n742 & n1458 ;
  assign n861 = n859 | n860 ;
  assign n1459 = ~n850 ;
  assign n862 = n1459 & n861 ;
  assign n1460 = ~n862 ;
  assign n863 = n849 & n1460 ;
  assign n864 = x28 | n863 ;
  assign n852 = n751 & n1413 ;
  assign n853 = n36 & n852 ;
  assign n1461 = ~n737 ;
  assign n854 = n1461 & n853 ;
  assign n1462 = ~n853 ;
  assign n855 = n737 & n1462 ;
  assign n856 = n854 | n855 ;
  assign n865 = x28 & n863 ;
  assign n1463 = ~n865 ;
  assign n866 = n856 & n1463 ;
  assign n1464 = ~n866 ;
  assign n867 = n864 & n1464 ;
  assign n868 = x29 | n867 ;
  assign n870 = x29 & n867 ;
  assign n871 = n56 | n870 ;
  assign n1465 = ~n871 ;
  assign n872 = n868 & n1465 ;
  assign n1466 = ~n872 ;
  assign n873 = n760 & n1466 ;
  assign n1467 = ~x31 ;
  assign n875 = n1467 & n873 ;
  assign n788 = n781 & n1428 ;
  assign n1468 = ~n760 ;
  assign n869 = n1468 & n868 ;
  assign n876 = n869 | n871 ;
  assign n35 = ~n876 ;
  assign n877 = n788 & n35 ;
  assign n1470 = ~n774 ;
  assign n878 = n1470 & n877 ;
  assign n1471 = ~n877 ;
  assign n879 = n774 & n1471 ;
  assign n880 = n878 | n879 ;
  assign n882 = n1273 & n880 ;
  assign n1472 = ~n880 ;
  assign n881 = x20 & n1472 ;
  assign n1473 = ~x1 ;
  assign n1583 = n1473 & x16 ;
  assign n50 = x17 | n1583 ;
  assign n49 = x17 & n1583 ;
  assign n884 = x16 & n35 ;
  assign n885 = x2 & n884 ;
  assign n886 = x2 | n884 ;
  assign n1474 = ~n885 ;
  assign n887 = n1474 & n886 ;
  assign n1475 = ~n49 ;
  assign n888 = n1475 & n887 ;
  assign n1476 = ~n888 ;
  assign n889 = n50 & n1476 ;
  assign n891 = x18 | n889 ;
  assign n890 = x18 & n889 ;
  assign n51 = n1421 & n1523 ;
  assign n897 = n51 & n35 ;
  assign n898 = n765 & n897 ;
  assign n899 = n765 | n897 ;
  assign n1477 = ~n898 ;
  assign n900 = n1477 & n899 ;
  assign n1478 = ~n890 ;
  assign n901 = n1478 & n900 ;
  assign n1479 = ~n901 ;
  assign n902 = n891 & n1479 ;
  assign n903 = x19 | n902 ;
  assign n904 = x19 & n902 ;
  assign n770 = n1424 & n769 ;
  assign n906 = n770 & n35 ;
  assign n1480 = ~n778 ;
  assign n907 = n1480 & n906 ;
  assign n1481 = ~n906 ;
  assign n908 = n778 & n1481 ;
  assign n909 = n907 | n908 ;
  assign n1482 = ~n904 ;
  assign n910 = n1482 & n909 ;
  assign n1483 = ~n910 ;
  assign n911 = n903 & n1483 ;
  assign n912 = n881 | n911 ;
  assign n1484 = ~n882 ;
  assign n913 = n1484 & n912 ;
  assign n914 = x21 | n913 ;
  assign n915 = x21 & n913 ;
  assign n787 = n785 & n1433 ;
  assign n919 = n787 & n35 ;
  assign n1485 = ~n792 ;
  assign n920 = n1485 & n919 ;
  assign n1486 = ~n919 ;
  assign n921 = n792 & n1486 ;
  assign n922 = n920 | n921 ;
  assign n1487 = ~n915 ;
  assign n923 = n1487 & n922 ;
  assign n1488 = ~n923 ;
  assign n924 = n914 & n1488 ;
  assign n925 = x22 | n924 ;
  assign n926 = x22 & n924 ;
  assign n797 = n795 & n1436 ;
  assign n928 = n797 & n35 ;
  assign n929 = n801 & n928 ;
  assign n930 = n801 | n928 ;
  assign n1489 = ~n929 ;
  assign n931 = n1489 & n930 ;
  assign n1490 = ~n926 ;
  assign n932 = n1490 & n931 ;
  assign n1491 = ~n932 ;
  assign n933 = n925 & n1491 ;
  assign n934 = x23 | n933 ;
  assign n935 = x23 & n933 ;
  assign n806 = n804 & n1439 ;
  assign n937 = n806 & n35 ;
  assign n1492 = ~n814 ;
  assign n938 = n1492 & n937 ;
  assign n1493 = ~n937 ;
  assign n939 = n814 & n1493 ;
  assign n940 = n938 | n939 ;
  assign n1494 = ~n935 ;
  assign n941 = n1494 & n940 ;
  assign n1495 = ~n941 ;
  assign n942 = n934 & n1495 ;
  assign n943 = x24 | n942 ;
  assign n944 = x24 & n942 ;
  assign n824 = n817 & n1443 ;
  assign n950 = n824 & n35 ;
  assign n1496 = ~n810 ;
  assign n951 = n1496 & n950 ;
  assign n1497 = ~n950 ;
  assign n952 = n810 & n1497 ;
  assign n953 = n951 | n952 ;
  assign n1498 = ~n944 ;
  assign n954 = n1498 & n953 ;
  assign n1499 = ~n954 ;
  assign n955 = n943 & n1499 ;
  assign n956 = x25 | n955 ;
  assign n957 = x25 & n955 ;
  assign n823 = n821 & n1447 ;
  assign n959 = n823 & n35 ;
  assign n1500 = ~n832 ;
  assign n960 = n1500 & n959 ;
  assign n1501 = ~n959 ;
  assign n961 = n832 & n1501 ;
  assign n962 = n960 | n961 ;
  assign n1502 = ~n957 ;
  assign n963 = n1502 & n962 ;
  assign n1503 = ~n963 ;
  assign n964 = n956 & n1503 ;
  assign n965 = x26 | n964 ;
  assign n842 = n835 & n1451 ;
  assign n893 = n842 & n35 ;
  assign n1504 = ~n828 ;
  assign n894 = n1504 & n893 ;
  assign n1505 = ~n893 ;
  assign n895 = n828 & n1505 ;
  assign n896 = n894 | n895 ;
  assign n966 = x26 & n964 ;
  assign n1506 = ~n966 ;
  assign n967 = n896 & n1506 ;
  assign n1507 = ~n967 ;
  assign n968 = n965 & n1507 ;
  assign n969 = x27 | n968 ;
  assign n841 = n839 & n1455 ;
  assign n946 = n841 & n35 ;
  assign n1508 = ~n846 ;
  assign n947 = n1508 & n946 ;
  assign n1509 = ~n946 ;
  assign n948 = n846 & n1509 ;
  assign n949 = n947 | n948 ;
  assign n970 = x27 & n968 ;
  assign n1510 = ~n970 ;
  assign n971 = n949 & n1510 ;
  assign n1511 = ~n971 ;
  assign n972 = n969 & n1511 ;
  assign n973 = x28 | n972 ;
  assign n974 = x28 & n972 ;
  assign n851 = n849 & n1459 ;
  assign n917 = n851 & n35 ;
  assign n1512 = ~n861 ;
  assign n918 = n1512 & n917 ;
  assign n1513 = ~n917 ;
  assign n983 = n861 & n1513 ;
  assign n984 = n918 | n983 ;
  assign n1514 = ~n974 ;
  assign n985 = n1514 & n984 ;
  assign n1515 = ~n985 ;
  assign n986 = n973 & n1515 ;
  assign n987 = x29 | n986 ;
  assign n978 = n864 & n1463 ;
  assign n979 = n35 & n978 ;
  assign n1516 = ~n856 ;
  assign n980 = n1516 & n979 ;
  assign n1517 = ~n979 ;
  assign n981 = n856 & n1517 ;
  assign n982 = n980 | n981 ;
  assign n988 = x29 & n986 ;
  assign n1518 = ~n988 ;
  assign n989 = n982 & n1518 ;
  assign n1519 = ~n989 ;
  assign n990 = n987 & n1519 ;
  assign n991 = x30 & n990 ;
  assign n992 = x30 | n990 ;
  assign n1520 = ~n991 ;
  assign n994 = n1520 & n992 ;
  assign n1521 = ~n994 ;
  assign n995 = n875 & n1521 ;
  assign n1522 = ~n873 ;
  assign n874 = x31 & n1522 ;
  assign n993 = n1522 & n992 ;
  assign n996 = x31 | n991 ;
  assign n997 = n993 | n996 ;
  assign n1095 = n987 & n1518 ;
  assign n34 = ~n997 ;
  assign n1096 = n34 & n1095 ;
  assign n1524 = ~n982 ;
  assign n1097 = n1524 & n1096 ;
  assign n1525 = ~n1096 ;
  assign n1098 = n982 & n1525 ;
  assign n1099 = n1097 | n1098 ;
  assign n1526 = ~n1099 ;
  assign n1100 = x30 & n1526 ;
  assign n1101 = n874 | n1100 ;
  assign n976 = n969 & n1510 ;
  assign n998 = n976 & n34 ;
  assign n1527 = ~n949 ;
  assign n999 = n1527 & n998 ;
  assign n1528 = ~n998 ;
  assign n1000 = n949 & n1528 ;
  assign n1001 = n999 | n1000 ;
  assign n1529 = ~x28 ;
  assign n1003 = n1529 & n1001 ;
  assign n977 = n965 & n1506 ;
  assign n1071 = n977 & n34 ;
  assign n1072 = n896 | n1071 ;
  assign n1073 = n896 & n1071 ;
  assign n1530 = ~n1073 ;
  assign n1074 = n1072 & n1530 ;
  assign n1531 = ~x27 ;
  assign n1075 = n1531 & n1074 ;
  assign n1076 = n1003 | n1075 ;
  assign n1532 = ~n1074 ;
  assign n1077 = x27 & n1532 ;
  assign n958 = n956 & n1502 ;
  assign n1054 = n958 & n34 ;
  assign n1533 = ~n962 ;
  assign n1055 = n1533 & n1054 ;
  assign n1534 = ~n1054 ;
  assign n1056 = n962 & n1534 ;
  assign n1057 = n1055 | n1056 ;
  assign n1535 = ~x26 ;
  assign n1060 = n1535 & n1057 ;
  assign n945 = n943 & n1498 ;
  assign n1038 = n945 & n34 ;
  assign n1536 = ~n953 ;
  assign n1039 = n1536 & n1038 ;
  assign n1537 = ~n1038 ;
  assign n1040 = n953 & n1537 ;
  assign n1041 = n1039 | n1040 ;
  assign n1538 = ~n1041 ;
  assign n1044 = x25 & n1538 ;
  assign n1539 = ~n1057 ;
  assign n1058 = x26 & n1539 ;
  assign n1059 = n1044 | n1058 ;
  assign n936 = n934 & n1494 ;
  assign n1004 = n936 & n34 ;
  assign n1005 = n940 | n1004 ;
  assign n1006 = n940 & n1004 ;
  assign n1540 = ~n1006 ;
  assign n1007 = n1005 & n1540 ;
  assign n1541 = ~x24 ;
  assign n1008 = n1541 & n1007 ;
  assign n1542 = ~x25 ;
  assign n1042 = n1542 & n1041 ;
  assign n1043 = n1008 | n1042 ;
  assign n1543 = ~n1007 ;
  assign n1009 = x24 & n1543 ;
  assign n927 = n925 & n1490 ;
  assign n1024 = n927 & n34 ;
  assign n1544 = ~n931 ;
  assign n1025 = n1544 & n1024 ;
  assign n1545 = ~n1024 ;
  assign n1026 = n931 & n1545 ;
  assign n1027 = n1025 | n1026 ;
  assign n1546 = ~n1027 ;
  assign n1028 = x23 & n1546 ;
  assign n1029 = n1009 | n1028 ;
  assign n1547 = ~x23 ;
  assign n1030 = n1547 & n1027 ;
  assign n916 = n914 & n1487 ;
  assign n1031 = n916 & n34 ;
  assign n1548 = ~n922 ;
  assign n1032 = n1548 & n1031 ;
  assign n1549 = ~n1031 ;
  assign n1033 = n922 & n1549 ;
  assign n1034 = n1032 | n1033 ;
  assign n1550 = ~x22 ;
  assign n1036 = n1550 & n1034 ;
  assign n1037 = n1030 | n1036 ;
  assign n1551 = ~n1034 ;
  assign n1035 = x22 & n1551 ;
  assign n883 = n881 | n882 ;
  assign n1053 = n911 & n34 ;
  assign n1078 = x20 & n997 ;
  assign n1079 = n1053 | n1078 ;
  assign n1552 = ~n883 ;
  assign n1080 = n1552 & n1079 ;
  assign n1553 = ~n1079 ;
  assign n1081 = n883 & n1553 ;
  assign n1082 = n1080 | n1081 ;
  assign n1554 = ~n1082 ;
  assign n1083 = x21 & n1554 ;
  assign n1084 = n1035 | n1083 ;
  assign n905 = n903 & n1482 ;
  assign n1012 = n905 & n34 ;
  assign n1013 = n909 & n1012 ;
  assign n1014 = n909 | n1012 ;
  assign n1555 = ~n1013 ;
  assign n1015 = n1555 & n1014 ;
  assign n1556 = ~n1015 ;
  assign n1016 = x20 & n1556 ;
  assign n52 = n1475 & n50 ;
  assign n1045 = n52 & n34 ;
  assign n1046 = n887 & n1045 ;
  assign n1047 = n887 | n1045 ;
  assign n1557 = ~n1046 ;
  assign n1048 = n1557 & n1047 ;
  assign n1049 = n1262 & n1048 ;
  assign n1558 = ~x0 ;
  assign n53 = n1558 & x16 ;
  assign n54 = x17 & n53 ;
  assign n1018 = x16 & n34 ;
  assign n1559 = ~n1018 ;
  assign n1019 = x1 & n1559 ;
  assign n55 = x17 | n53 ;
  assign n1020 = n1473 & n1018 ;
  assign n1560 = ~n1020 ;
  assign n1021 = n55 & n1560 ;
  assign n1561 = ~n1019 ;
  assign n1022 = n1561 & n1021 ;
  assign n1023 = n54 | n1022 ;
  assign n1562 = ~n1048 ;
  assign n1050 = x18 & n1562 ;
  assign n1051 = n1023 | n1050 ;
  assign n1563 = ~n1049 ;
  assign n1052 = n1563 & n1051 ;
  assign n892 = n1478 & n891 ;
  assign n1061 = n892 & n34 ;
  assign n1564 = ~n900 ;
  assign n1062 = n1564 & n1061 ;
  assign n1565 = ~n1061 ;
  assign n1063 = n900 & n1565 ;
  assign n1064 = n1062 | n1063 ;
  assign n1566 = ~n1064 ;
  assign n1065 = x19 & n1566 ;
  assign n1066 = n1052 | n1065 ;
  assign n1017 = n1273 & n1015 ;
  assign n1067 = n1207 & n1064 ;
  assign n1068 = n1017 | n1067 ;
  assign n1567 = ~n1068 ;
  assign n1069 = n1066 & n1567 ;
  assign n1070 = n1016 | n1069 ;
  assign n1568 = ~x21 ;
  assign n1085 = n1568 & n1082 ;
  assign n1569 = ~n1085 ;
  assign n1086 = n1070 & n1569 ;
  assign n1087 = n1084 | n1086 ;
  assign n1570 = ~n1037 ;
  assign n1088 = n1570 & n1087 ;
  assign n1089 = n1029 | n1088 ;
  assign n1571 = ~n1043 ;
  assign n1090 = n1571 & n1089 ;
  assign n1091 = n1059 | n1090 ;
  assign n1572 = ~n1060 ;
  assign n1092 = n1572 & n1091 ;
  assign n1093 = n1077 | n1092 ;
  assign n1573 = ~n1076 ;
  assign n1094 = n1573 & n1093 ;
  assign n1574 = ~n1001 ;
  assign n1002 = x28 & n1574 ;
  assign n975 = n973 & n1514 ;
  assign n1010 = n975 & n34 ;
  assign n1575 = ~n984 ;
  assign n1011 = n1575 & n1010 ;
  assign n1576 = ~n1010 ;
  assign n1103 = n984 & n1576 ;
  assign n1104 = n1011 | n1103 ;
  assign n1577 = ~n1104 ;
  assign n1105 = x29 & n1577 ;
  assign n1106 = n1002 | n1105 ;
  assign n1107 = n1094 | n1106 ;
  assign n1578 = ~x30 ;
  assign n1102 = n1578 & n1099 ;
  assign n1579 = ~x29 ;
  assign n1108 = n1579 & n1104 ;
  assign n1109 = n1102 | n1108 ;
  assign n1580 = ~n1109 ;
  assign n1110 = n1107 & n1580 ;
  assign n1111 = n1101 | n1110 ;
  assign n1581 = ~n995 ;
  assign n1112 = n1581 & n1111 ;
  assign n70 = n1119 & x16 ;
  assign n71 = n69 | n70 ;
  assign n33 = ~n1112 ;
  assign n48 = ~n71 ;
  assign y0 = n33 ;
  assign y1 = n34 ;
  assign y2 = n35 ;
  assign y3 = n36 ;
  assign y4 = n37 ;
  assign y5 = n38 ;
  assign y6 = n39 ;
  assign y7 = n40 ;
  assign y8 = n41 ;
  assign y9 = n42 ;
  assign y10 = n43 ;
  assign y11 = n44 ;
  assign y12 = n45 ;
  assign y13 = n46 ;
  assign y14 = n47 ;
  assign y15 = n48 ;
endmodule
