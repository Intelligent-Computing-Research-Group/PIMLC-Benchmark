module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 ;
  assign n65 = x0 & x32 ;
  assign n1324 = x1 & x32 ;
  assign n530 = x0 & x33 ;
  assign n4273 = ~n530 ;
  assign n757 = n1324 & n4273 ;
  assign n4274 = ~n1324 ;
  assign n4247 = n4274 & n530 ;
  assign n66 = n757 | n4247 ;
  assign n526 = x0 & x34 ;
  assign n527 = x1 & x33 ;
  assign n4249 = x32 | n527 ;
  assign n4275 = ~x2 ;
  assign n4250 = n4275 & n65 ;
  assign n4276 = ~n4250 ;
  assign n4251 = n4249 & n4276 ;
  assign n4252 = n526 & n4251 ;
  assign n4255 = x34 | n4251 ;
  assign n528 = x2 & x32 ;
  assign n4277 = ~n528 ;
  assign n753 = n527 & n4277 ;
  assign n4278 = ~n527 ;
  assign n4253 = n4278 & n528 ;
  assign n4254 = x0 | n4253 ;
  assign n4256 = n753 | n4254 ;
  assign n4257 = n4255 & n4256 ;
  assign n4279 = ~n4252 ;
  assign n67 = n4279 & n4257 ;
  assign n529 = x1 & x34 ;
  assign n771 = x2 & x34 ;
  assign n754 = n771 | n753 ;
  assign n755 = n65 & n754 ;
  assign n756 = n529 | n755 ;
  assign n758 = n530 | n755 ;
  assign n759 = n529 & n758 ;
  assign n4280 = ~n759 ;
  assign n760 = n756 & n4280 ;
  assign n1417 = x0 & x35 ;
  assign n1519 = x3 & x32 ;
  assign n531 = n1417 & n1519 ;
  assign n761 = n1417 | n1519 ;
  assign n4281 = ~n531 ;
  assign n762 = n4281 & n761 ;
  assign n764 = n1324 & n762 ;
  assign n1630 = x2 & x33 ;
  assign n763 = n1630 & n762 ;
  assign n765 = n1630 | n762 ;
  assign n4282 = ~n763 ;
  assign n766 = n4282 & n765 ;
  assign n767 = n4274 & n766 ;
  assign n768 = n764 | n767 ;
  assign n4283 = ~n760 ;
  assign n769 = n4283 & n768 ;
  assign n4284 = ~n768 ;
  assign n770 = n760 & n4284 ;
  assign n68 = n769 | n770 ;
  assign n4285 = ~n1630 ;
  assign n1169 = n4285 & n762 ;
  assign n4286 = ~n1169 ;
  assign n1170 = n761 & n4286 ;
  assign n139 = x0 & x36 ;
  assign n140 = n771 & n139 ;
  assign n1171 = n771 | n139 ;
  assign n4287 = ~n140 ;
  assign n1172 = n4287 & n1171 ;
  assign n1173 = n1170 & n1172 ;
  assign n1174 = n1170 | n1172 ;
  assign n4288 = ~n1173 ;
  assign n1175 = n4288 & n1174 ;
  assign n564 = x3 & x33 ;
  assign n135 = x4 & x35 ;
  assign n567 = n1324 & n135 ;
  assign n565 = x4 & x32 ;
  assign n566 = x1 & x35 ;
  assign n1130 = n565 | n566 ;
  assign n4289 = ~n567 ;
  assign n1131 = n4289 & n1130 ;
  assign n4290 = ~n564 ;
  assign n1132 = n4290 & n1131 ;
  assign n4291 = ~n1131 ;
  assign n1176 = n564 & n4291 ;
  assign n1177 = n1132 | n1176 ;
  assign n1178 = n1175 | n1177 ;
  assign n1179 = n1175 & n1177 ;
  assign n4292 = ~n1179 ;
  assign n1198 = n1178 & n4292 ;
  assign n569 = n1324 & n1630 ;
  assign n4293 = ~n68 ;
  assign n1194 = n569 & n4293 ;
  assign n1195 = n756 & n766 ;
  assign n1196 = n759 | n1195 ;
  assign n1197 = n1194 | n1196 ;
  assign n1199 = n1194 & n1196 ;
  assign n4294 = ~n1199 ;
  assign n4259 = n1197 & n4294 ;
  assign n4260 = n1198 & n4259 ;
  assign n4261 = n1198 | n4259 ;
  assign n4295 = ~n4260 ;
  assign n69 = n4295 & n4261 ;
  assign n1200 = n1198 | n1199 ;
  assign n1201 = n1197 & n1200 ;
  assign n561 = x4 & x33 ;
  assign n130 = x5 & x32 ;
  assign n131 = x2 & x35 ;
  assign n562 = n130 & n131 ;
  assign n1090 = n130 | n131 ;
  assign n4296 = ~n562 ;
  assign n1091 = n4296 & n1090 ;
  assign n4297 = ~n561 ;
  assign n1092 = n4297 & n1091 ;
  assign n4298 = ~n1091 ;
  assign n1141 = n561 & n4298 ;
  assign n1142 = n1092 | n1141 ;
  assign n1133 = n564 & n1131 ;
  assign n1134 = n567 | n1133 ;
  assign n138 = x3 & x34 ;
  assign n136 = x0 & x37 ;
  assign n137 = x1 & x36 ;
  assign n568 = n136 & n137 ;
  assign n1135 = n136 | n137 ;
  assign n4299 = ~n568 ;
  assign n1136 = n4299 & n1135 ;
  assign n1137 = n138 & n1136 ;
  assign n1138 = n138 | n1136 ;
  assign n4300 = ~n1137 ;
  assign n1139 = n4300 & n1138 ;
  assign n1140 = n1134 | n1139 ;
  assign n1143 = n1134 & n1139 ;
  assign n4301 = ~n1143 ;
  assign n1144 = n1140 & n4301 ;
  assign n4302 = ~n1142 ;
  assign n1145 = n4302 & n1144 ;
  assign n4303 = ~n1144 ;
  assign n1181 = n1142 & n4303 ;
  assign n1182 = n1145 | n1181 ;
  assign n1180 = n140 & n1179 ;
  assign n1183 = n140 | n1179 ;
  assign n4304 = ~n1180 ;
  assign n1184 = n4304 & n1183 ;
  assign n1185 = n1173 | n1184 ;
  assign n1186 = n1182 | n1185 ;
  assign n1187 = n1182 & n1185 ;
  assign n4305 = ~n1187 ;
  assign n1202 = n1186 & n4305 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = n1201 & n1202 ;
  assign n4306 = ~n1204 ;
  assign n70 = n1203 & n4306 ;
  assign n1188 = n1180 | n1187 ;
  assign n126 = x0 & x38 ;
  assign n4307 = ~n138 ;
  assign n1148 = n4307 & n1136 ;
  assign n4308 = ~n1148 ;
  assign n1149 = n1135 & n4308 ;
  assign n1150 = n126 & n1149 ;
  assign n1161 = n126 | n1149 ;
  assign n4309 = ~n1150 ;
  assign n1162 = n4309 & n1161 ;
  assign n132 = x2 & x36 ;
  assign n133 = x1 & x37 ;
  assign n134 = x4 & x34 ;
  assign n563 = n133 & n134 ;
  assign n1097 = n133 | n134 ;
  assign n4310 = ~n563 ;
  assign n1098 = n4310 & n1097 ;
  assign n1099 = n132 & n1098 ;
  assign n1100 = n132 | n1098 ;
  assign n4311 = ~n1099 ;
  assign n1101 = n4311 & n1100 ;
  assign n4312 = ~n1092 ;
  assign n1093 = n1090 & n4312 ;
  assign n129 = x3 & x35 ;
  assign n127 = x5 & x33 ;
  assign n128 = x6 & x32 ;
  assign n560 = n127 & n128 ;
  assign n1049 = n127 | n128 ;
  assign n4313 = ~n560 ;
  assign n1050 = n4313 & n1049 ;
  assign n1051 = n129 & n1050 ;
  assign n1094 = n129 | n1050 ;
  assign n4314 = ~n1051 ;
  assign n1095 = n4314 & n1094 ;
  assign n1096 = n1093 | n1095 ;
  assign n1102 = n1093 & n1095 ;
  assign n4315 = ~n1102 ;
  assign n1103 = n1096 & n4315 ;
  assign n4316 = ~n1101 ;
  assign n1104 = n4316 & n1103 ;
  assign n4317 = ~n1103 ;
  assign n1128 = n1101 & n4317 ;
  assign n1129 = n1104 | n1128 ;
  assign n4318 = ~n1145 ;
  assign n1146 = n1140 & n4318 ;
  assign n1147 = n1129 & n1146 ;
  assign n1160 = n1129 | n1146 ;
  assign n4319 = ~n1147 ;
  assign n1189 = n4319 & n1160 ;
  assign n4320 = ~n1189 ;
  assign n1190 = n1162 & n4320 ;
  assign n4321 = ~n1162 ;
  assign n1191 = n4321 & n1189 ;
  assign n1192 = n1190 | n1191 ;
  assign n1193 = n1188 | n1192 ;
  assign n1205 = n1188 & n1192 ;
  assign n4322 = ~n1205 ;
  assign n1206 = n1193 & n4322 ;
  assign n1207 = n4306 & n1206 ;
  assign n4323 = ~n1206 ;
  assign n4264 = n1204 & n4323 ;
  assign n71 = n1207 | n4264 ;
  assign n4324 = ~n1207 ;
  assign n1208 = n1193 & n4324 ;
  assign n119 = x6 & x33 ;
  assign n120 = x7 & x32 ;
  assign n557 = n119 & n120 ;
  assign n984 = n119 | n120 ;
  assign n4325 = ~n557 ;
  assign n985 = n4325 & n984 ;
  assign n4326 = ~n135 ;
  assign n986 = n4326 & n985 ;
  assign n4327 = ~n985 ;
  assign n1047 = n135 & n4327 ;
  assign n1048 = n986 | n1047 ;
  assign n4328 = ~n129 ;
  assign n1052 = n4328 & n1050 ;
  assign n4329 = ~n1052 ;
  assign n1053 = n1049 & n4329 ;
  assign n4330 = ~n1048 ;
  assign n1054 = n4330 & n1053 ;
  assign n4331 = ~n1053 ;
  assign n1056 = n1048 & n4331 ;
  assign n1057 = n1054 | n1056 ;
  assign n123 = x3 & x36 ;
  assign n121 = x2 & x37 ;
  assign n122 = x5 & x34 ;
  assign n558 = n121 & n122 ;
  assign n1028 = n121 | n122 ;
  assign n4332 = ~n558 ;
  assign n1029 = n4332 & n1028 ;
  assign n4333 = ~n1029 ;
  assign n1030 = n123 & n4333 ;
  assign n4334 = ~n123 ;
  assign n1031 = n4334 & n1029 ;
  assign n1058 = n1030 | n1031 ;
  assign n4335 = ~n1058 ;
  assign n1059 = n1057 & n4335 ;
  assign n4336 = ~n1057 ;
  assign n1088 = n4336 & n1058 ;
  assign n1089 = n1059 | n1088 ;
  assign n4337 = ~n1104 ;
  assign n1105 = n1096 & n4337 ;
  assign n4338 = ~n1089 ;
  assign n1106 = n4338 & n1105 ;
  assign n4339 = ~n1105 ;
  assign n1112 = n1089 & n4339 ;
  assign n1113 = n1106 | n1112 ;
  assign n124 = x0 & x39 ;
  assign n125 = x1 & x38 ;
  assign n559 = n124 & n125 ;
  assign n1033 = n124 | n125 ;
  assign n4340 = ~n559 ;
  assign n1034 = n4340 & n1033 ;
  assign n4341 = ~n132 ;
  assign n1108 = n4341 & n1098 ;
  assign n4342 = ~n1108 ;
  assign n1109 = n1097 & n4342 ;
  assign n1110 = n1034 & n1109 ;
  assign n1111 = n1034 | n1109 ;
  assign n4343 = ~n1110 ;
  assign n1156 = n4343 & n1111 ;
  assign n1157 = n1113 | n1156 ;
  assign n1158 = n1113 & n1156 ;
  assign n4344 = ~n1158 ;
  assign n1159 = n1157 & n4344 ;
  assign n1151 = n1147 & n1150 ;
  assign n1163 = n1147 | n1162 ;
  assign n1164 = n1160 & n1163 ;
  assign n1165 = n1150 | n1164 ;
  assign n4345 = ~n1151 ;
  assign n1166 = n4345 & n1165 ;
  assign n1167 = n1159 & n1166 ;
  assign n1168 = n1159 | n1166 ;
  assign n4346 = ~n1167 ;
  assign n1209 = n4346 & n1168 ;
  assign n4347 = ~n1209 ;
  assign n1210 = n1208 & n4347 ;
  assign n4348 = ~n1208 ;
  assign n1211 = n4348 & n1209 ;
  assign n72 = n1210 | n1211 ;
  assign n4349 = ~n1211 ;
  assign n1212 = n1168 & n4349 ;
  assign n1055 = n1048 & n1053 ;
  assign n1060 = n1057 & n1058 ;
  assign n1061 = n1055 | n1060 ;
  assign n4350 = ~n1031 ;
  assign n1032 = n1028 & n4350 ;
  assign n115 = x1 & x39 ;
  assign n113 = x0 & x40 ;
  assign n114 = x2 & x38 ;
  assign n966 = n113 | n114 ;
  assign n967 = n115 & n966 ;
  assign n1035 = n967 & n1034 ;
  assign n2815 = x2 & x40 ;
  assign n4351 = ~n2815 ;
  assign n1036 = n4351 & n966 ;
  assign n4352 = ~n1036 ;
  assign n1037 = n126 & n4352 ;
  assign n1038 = n115 | n966 ;
  assign n4353 = ~n1037 ;
  assign n1039 = n4353 & n1038 ;
  assign n4354 = ~n1035 ;
  assign n1040 = n4354 & n1039 ;
  assign n1041 = n1032 & n1040 ;
  assign n1042 = n1032 | n1040 ;
  assign n4355 = ~n1041 ;
  assign n1043 = n4355 & n1042 ;
  assign n118 = x4 & x36 ;
  assign n116 = x6 & x34 ;
  assign n117 = x3 & x37 ;
  assign n556 = n116 & n117 ;
  assign n972 = n116 | n117 ;
  assign n4356 = ~n556 ;
  assign n973 = n4356 & n972 ;
  assign n974 = n118 & n973 ;
  assign n992 = n118 | n973 ;
  assign n4357 = ~n974 ;
  assign n993 = n4357 & n992 ;
  assign n4358 = ~n986 ;
  assign n987 = n984 & n4358 ;
  assign n552 = x7 & x33 ;
  assign n109 = x5 & x35 ;
  assign n110 = x8 & x32 ;
  assign n553 = n109 & n110 ;
  assign n925 = n109 | n110 ;
  assign n4359 = ~n553 ;
  assign n926 = n4359 & n925 ;
  assign n4360 = ~n552 ;
  assign n927 = n4360 & n926 ;
  assign n4361 = ~n926 ;
  assign n988 = n552 & n4361 ;
  assign n989 = n927 | n988 ;
  assign n990 = n987 | n989 ;
  assign n991 = n987 & n989 ;
  assign n4362 = ~n991 ;
  assign n994 = n990 & n4362 ;
  assign n995 = n993 & n994 ;
  assign n1044 = n993 | n994 ;
  assign n4363 = ~n995 ;
  assign n1045 = n4363 & n1044 ;
  assign n1046 = n1043 & n1045 ;
  assign n1062 = n1043 | n1045 ;
  assign n4364 = ~n1046 ;
  assign n1063 = n4364 & n1062 ;
  assign n1064 = n1061 & n1063 ;
  assign n1117 = n1061 | n1063 ;
  assign n4365 = ~n1064 ;
  assign n1118 = n4365 & n1117 ;
  assign n1107 = n1089 & n1105 ;
  assign n1115 = n1107 & n4343 ;
  assign n1114 = n1110 | n1113 ;
  assign n1116 = n1111 & n1114 ;
  assign n4366 = ~n1107 ;
  assign n1119 = n4366 & n1116 ;
  assign n1120 = n1115 | n1119 ;
  assign n4367 = ~n1118 ;
  assign n1121 = n4367 & n1120 ;
  assign n4368 = ~n1120 ;
  assign n1152 = n1118 & n4368 ;
  assign n1153 = n1121 | n1152 ;
  assign n4369 = ~n1153 ;
  assign n1154 = n1151 & n4369 ;
  assign n1213 = n4345 & n1153 ;
  assign n1214 = n1154 | n1213 ;
  assign n1215 = n1212 | n1214 ;
  assign n1216 = n1212 & n1214 ;
  assign n4370 = ~n1216 ;
  assign n73 = n1215 & n4370 ;
  assign n1155 = n1151 & n1153 ;
  assign n1217 = n1155 | n1216 ;
  assign n1122 = n1107 | n1116 ;
  assign n4371 = ~n1121 ;
  assign n1123 = n4371 & n1122 ;
  assign n102 = x8 & x33 ;
  assign n100 = x9 & x32 ;
  assign n101 = x6 & x35 ;
  assign n549 = n100 & n101 ;
  assign n877 = n100 | n101 ;
  assign n4372 = ~n549 ;
  assign n878 = n4372 & n877 ;
  assign n879 = n102 & n878 ;
  assign n932 = n102 | n878 ;
  assign n4373 = ~n879 ;
  assign n933 = n4373 & n932 ;
  assign n4374 = ~n927 ;
  assign n928 = n925 & n4374 ;
  assign n108 = x5 & x36 ;
  assign n106 = x4 & x37 ;
  assign n107 = x7 & x34 ;
  assign n551 = n106 & n107 ;
  assign n912 = n106 | n107 ;
  assign n4375 = ~n551 ;
  assign n913 = n4375 & n912 ;
  assign n914 = n108 & n913 ;
  assign n929 = n108 | n913 ;
  assign n4376 = ~n914 ;
  assign n930 = n4376 & n929 ;
  assign n931 = n928 | n930 ;
  assign n934 = n928 & n930 ;
  assign n4377 = ~n934 ;
  assign n935 = n931 & n4377 ;
  assign n4378 = ~n933 ;
  assign n936 = n4378 & n935 ;
  assign n4379 = ~n935 ;
  assign n998 = n933 & n4379 ;
  assign n999 = n936 | n998 ;
  assign n4380 = ~n118 ;
  assign n975 = n4380 & n973 ;
  assign n4381 = ~n975 ;
  assign n976 = n972 & n4381 ;
  assign n555 = n113 & n114 ;
  assign n968 = n555 | n967 ;
  assign n105 = x1 & x40 ;
  assign n103 = x2 & x39 ;
  assign n104 = x3 & x38 ;
  assign n550 = n103 & n104 ;
  assign n907 = n103 | n104 ;
  assign n4382 = ~n550 ;
  assign n908 = n4382 & n907 ;
  assign n4383 = ~n908 ;
  assign n909 = n105 & n4383 ;
  assign n4384 = ~n105 ;
  assign n910 = n4384 & n908 ;
  assign n969 = n909 | n910 ;
  assign n970 = n968 | n969 ;
  assign n971 = n968 & n969 ;
  assign n4385 = ~n971 ;
  assign n977 = n970 & n4385 ;
  assign n978 = n976 & n977 ;
  assign n982 = n976 | n977 ;
  assign n4386 = ~n978 ;
  assign n983 = n4386 & n982 ;
  assign n996 = n991 | n995 ;
  assign n997 = n983 | n996 ;
  assign n1000 = n983 & n996 ;
  assign n4387 = ~n1000 ;
  assign n1001 = n997 & n4387 ;
  assign n4388 = ~n999 ;
  assign n1002 = n4388 & n1001 ;
  assign n4389 = ~n1001 ;
  assign n1026 = n999 & n4389 ;
  assign n1027 = n1002 | n1026 ;
  assign n1065 = n1046 | n1064 ;
  assign n1066 = n1027 | n1065 ;
  assign n1067 = n1027 & n1065 ;
  assign n4390 = ~n1067 ;
  assign n1073 = n1066 & n4390 ;
  assign n536 = x0 & x41 ;
  assign n1068 = n115 & n1037 ;
  assign n1069 = n1041 | n1068 ;
  assign n1070 = n536 | n1069 ;
  assign n1071 = n536 & n1069 ;
  assign n4391 = ~n1071 ;
  assign n1074 = n1070 & n4391 ;
  assign n1075 = n1073 & n1074 ;
  assign n1124 = n1073 | n1074 ;
  assign n4392 = ~n1075 ;
  assign n1125 = n4392 & n1124 ;
  assign n4393 = ~n1123 ;
  assign n1126 = n4393 & n1125 ;
  assign n4394 = ~n1125 ;
  assign n1218 = n1123 & n4394 ;
  assign n1219 = n1126 | n1218 ;
  assign n4395 = ~n1219 ;
  assign n1220 = n1217 & n4395 ;
  assign n4396 = ~n1217 ;
  assign n1221 = n4396 & n1219 ;
  assign n74 = n1220 | n1221 ;
  assign n1127 = n1123 | n1125 ;
  assign n4397 = ~n1221 ;
  assign n1222 = n1127 & n4397 ;
  assign n1072 = n1067 & n1071 ;
  assign n1076 = n1067 | n1071 ;
  assign n4398 = ~n1072 ;
  assign n1077 = n4398 & n1076 ;
  assign n1078 = n1075 | n1077 ;
  assign n1003 = n999 & n1001 ;
  assign n1004 = n1000 | n1003 ;
  assign n3797 = x5 & x37 ;
  assign n3394 = x8 & x34 ;
  assign n3592 = x6 & x36 ;
  assign n540 = n3394 & n3592 ;
  assign n799 = n3394 | n3592 ;
  assign n4399 = ~n540 ;
  assign n800 = n4399 & n799 ;
  assign n801 = n3797 & n800 ;
  assign n885 = n3797 | n800 ;
  assign n4400 = ~n801 ;
  assign n886 = n4400 & n885 ;
  assign n4401 = ~n102 ;
  assign n880 = n4401 & n878 ;
  assign n4402 = ~n880 ;
  assign n881 = n877 & n4402 ;
  assign n4248 = x9 & x33 ;
  assign n4007 = x7 & x35 ;
  assign n4246 = x10 & x32 ;
  assign n541 = n4007 & n4246 ;
  assign n816 = n4007 | n4246 ;
  assign n4403 = ~n541 ;
  assign n817 = n4403 & n816 ;
  assign n818 = n4248 & n817 ;
  assign n882 = n4248 | n817 ;
  assign n4404 = ~n818 ;
  assign n883 = n4404 & n882 ;
  assign n884 = n881 | n883 ;
  assign n887 = n881 & n883 ;
  assign n4405 = ~n887 ;
  assign n888 = n884 & n4405 ;
  assign n889 = n886 & n888 ;
  assign n939 = n886 | n888 ;
  assign n4406 = ~n889 ;
  assign n940 = n4406 & n939 ;
  assign n4407 = ~n910 ;
  assign n911 = n907 & n4407 ;
  assign n4408 = ~n108 ;
  assign n915 = n4408 & n913 ;
  assign n4409 = ~n915 ;
  assign n916 = n912 & n4409 ;
  assign n4410 = ~n911 ;
  assign n917 = n4410 & n916 ;
  assign n4411 = ~n916 ;
  assign n918 = n911 & n4411 ;
  assign n919 = n917 | n918 ;
  assign n2463 = x3 & x39 ;
  assign n2639 = x4 & x38 ;
  assign n537 = n2463 & n2639 ;
  assign n788 = n2463 | n2639 ;
  assign n4412 = ~n537 ;
  assign n789 = n4412 & n788 ;
  assign n790 = n4351 & n789 ;
  assign n4413 = ~n789 ;
  assign n920 = n2815 & n4413 ;
  assign n921 = n790 | n920 ;
  assign n922 = n919 | n921 ;
  assign n923 = n919 & n921 ;
  assign n4414 = ~n923 ;
  assign n924 = n922 & n4414 ;
  assign n4415 = ~n936 ;
  assign n937 = n931 & n4415 ;
  assign n938 = n924 & n937 ;
  assign n941 = n924 | n937 ;
  assign n4416 = ~n938 ;
  assign n942 = n4416 & n941 ;
  assign n943 = n940 & n942 ;
  assign n1005 = n940 | n942 ;
  assign n4417 = ~n943 ;
  assign n1006 = n4417 & n1005 ;
  assign n111 = x0 & x42 ;
  assign n112 = x1 & x41 ;
  assign n554 = n111 & n112 ;
  assign n949 = n111 | n112 ;
  assign n4418 = ~n554 ;
  assign n950 = n4418 & n949 ;
  assign n979 = n971 | n978 ;
  assign n4419 = ~n979 ;
  assign n980 = n950 & n4419 ;
  assign n4420 = ~n950 ;
  assign n1007 = n4420 & n979 ;
  assign n1008 = n980 | n1007 ;
  assign n1009 = n1006 & n1008 ;
  assign n1010 = n1006 | n1008 ;
  assign n4421 = ~n1009 ;
  assign n1079 = n4421 & n1010 ;
  assign n1080 = n1004 & n1079 ;
  assign n1081 = n1004 | n1079 ;
  assign n4422 = ~n1080 ;
  assign n1082 = n4422 & n1081 ;
  assign n4423 = ~n1078 ;
  assign n1083 = n4423 & n1082 ;
  assign n4424 = ~n1082 ;
  assign n1223 = n1078 & n4424 ;
  assign n1224 = n1083 | n1223 ;
  assign n1225 = n1222 | n1224 ;
  assign n1226 = n1222 & n1224 ;
  assign n4425 = ~n1226 ;
  assign n75 = n1225 & n4425 ;
  assign n4265 = x11 & x32 ;
  assign n4266 = x8 & x35 ;
  assign n4267 = x10 & x33 ;
  assign n543 = n4266 & n4267 ;
  assign n827 = n4266 | n4267 ;
  assign n4426 = ~n543 ;
  assign n828 = n4426 & n827 ;
  assign n829 = n4265 & n828 ;
  assign n831 = n4265 | n828 ;
  assign n4427 = ~n829 ;
  assign n832 = n4427 & n831 ;
  assign n4428 = ~n4248 ;
  assign n819 = n4428 & n817 ;
  assign n4429 = ~n819 ;
  assign n820 = n816 & n4429 ;
  assign n4263 = x7 & x36 ;
  assign n4258 = x6 & x37 ;
  assign n4262 = x9 & x34 ;
  assign n542 = n4258 & n4262 ;
  assign n821 = n4258 | n4262 ;
  assign n4430 = ~n542 ;
  assign n822 = n4430 & n821 ;
  assign n823 = n4263 & n822 ;
  assign n824 = n4263 | n822 ;
  assign n4431 = ~n823 ;
  assign n825 = n4431 & n824 ;
  assign n826 = n820 | n825 ;
  assign n833 = n820 & n825 ;
  assign n4432 = ~n833 ;
  assign n834 = n826 & n4432 ;
  assign n835 = n832 & n834 ;
  assign n893 = n832 | n834 ;
  assign n4433 = ~n835 ;
  assign n894 = n4433 & n893 ;
  assign n4434 = ~n3797 ;
  assign n802 = n4434 & n800 ;
  assign n4435 = ~n802 ;
  assign n803 = n799 & n4435 ;
  assign n4436 = ~n790 ;
  assign n791 = n788 & n4436 ;
  assign n538 = x4 & x39 ;
  assign n3004 = x3 & x40 ;
  assign n3199 = x5 & x38 ;
  assign n539 = n3004 & n3199 ;
  assign n792 = n3004 | n3199 ;
  assign n4437 = ~n539 ;
  assign n793 = n4437 & n792 ;
  assign n4438 = ~n538 ;
  assign n794 = n4438 & n793 ;
  assign n4439 = ~n793 ;
  assign n795 = n538 & n4439 ;
  assign n796 = n794 | n795 ;
  assign n797 = n791 | n796 ;
  assign n798 = n791 & n796 ;
  assign n4440 = ~n798 ;
  assign n804 = n797 & n4440 ;
  assign n805 = n803 & n804 ;
  assign n875 = n803 | n804 ;
  assign n4441 = ~n805 ;
  assign n876 = n4441 & n875 ;
  assign n4442 = ~n886 ;
  assign n890 = n4442 & n888 ;
  assign n4443 = ~n890 ;
  assign n891 = n884 & n4443 ;
  assign n892 = n876 & n891 ;
  assign n895 = n876 | n891 ;
  assign n4444 = ~n892 ;
  assign n896 = n4444 & n895 ;
  assign n897 = n894 & n896 ;
  assign n905 = n894 | n896 ;
  assign n4445 = ~n897 ;
  assign n906 = n4445 & n905 ;
  assign n944 = n938 | n943 ;
  assign n4446 = ~n944 ;
  assign n945 = n906 & n4446 ;
  assign n4447 = ~n906 ;
  assign n957 = n4447 & n944 ;
  assign n958 = n945 | n957 ;
  assign n947 = n911 & n916 ;
  assign n948 = n923 | n947 ;
  assign n535 = x1 & x42 ;
  assign n533 = x0 & x43 ;
  assign n534 = x2 & x41 ;
  assign n777 = n533 | n534 ;
  assign n779 = n535 & n777 ;
  assign n951 = n779 & n950 ;
  assign n778 = n535 | n777 ;
  assign n2155 = x2 & x43 ;
  assign n4448 = ~n2155 ;
  assign n810 = n4448 & n777 ;
  assign n4449 = ~n810 ;
  assign n811 = n536 & n4449 ;
  assign n4450 = ~n811 ;
  assign n952 = n778 & n4450 ;
  assign n4451 = ~n951 ;
  assign n953 = n4451 & n952 ;
  assign n954 = n948 & n953 ;
  assign n956 = n948 | n953 ;
  assign n4452 = ~n954 ;
  assign n1013 = n4452 & n956 ;
  assign n4453 = ~n958 ;
  assign n1014 = n4453 & n1013 ;
  assign n4454 = ~n1013 ;
  assign n1015 = n958 & n4454 ;
  assign n1016 = n1014 | n1015 ;
  assign n981 = n950 & n979 ;
  assign n1011 = n1004 & n1010 ;
  assign n1012 = n981 & n1011 ;
  assign n1017 = n981 | n1011 ;
  assign n4455 = ~n1012 ;
  assign n1018 = n4455 & n1017 ;
  assign n1019 = n1009 | n1018 ;
  assign n1020 = n1016 | n1019 ;
  assign n1021 = n1016 & n1019 ;
  assign n4456 = ~n1021 ;
  assign n1025 = n1020 & n4456 ;
  assign n1084 = n1078 & n1082 ;
  assign n1085 = n1072 | n1084 ;
  assign n1086 = n1025 | n1085 ;
  assign n1087 = n1025 & n1085 ;
  assign n4457 = ~n1087 ;
  assign n1227 = n1086 & n4457 ;
  assign n1228 = n1226 | n1227 ;
  assign n1229 = n1226 & n1227 ;
  assign n4458 = ~n1229 ;
  assign n76 = n1228 & n4458 ;
  assign n1230 = n1087 | n1229 ;
  assign n1751 = x2 & x42 ;
  assign n1883 = x3 & x41 ;
  assign n2018 = x1 & x43 ;
  assign n532 = n1883 & n2018 ;
  assign n772 = n1883 | n2018 ;
  assign n4459 = ~n532 ;
  assign n773 = n4459 & n772 ;
  assign n774 = n1751 & n773 ;
  assign n775 = n1751 | n773 ;
  assign n4460 = ~n774 ;
  assign n776 = n4460 & n775 ;
  assign n2312 = x0 & x44 ;
  assign n780 = n2155 & n536 ;
  assign n781 = n779 | n780 ;
  assign n782 = n2312 & n781 ;
  assign n783 = n2312 | n781 ;
  assign n4461 = ~n782 ;
  assign n784 = n4461 & n783 ;
  assign n4462 = ~n776 ;
  assign n785 = n4462 & n784 ;
  assign n4463 = ~n784 ;
  assign n786 = n776 & n4463 ;
  assign n787 = n785 | n786 ;
  assign n806 = n798 | n805 ;
  assign n4464 = ~n806 ;
  assign n807 = n787 & n4464 ;
  assign n4465 = ~n787 ;
  assign n808 = n4465 & n806 ;
  assign n809 = n807 | n808 ;
  assign n812 = n535 & n811 ;
  assign n4466 = ~n809 ;
  assign n813 = n4466 & n812 ;
  assign n4467 = ~n812 ;
  assign n814 = n809 & n4467 ;
  assign n815 = n813 | n814 ;
  assign n4468 = ~n832 ;
  assign n836 = n4468 & n834 ;
  assign n4469 = ~n836 ;
  assign n837 = n826 & n4469 ;
  assign n4470 = ~n794 ;
  assign n838 = n792 & n4470 ;
  assign n4471 = ~n4263 ;
  assign n839 = n4471 & n822 ;
  assign n4472 = ~n839 ;
  assign n840 = n821 & n4472 ;
  assign n841 = n838 & n840 ;
  assign n842 = n838 | n840 ;
  assign n4473 = ~n841 ;
  assign n843 = n4473 & n842 ;
  assign n4270 = x5 & x39 ;
  assign n4268 = x4 & x40 ;
  assign n4269 = x6 & x38 ;
  assign n544 = n4268 & n4269 ;
  assign n844 = n4268 | n4269 ;
  assign n4474 = ~n544 ;
  assign n845 = n4474 & n844 ;
  assign n4475 = ~n845 ;
  assign n846 = n4270 & n4475 ;
  assign n4476 = ~n4270 ;
  assign n847 = n4476 & n845 ;
  assign n848 = n846 | n847 ;
  assign n4477 = ~n848 ;
  assign n849 = n843 & n4477 ;
  assign n4478 = ~n843 ;
  assign n850 = n4478 & n848 ;
  assign n851 = n849 | n850 ;
  assign n4479 = ~n4265 ;
  assign n830 = n4479 & n828 ;
  assign n4480 = ~n830 ;
  assign n852 = n827 & n4480 ;
  assign n545 = x7 & x37 ;
  assign n4272 = x8 & x36 ;
  assign n97 = x10 & x34 ;
  assign n546 = n4272 & n97 ;
  assign n853 = n4272 | n97 ;
  assign n4481 = ~n546 ;
  assign n854 = n4481 & n853 ;
  assign n4482 = ~n545 ;
  assign n855 = n4482 & n854 ;
  assign n4483 = ~n854 ;
  assign n856 = n545 & n4483 ;
  assign n857 = n855 | n856 ;
  assign n547 = x9 & x35 ;
  assign n98 = x11 & x33 ;
  assign n99 = x12 & x32 ;
  assign n548 = n98 & n99 ;
  assign n858 = n98 | n99 ;
  assign n4484 = ~n548 ;
  assign n859 = n4484 & n858 ;
  assign n4485 = ~n547 ;
  assign n860 = n4485 & n859 ;
  assign n4486 = ~n859 ;
  assign n861 = n547 & n4486 ;
  assign n862 = n860 | n861 ;
  assign n863 = n857 | n862 ;
  assign n864 = n857 & n862 ;
  assign n4487 = ~n864 ;
  assign n865 = n863 & n4487 ;
  assign n866 = n852 & n865 ;
  assign n867 = n852 | n865 ;
  assign n4488 = ~n866 ;
  assign n868 = n4488 & n867 ;
  assign n869 = n851 & n868 ;
  assign n870 = n851 | n868 ;
  assign n4489 = ~n869 ;
  assign n871 = n4489 & n870 ;
  assign n872 = n837 & n871 ;
  assign n873 = n837 | n871 ;
  assign n4490 = ~n872 ;
  assign n874 = n4490 & n873 ;
  assign n898 = n892 | n897 ;
  assign n899 = n874 | n898 ;
  assign n900 = n874 & n898 ;
  assign n4491 = ~n900 ;
  assign n901 = n899 & n4491 ;
  assign n902 = n815 & n901 ;
  assign n903 = n815 | n901 ;
  assign n4492 = ~n902 ;
  assign n904 = n4492 & n903 ;
  assign n946 = n906 & n944 ;
  assign n955 = n946 & n4452 ;
  assign n959 = n954 | n958 ;
  assign n960 = n956 & n959 ;
  assign n4493 = ~n946 ;
  assign n961 = n4493 & n960 ;
  assign n962 = n955 | n961 ;
  assign n4494 = ~n904 ;
  assign n963 = n4494 & n962 ;
  assign n4495 = ~n962 ;
  assign n964 = n904 & n4495 ;
  assign n965 = n963 | n964 ;
  assign n1022 = n1012 | n1021 ;
  assign n1023 = n965 | n1022 ;
  assign n1024 = n965 & n1022 ;
  assign n4496 = ~n1024 ;
  assign n1231 = n1023 & n4496 ;
  assign n1232 = n1230 & n1231 ;
  assign n4271 = n1230 | n1231 ;
  assign n4497 = ~n1232 ;
  assign n77 = n4497 & n4271 ;
  assign n1233 = n1024 | n1232 ;
  assign n4498 = ~n855 ;
  assign n1234 = n853 & n4498 ;
  assign n4499 = ~n847 ;
  assign n1235 = n844 & n4499 ;
  assign n1236 = n1234 & n1235 ;
  assign n1237 = n1234 | n1235 ;
  assign n4500 = ~n1236 ;
  assign n1238 = n4500 & n1237 ;
  assign n570 = x5 & x40 ;
  assign n141 = x6 & x39 ;
  assign n142 = x7 & x38 ;
  assign n571 = n141 & n142 ;
  assign n1239 = n141 | n142 ;
  assign n4501 = ~n571 ;
  assign n1240 = n4501 & n1239 ;
  assign n4502 = ~n570 ;
  assign n1241 = n4502 & n1240 ;
  assign n4503 = ~n1240 ;
  assign n1242 = n570 & n4503 ;
  assign n1243 = n1241 | n1242 ;
  assign n4504 = ~n1243 ;
  assign n1244 = n1238 & n4504 ;
  assign n4505 = ~n1238 ;
  assign n1245 = n4505 & n1243 ;
  assign n1246 = n1244 | n1245 ;
  assign n572 = x9 & x36 ;
  assign n143 = x11 & x34 ;
  assign n144 = x8 & x37 ;
  assign n573 = n143 & n144 ;
  assign n1247 = n143 | n144 ;
  assign n4506 = ~n573 ;
  assign n1248 = n4506 & n1247 ;
  assign n4507 = ~n572 ;
  assign n1249 = n4507 & n1248 ;
  assign n4508 = ~n1248 ;
  assign n1250 = n572 & n4508 ;
  assign n1251 = n1249 | n1250 ;
  assign n4509 = ~n860 ;
  assign n1252 = n858 & n4509 ;
  assign n574 = x12 & x33 ;
  assign n145 = x10 & x35 ;
  assign n146 = x13 & x32 ;
  assign n575 = n145 & n146 ;
  assign n1253 = n145 | n146 ;
  assign n4510 = ~n575 ;
  assign n1254 = n4510 & n1253 ;
  assign n4511 = ~n574 ;
  assign n1255 = n4511 & n1254 ;
  assign n4512 = ~n1254 ;
  assign n1256 = n574 & n4512 ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = n1252 | n1257 ;
  assign n1259 = n1252 & n1257 ;
  assign n4513 = ~n1259 ;
  assign n1260 = n1258 & n4513 ;
  assign n4514 = ~n1251 ;
  assign n1261 = n4514 & n1260 ;
  assign n4515 = ~n1260 ;
  assign n1262 = n1251 & n4515 ;
  assign n1263 = n1261 | n1262 ;
  assign n1264 = n864 | n866 ;
  assign n1265 = n1263 | n1264 ;
  assign n1266 = n1263 & n1264 ;
  assign n4516 = ~n1266 ;
  assign n1267 = n1265 & n4516 ;
  assign n4517 = ~n1246 ;
  assign n1268 = n4517 & n1267 ;
  assign n4518 = ~n1267 ;
  assign n1269 = n1246 & n4518 ;
  assign n1270 = n1268 | n1269 ;
  assign n1271 = n776 & n784 ;
  assign n1272 = n782 | n1271 ;
  assign n4519 = ~n1751 ;
  assign n1273 = n4519 & n773 ;
  assign n4520 = ~n1273 ;
  assign n1274 = n772 & n4520 ;
  assign n576 = x1 & x44 ;
  assign n577 = x0 & x45 ;
  assign n1275 = n576 | n577 ;
  assign n578 = x1 & x45 ;
  assign n1276 = n2312 & n578 ;
  assign n4521 = ~n1276 ;
  assign n1277 = n1275 & n4521 ;
  assign n147 = x3 & x42 ;
  assign n148 = x4 & x41 ;
  assign n579 = n147 & n148 ;
  assign n1278 = n147 | n148 ;
  assign n4522 = ~n579 ;
  assign n1279 = n4522 & n1278 ;
  assign n1280 = n2155 & n1279 ;
  assign n1281 = n2155 | n1279 ;
  assign n4523 = ~n1280 ;
  assign n1282 = n4523 & n1281 ;
  assign n1283 = n1277 & n1282 ;
  assign n1284 = n1277 | n1282 ;
  assign n4524 = ~n1283 ;
  assign n1285 = n4524 & n1284 ;
  assign n4525 = ~n1274 ;
  assign n1286 = n4525 & n1285 ;
  assign n4526 = ~n1285 ;
  assign n1287 = n1274 & n4526 ;
  assign n1288 = n1286 | n1287 ;
  assign n1289 = n843 & n848 ;
  assign n1290 = n841 | n1289 ;
  assign n1291 = n1288 | n1290 ;
  assign n1292 = n1288 & n1290 ;
  assign n4527 = ~n1292 ;
  assign n1293 = n1291 & n4527 ;
  assign n1294 = n1272 & n1293 ;
  assign n1295 = n1272 | n1293 ;
  assign n4528 = ~n1294 ;
  assign n1296 = n4528 & n1295 ;
  assign n4529 = ~n837 ;
  assign n1297 = n4529 & n871 ;
  assign n4530 = ~n1297 ;
  assign n1298 = n870 & n4530 ;
  assign n1299 = n1296 & n1298 ;
  assign n1300 = n1296 | n1298 ;
  assign n4531 = ~n1299 ;
  assign n1301 = n4531 & n1300 ;
  assign n1302 = n1270 & n1301 ;
  assign n1303 = n1270 | n1301 ;
  assign n4532 = ~n1302 ;
  assign n1304 = n4532 & n1303 ;
  assign n4533 = ~n815 ;
  assign n1305 = n4533 & n901 ;
  assign n4534 = ~n1305 ;
  assign n1306 = n899 & n4534 ;
  assign n1307 = n787 & n806 ;
  assign n1308 = n809 & n812 ;
  assign n1309 = n1307 | n1308 ;
  assign n1310 = n1306 | n1309 ;
  assign n1311 = n1306 & n1309 ;
  assign n4535 = ~n1311 ;
  assign n1312 = n1310 & n4535 ;
  assign n4536 = ~n1304 ;
  assign n1313 = n4536 & n1312 ;
  assign n4537 = ~n1312 ;
  assign n1314 = n1304 & n4537 ;
  assign n1315 = n1313 | n1314 ;
  assign n1316 = n946 & n954 ;
  assign n1317 = n904 & n962 ;
  assign n1318 = n1316 | n1317 ;
  assign n1319 = n1315 | n1318 ;
  assign n1320 = n1315 & n1318 ;
  assign n4538 = ~n1320 ;
  assign n1321 = n1319 & n4538 ;
  assign n4539 = ~n1233 ;
  assign n1322 = n4539 & n1321 ;
  assign n4540 = ~n1321 ;
  assign n1323 = n1233 & n4540 ;
  assign n78 = n1322 | n1323 ;
  assign n4541 = ~n1322 ;
  assign n1325 = n1319 & n4541 ;
  assign n1326 = n1292 | n1294 ;
  assign n4542 = ~n1326 ;
  assign n1327 = n1276 & n4542 ;
  assign n1328 = n4521 & n1326 ;
  assign n1329 = n1327 | n1328 ;
  assign n1330 = n1299 | n1302 ;
  assign n1331 = n1329 | n1330 ;
  assign n1332 = n1329 & n1330 ;
  assign n4543 = ~n1332 ;
  assign n1333 = n1331 & n4543 ;
  assign n1334 = n1251 & n1260 ;
  assign n1335 = n1259 | n1334 ;
  assign n4544 = ~n1241 ;
  assign n1336 = n1239 & n4544 ;
  assign n4545 = ~n1249 ;
  assign n1337 = n1247 & n4545 ;
  assign n1338 = n1336 & n1337 ;
  assign n1339 = n1336 | n1337 ;
  assign n4546 = ~n1338 ;
  assign n1340 = n4546 & n1339 ;
  assign n580 = x6 & x40 ;
  assign n149 = x7 & x39 ;
  assign n150 = x8 & x38 ;
  assign n581 = n149 & n150 ;
  assign n1341 = n149 | n150 ;
  assign n4547 = ~n581 ;
  assign n1342 = n4547 & n1341 ;
  assign n4548 = ~n580 ;
  assign n1343 = n4548 & n1342 ;
  assign n4549 = ~n1342 ;
  assign n1344 = n580 & n4549 ;
  assign n1345 = n1343 | n1344 ;
  assign n4550 = ~n1345 ;
  assign n1346 = n1340 & n4550 ;
  assign n4551 = ~n1340 ;
  assign n1347 = n4551 & n1345 ;
  assign n1348 = n1346 | n1347 ;
  assign n151 = x13 & x33 ;
  assign n152 = x14 & x32 ;
  assign n153 = x11 & x35 ;
  assign n582 = n152 & n153 ;
  assign n1349 = n152 | n153 ;
  assign n4552 = ~n582 ;
  assign n1350 = n4552 & n1349 ;
  assign n1351 = n151 & n1350 ;
  assign n1352 = n151 | n1350 ;
  assign n4553 = ~n1351 ;
  assign n1353 = n4553 & n1352 ;
  assign n4554 = ~n1255 ;
  assign n1354 = n1253 & n4554 ;
  assign n583 = x10 & x36 ;
  assign n154 = x9 & x37 ;
  assign n155 = x12 & x34 ;
  assign n584 = n154 & n155 ;
  assign n1355 = n154 | n155 ;
  assign n4555 = ~n584 ;
  assign n1356 = n4555 & n1355 ;
  assign n4556 = ~n583 ;
  assign n1357 = n4556 & n1356 ;
  assign n4557 = ~n1356 ;
  assign n1358 = n583 & n4557 ;
  assign n1359 = n1357 | n1358 ;
  assign n1360 = n1354 | n1359 ;
  assign n1361 = n1354 & n1359 ;
  assign n4558 = ~n1361 ;
  assign n1362 = n1360 & n4558 ;
  assign n1363 = n1353 & n1362 ;
  assign n1364 = n1353 | n1362 ;
  assign n4559 = ~n1363 ;
  assign n1365 = n4559 & n1364 ;
  assign n1366 = n1348 & n1365 ;
  assign n1367 = n1348 | n1365 ;
  assign n4560 = ~n1366 ;
  assign n1368 = n4560 & n1367 ;
  assign n4561 = ~n1335 ;
  assign n1369 = n4561 & n1368 ;
  assign n4562 = ~n1368 ;
  assign n1370 = n1335 & n4562 ;
  assign n1371 = n1369 | n1370 ;
  assign n1372 = n1274 & n1285 ;
  assign n1373 = n1283 | n1372 ;
  assign n1374 = n4448 & n1279 ;
  assign n4563 = ~n1374 ;
  assign n1375 = n1278 & n4563 ;
  assign n156 = x2 & x44 ;
  assign n157 = x0 & x46 ;
  assign n585 = n156 & n157 ;
  assign n1376 = n156 | n157 ;
  assign n4564 = ~n585 ;
  assign n1377 = n4564 & n1376 ;
  assign n4565 = ~n578 ;
  assign n1378 = n4565 & n1377 ;
  assign n4566 = ~n1377 ;
  assign n1379 = n578 & n4566 ;
  assign n1380 = n1378 | n1379 ;
  assign n586 = x3 & x43 ;
  assign n158 = x4 & x42 ;
  assign n159 = x5 & x41 ;
  assign n587 = n158 & n159 ;
  assign n1381 = n158 | n159 ;
  assign n4567 = ~n587 ;
  assign n1382 = n4567 & n1381 ;
  assign n4568 = ~n586 ;
  assign n1383 = n4568 & n1382 ;
  assign n4569 = ~n1382 ;
  assign n1384 = n586 & n4569 ;
  assign n1385 = n1383 | n1384 ;
  assign n1386 = n1380 | n1385 ;
  assign n1387 = n1380 & n1385 ;
  assign n4570 = ~n1387 ;
  assign n1388 = n1386 & n4570 ;
  assign n4571 = ~n1375 ;
  assign n1389 = n4571 & n1388 ;
  assign n4572 = ~n1388 ;
  assign n1390 = n1375 & n4572 ;
  assign n1391 = n1389 | n1390 ;
  assign n1392 = n1238 & n1243 ;
  assign n1393 = n1236 | n1392 ;
  assign n1394 = n1391 | n1393 ;
  assign n1395 = n1391 & n1393 ;
  assign n4573 = ~n1395 ;
  assign n1396 = n1394 & n4573 ;
  assign n4574 = ~n1373 ;
  assign n1397 = n4574 & n1396 ;
  assign n4575 = ~n1396 ;
  assign n1398 = n1373 & n4575 ;
  assign n1399 = n1397 | n1398 ;
  assign n4576 = ~n1268 ;
  assign n1400 = n1265 & n4576 ;
  assign n1401 = n1399 & n1400 ;
  assign n1402 = n1399 | n1400 ;
  assign n4577 = ~n1401 ;
  assign n1403 = n4577 & n1402 ;
  assign n1404 = n1371 & n1403 ;
  assign n1406 = n1371 | n1403 ;
  assign n4578 = ~n1404 ;
  assign n1407 = n4578 & n1406 ;
  assign n4579 = ~n1407 ;
  assign n1408 = n1333 & n4579 ;
  assign n4580 = ~n1333 ;
  assign n1409 = n4580 & n1407 ;
  assign n1410 = n1408 | n1409 ;
  assign n4581 = ~n1313 ;
  assign n1411 = n1310 & n4581 ;
  assign n1412 = n1410 & n1411 ;
  assign n1413 = n1410 | n1411 ;
  assign n4582 = ~n1412 ;
  assign n1414 = n4582 & n1413 ;
  assign n1415 = n1325 & n1414 ;
  assign n1416 = n1325 | n1414 ;
  assign n4583 = ~n1415 ;
  assign n79 = n4583 & n1416 ;
  assign n1418 = n1412 | n1415 ;
  assign n4584 = ~n1371 ;
  assign n1405 = n4584 & n1403 ;
  assign n4585 = ~n1405 ;
  assign n1419 = n1402 & n4585 ;
  assign n1420 = n1373 & n1396 ;
  assign n1421 = n1395 | n1420 ;
  assign n160 = x0 & x47 ;
  assign n4586 = ~n1378 ;
  assign n1422 = n1376 & n4586 ;
  assign n1423 = n160 & n1422 ;
  assign n1424 = n160 | n1422 ;
  assign n4587 = ~n1423 ;
  assign n1425 = n4587 & n1424 ;
  assign n1426 = n1421 & n1425 ;
  assign n1427 = n1421 | n1425 ;
  assign n4588 = ~n1426 ;
  assign n1428 = n4588 & n1427 ;
  assign n1429 = n1419 & n1428 ;
  assign n1430 = n1419 | n1428 ;
  assign n4589 = ~n1429 ;
  assign n1431 = n4589 & n1430 ;
  assign n588 = x15 & x32 ;
  assign n161 = x14 & x33 ;
  assign n162 = x12 & x35 ;
  assign n589 = n161 & n162 ;
  assign n1432 = n161 | n162 ;
  assign n4590 = ~n589 ;
  assign n1433 = n4590 & n1432 ;
  assign n4591 = ~n588 ;
  assign n1434 = n4591 & n1433 ;
  assign n4592 = ~n1433 ;
  assign n1435 = n588 & n4592 ;
  assign n1436 = n1434 | n1435 ;
  assign n4593 = ~n151 ;
  assign n1437 = n4593 & n1350 ;
  assign n4594 = ~n1437 ;
  assign n1438 = n1349 & n4594 ;
  assign n165 = x13 & x34 ;
  assign n163 = x10 & x37 ;
  assign n164 = x11 & x36 ;
  assign n590 = n163 & n164 ;
  assign n1439 = n163 | n164 ;
  assign n4595 = ~n590 ;
  assign n1440 = n4595 & n1439 ;
  assign n1441 = n165 & n1440 ;
  assign n1442 = n165 | n1440 ;
  assign n4596 = ~n1441 ;
  assign n1443 = n4596 & n1442 ;
  assign n1444 = n1438 | n1443 ;
  assign n1445 = n1438 & n1443 ;
  assign n4597 = ~n1445 ;
  assign n1446 = n1444 & n4597 ;
  assign n4598 = ~n1436 ;
  assign n1447 = n4598 & n1446 ;
  assign n4599 = ~n1446 ;
  assign n1448 = n1436 & n4599 ;
  assign n1449 = n1447 | n1448 ;
  assign n4600 = ~n1357 ;
  assign n1450 = n1355 & n4600 ;
  assign n4601 = ~n1343 ;
  assign n1451 = n1341 & n4601 ;
  assign n168 = x7 & x40 ;
  assign n166 = x8 & x39 ;
  assign n167 = x9 & x38 ;
  assign n591 = n166 & n167 ;
  assign n1452 = n166 | n167 ;
  assign n4602 = ~n591 ;
  assign n1453 = n4602 & n1452 ;
  assign n4603 = ~n1453 ;
  assign n1454 = n168 & n4603 ;
  assign n4604 = ~n168 ;
  assign n1455 = n4604 & n1453 ;
  assign n1456 = n1454 | n1455 ;
  assign n1457 = n1451 | n1456 ;
  assign n1458 = n1451 & n1456 ;
  assign n4605 = ~n1458 ;
  assign n1459 = n1457 & n4605 ;
  assign n4606 = ~n1450 ;
  assign n1460 = n4606 & n1459 ;
  assign n4607 = ~n1459 ;
  assign n1461 = n1450 & n4607 ;
  assign n1462 = n1460 | n1461 ;
  assign n1463 = n1361 | n1363 ;
  assign n1464 = n1462 | n1463 ;
  assign n1465 = n1462 & n1463 ;
  assign n4608 = ~n1465 ;
  assign n1466 = n1464 & n4608 ;
  assign n4609 = ~n1449 ;
  assign n1467 = n4609 & n1466 ;
  assign n4610 = ~n1466 ;
  assign n1468 = n1449 & n4610 ;
  assign n1469 = n1467 | n1468 ;
  assign n169 = x1 & x46 ;
  assign n170 = x3 & x44 ;
  assign n171 = x2 & x45 ;
  assign n592 = n170 & n171 ;
  assign n1470 = n170 | n171 ;
  assign n4611 = ~n592 ;
  assign n1471 = n4611 & n1470 ;
  assign n1472 = n169 & n1471 ;
  assign n1473 = n169 | n1471 ;
  assign n4612 = ~n1472 ;
  assign n1474 = n4612 & n1473 ;
  assign n4613 = ~n1383 ;
  assign n1475 = n1381 & n4613 ;
  assign n174 = x4 & x43 ;
  assign n172 = x5 & x42 ;
  assign n173 = x6 & x41 ;
  assign n593 = n172 & n173 ;
  assign n1476 = n172 | n173 ;
  assign n4614 = ~n593 ;
  assign n1477 = n4614 & n1476 ;
  assign n4615 = ~n1477 ;
  assign n1478 = n174 & n4615 ;
  assign n4616 = ~n174 ;
  assign n1479 = n4616 & n1477 ;
  assign n1480 = n1478 | n1479 ;
  assign n1481 = n1475 | n1480 ;
  assign n1482 = n1475 & n1480 ;
  assign n4617 = ~n1482 ;
  assign n1483 = n1481 & n4617 ;
  assign n4618 = ~n1474 ;
  assign n1484 = n4618 & n1483 ;
  assign n4619 = ~n1483 ;
  assign n1485 = n1474 & n4619 ;
  assign n1486 = n1484 | n1485 ;
  assign n1487 = n1375 & n1388 ;
  assign n1488 = n1387 | n1487 ;
  assign n1489 = n1340 & n1345 ;
  assign n1490 = n1338 | n1489 ;
  assign n1491 = n1488 | n1490 ;
  assign n1492 = n1488 & n1490 ;
  assign n4620 = ~n1492 ;
  assign n1493 = n1491 & n4620 ;
  assign n4621 = ~n1486 ;
  assign n1494 = n4621 & n1493 ;
  assign n4622 = ~n1493 ;
  assign n1495 = n1486 & n4622 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = n1335 & n1368 ;
  assign n1498 = n1366 | n1497 ;
  assign n1499 = n1496 | n1498 ;
  assign n1500 = n1496 & n1498 ;
  assign n4623 = ~n1500 ;
  assign n1501 = n1499 & n4623 ;
  assign n4624 = ~n1469 ;
  assign n1502 = n4624 & n1501 ;
  assign n4625 = ~n1501 ;
  assign n1503 = n1469 & n4625 ;
  assign n1504 = n1502 | n1503 ;
  assign n4626 = ~n1504 ;
  assign n1505 = n1431 & n4626 ;
  assign n4627 = ~n1431 ;
  assign n1506 = n4627 & n1504 ;
  assign n1507 = n1505 | n1506 ;
  assign n1509 = n1333 & n1407 ;
  assign n1508 = n1276 & n1326 ;
  assign n1510 = n1332 | n1508 ;
  assign n4628 = ~n1509 ;
  assign n1511 = n4628 & n1510 ;
  assign n4629 = ~n1508 ;
  assign n1512 = n4629 & n1509 ;
  assign n1513 = n1511 | n1512 ;
  assign n4630 = ~n1507 ;
  assign n1514 = n4630 & n1513 ;
  assign n4631 = ~n1513 ;
  assign n1515 = n1507 & n4631 ;
  assign n1516 = n1514 | n1515 ;
  assign n1517 = n1418 | n1516 ;
  assign n1518 = n1418 & n1516 ;
  assign n4632 = ~n1518 ;
  assign n80 = n1517 & n4632 ;
  assign n1520 = n1431 & n1504 ;
  assign n4633 = ~n1447 ;
  assign n1521 = n1444 & n4633 ;
  assign n4634 = ~n1455 ;
  assign n1522 = n1452 & n4634 ;
  assign n4635 = ~n165 ;
  assign n1523 = n4635 & n1440 ;
  assign n4636 = ~n1523 ;
  assign n1524 = n1439 & n4636 ;
  assign n177 = x8 & x40 ;
  assign n175 = x9 & x39 ;
  assign n176 = x10 & x38 ;
  assign n594 = n175 & n176 ;
  assign n1525 = n175 | n176 ;
  assign n4637 = ~n594 ;
  assign n1526 = n4637 & n1525 ;
  assign n4638 = ~n1526 ;
  assign n1527 = n177 & n4638 ;
  assign n4639 = ~n177 ;
  assign n1528 = n4639 & n1526 ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = n1524 | n1529 ;
  assign n1531 = n1524 & n1529 ;
  assign n4640 = ~n1531 ;
  assign n1532 = n1530 & n4640 ;
  assign n1533 = n1522 & n1532 ;
  assign n1534 = n1522 | n1532 ;
  assign n4641 = ~n1533 ;
  assign n1535 = n4641 & n1534 ;
  assign n4642 = ~n1434 ;
  assign n1536 = n1432 & n4642 ;
  assign n178 = x14 & x34 ;
  assign n179 = x11 & x37 ;
  assign n180 = x12 & x36 ;
  assign n595 = n179 & n180 ;
  assign n1537 = n179 | n180 ;
  assign n4643 = ~n595 ;
  assign n1538 = n4643 & n1537 ;
  assign n1539 = n178 & n1538 ;
  assign n1540 = n178 | n1538 ;
  assign n4644 = ~n1539 ;
  assign n1541 = n4644 & n1540 ;
  assign n596 = x13 & x35 ;
  assign n181 = x15 & x33 ;
  assign n182 = x16 & x32 ;
  assign n597 = n181 & n182 ;
  assign n1542 = n181 | n182 ;
  assign n4645 = ~n597 ;
  assign n1543 = n4645 & n1542 ;
  assign n4646 = ~n596 ;
  assign n1544 = n4646 & n1543 ;
  assign n4647 = ~n1543 ;
  assign n1545 = n596 & n4647 ;
  assign n1546 = n1544 | n1545 ;
  assign n1547 = n1541 | n1546 ;
  assign n1548 = n1541 & n1546 ;
  assign n4648 = ~n1548 ;
  assign n1549 = n1547 & n4648 ;
  assign n1550 = n1536 & n1549 ;
  assign n1551 = n1536 | n1549 ;
  assign n4649 = ~n1550 ;
  assign n1552 = n4649 & n1551 ;
  assign n1553 = n1535 & n1552 ;
  assign n1554 = n1535 | n1552 ;
  assign n4650 = ~n1553 ;
  assign n1555 = n4650 & n1554 ;
  assign n4651 = ~n1521 ;
  assign n1556 = n4651 & n1555 ;
  assign n4652 = ~n1555 ;
  assign n1557 = n1521 & n4652 ;
  assign n1558 = n1556 | n1557 ;
  assign n1559 = n1474 & n1483 ;
  assign n1560 = n1482 | n1559 ;
  assign n4653 = ~n1479 ;
  assign n1561 = n1476 & n4653 ;
  assign n183 = x5 & x43 ;
  assign n184 = x6 & x42 ;
  assign n185 = x7 & x41 ;
  assign n598 = n184 & n185 ;
  assign n1562 = n184 | n185 ;
  assign n4654 = ~n598 ;
  assign n1563 = n4654 & n1562 ;
  assign n1564 = n183 & n1563 ;
  assign n1566 = n183 | n1563 ;
  assign n4655 = ~n1564 ;
  assign n1567 = n4655 & n1566 ;
  assign n188 = x4 & x44 ;
  assign n186 = x2 & x46 ;
  assign n187 = x3 & x45 ;
  assign n599 = n186 & n187 ;
  assign n1568 = n186 | n187 ;
  assign n4656 = ~n599 ;
  assign n1569 = n4656 & n1568 ;
  assign n4657 = ~n1569 ;
  assign n1570 = n188 & n4657 ;
  assign n4658 = ~n188 ;
  assign n1571 = n4658 & n1569 ;
  assign n1572 = n1570 | n1571 ;
  assign n1573 = n1567 | n1572 ;
  assign n1574 = n1567 & n1572 ;
  assign n4659 = ~n1574 ;
  assign n1575 = n1573 & n4659 ;
  assign n4660 = ~n1561 ;
  assign n1576 = n4660 & n1575 ;
  assign n4661 = ~n1575 ;
  assign n1577 = n1561 & n4661 ;
  assign n1578 = n1576 | n1577 ;
  assign n1579 = n1450 & n1459 ;
  assign n1580 = n1458 | n1579 ;
  assign n1581 = n1578 | n1580 ;
  assign n1582 = n1578 & n1580 ;
  assign n4662 = ~n1582 ;
  assign n1583 = n1581 & n4662 ;
  assign n4663 = ~n1560 ;
  assign n1584 = n4663 & n1583 ;
  assign n4664 = ~n1583 ;
  assign n1585 = n1560 & n4664 ;
  assign n1586 = n1584 | n1585 ;
  assign n1587 = n1449 & n1466 ;
  assign n1588 = n1465 | n1587 ;
  assign n1589 = n1586 | n1588 ;
  assign n1590 = n1586 & n1588 ;
  assign n4665 = ~n1590 ;
  assign n1591 = n1589 & n4665 ;
  assign n1592 = n1558 & n1591 ;
  assign n1593 = n1558 | n1591 ;
  assign n4666 = ~n1592 ;
  assign n1594 = n4666 & n1593 ;
  assign n4667 = ~n169 ;
  assign n1595 = n4667 & n1471 ;
  assign n4668 = ~n1595 ;
  assign n1596 = n1470 & n4668 ;
  assign n189 = x1 & x48 ;
  assign n602 = n160 & n189 ;
  assign n600 = x1 & x47 ;
  assign n601 = x0 & x48 ;
  assign n1597 = n600 | n601 ;
  assign n4669 = ~n602 ;
  assign n1598 = n4669 & n1597 ;
  assign n4670 = ~n1596 ;
  assign n1599 = n4670 & n1598 ;
  assign n4671 = ~n1598 ;
  assign n1600 = n1596 & n4671 ;
  assign n1601 = n1599 | n1600 ;
  assign n1602 = n1423 & n1601 ;
  assign n1603 = n1423 | n1601 ;
  assign n4672 = ~n1602 ;
  assign n1604 = n4672 & n1603 ;
  assign n4673 = ~n1494 ;
  assign n1605 = n1491 & n4673 ;
  assign n1606 = n1604 & n1605 ;
  assign n1607 = n1604 | n1605 ;
  assign n4674 = ~n1606 ;
  assign n1608 = n4674 & n1607 ;
  assign n4675 = ~n1502 ;
  assign n1609 = n1499 & n4675 ;
  assign n1610 = n1608 & n1609 ;
  assign n1611 = n1608 | n1609 ;
  assign n4676 = ~n1610 ;
  assign n1612 = n4676 & n1611 ;
  assign n4677 = ~n1594 ;
  assign n1613 = n4677 & n1612 ;
  assign n4678 = ~n1612 ;
  assign n1614 = n1594 & n4678 ;
  assign n1615 = n1613 | n1614 ;
  assign n1616 = n1426 | n1429 ;
  assign n1617 = n1615 | n1616 ;
  assign n1618 = n1615 & n1616 ;
  assign n4679 = ~n1618 ;
  assign n1619 = n1617 & n4679 ;
  assign n1620 = n1520 & n1619 ;
  assign n1621 = n1520 | n1619 ;
  assign n4680 = ~n1620 ;
  assign n1622 = n4680 & n1621 ;
  assign n1623 = n1509 | n1510 ;
  assign n4681 = ~n1514 ;
  assign n1624 = n4681 & n1623 ;
  assign n1625 = n1622 & n1624 ;
  assign n1626 = n1622 | n1624 ;
  assign n4682 = ~n1625 ;
  assign n1627 = n4682 & n1626 ;
  assign n1628 = n1518 & n1627 ;
  assign n1629 = n1518 | n1627 ;
  assign n4683 = ~n1628 ;
  assign n81 = n4683 & n1629 ;
  assign n1631 = n4632 & n1627 ;
  assign n4684 = ~n1631 ;
  assign n1632 = n1626 & n4684 ;
  assign n4685 = ~n1520 ;
  assign n1633 = n4685 & n1619 ;
  assign n4686 = ~n1633 ;
  assign n1634 = n1617 & n4686 ;
  assign n190 = x3 & x46 ;
  assign n191 = x5 & x44 ;
  assign n192 = x4 & x45 ;
  assign n603 = n191 & n192 ;
  assign n1635 = n191 | n192 ;
  assign n4687 = ~n603 ;
  assign n1636 = n4687 & n1635 ;
  assign n1637 = n190 & n1636 ;
  assign n1639 = n190 | n1636 ;
  assign n4688 = ~n1637 ;
  assign n1640 = n4688 & n1639 ;
  assign n4689 = ~n183 ;
  assign n1565 = n4689 & n1563 ;
  assign n4690 = ~n1565 ;
  assign n1641 = n1562 & n4690 ;
  assign n195 = x6 & x43 ;
  assign n193 = x7 & x42 ;
  assign n194 = x8 & x41 ;
  assign n604 = n193 & n194 ;
  assign n1642 = n193 | n194 ;
  assign n4691 = ~n604 ;
  assign n1643 = n4691 & n1642 ;
  assign n1644 = n195 & n1643 ;
  assign n1645 = n195 | n1643 ;
  assign n4692 = ~n1644 ;
  assign n1646 = n4692 & n1645 ;
  assign n4693 = ~n1646 ;
  assign n1647 = n1641 & n4693 ;
  assign n4694 = ~n1641 ;
  assign n1648 = n4694 & n1646 ;
  assign n1649 = n1647 | n1648 ;
  assign n4695 = ~n1640 ;
  assign n1650 = n4695 & n1649 ;
  assign n4696 = ~n1649 ;
  assign n1651 = n1640 & n4696 ;
  assign n1652 = n1650 | n1651 ;
  assign n1653 = n1561 & n1575 ;
  assign n1654 = n1574 | n1653 ;
  assign n1655 = n1531 | n1533 ;
  assign n1656 = n1654 | n1655 ;
  assign n1657 = n1654 & n1655 ;
  assign n4697 = ~n1657 ;
  assign n1658 = n1656 & n4697 ;
  assign n4698 = ~n1652 ;
  assign n1659 = n4698 & n1658 ;
  assign n4699 = ~n1658 ;
  assign n1660 = n1652 & n4699 ;
  assign n1661 = n1659 | n1660 ;
  assign n196 = x14 & x35 ;
  assign n197 = x16 & x33 ;
  assign n198 = x17 & x32 ;
  assign n605 = n197 & n198 ;
  assign n1662 = n197 | n198 ;
  assign n4700 = ~n605 ;
  assign n1663 = n4700 & n1662 ;
  assign n1664 = n196 & n1663 ;
  assign n1665 = n196 | n1663 ;
  assign n4701 = ~n1664 ;
  assign n1666 = n4701 & n1665 ;
  assign n4702 = ~n1544 ;
  assign n1667 = n1542 & n4702 ;
  assign n199 = x12 & x37 ;
  assign n200 = x13 & x36 ;
  assign n201 = x15 & x34 ;
  assign n606 = n200 & n201 ;
  assign n1668 = n200 | n201 ;
  assign n4703 = ~n606 ;
  assign n1669 = n4703 & n1668 ;
  assign n1670 = n199 & n1669 ;
  assign n1672 = n199 | n1669 ;
  assign n4704 = ~n1670 ;
  assign n1673 = n4704 & n1672 ;
  assign n1674 = n1667 | n1673 ;
  assign n1675 = n1667 & n1673 ;
  assign n4705 = ~n1675 ;
  assign n1676 = n1674 & n4705 ;
  assign n1677 = n1666 & n1676 ;
  assign n1678 = n1666 | n1676 ;
  assign n4706 = ~n1677 ;
  assign n1679 = n4706 & n1678 ;
  assign n4707 = ~n178 ;
  assign n1680 = n4707 & n1538 ;
  assign n4708 = ~n1680 ;
  assign n1681 = n1537 & n4708 ;
  assign n4709 = ~n1528 ;
  assign n1682 = n1525 & n4709 ;
  assign n204 = x9 & x40 ;
  assign n202 = x10 & x39 ;
  assign n203 = x11 & x38 ;
  assign n607 = n202 & n203 ;
  assign n1683 = n202 | n203 ;
  assign n4710 = ~n607 ;
  assign n1684 = n4710 & n1683 ;
  assign n4711 = ~n1684 ;
  assign n1685 = n204 & n4711 ;
  assign n4712 = ~n204 ;
  assign n1686 = n4712 & n1684 ;
  assign n1687 = n1685 | n1686 ;
  assign n1688 = n1682 | n1687 ;
  assign n1689 = n1682 & n1687 ;
  assign n4713 = ~n1689 ;
  assign n1690 = n1688 & n4713 ;
  assign n4714 = ~n1681 ;
  assign n1691 = n4714 & n1690 ;
  assign n4715 = ~n1690 ;
  assign n1692 = n1681 & n4715 ;
  assign n1693 = n1691 | n1692 ;
  assign n1694 = n1548 | n1550 ;
  assign n1695 = n1693 | n1694 ;
  assign n1696 = n1693 & n1694 ;
  assign n4716 = ~n1696 ;
  assign n1697 = n1695 & n4716 ;
  assign n1698 = n1679 & n1697 ;
  assign n1699 = n1679 | n1697 ;
  assign n4717 = ~n1698 ;
  assign n1700 = n4717 & n1699 ;
  assign n4718 = ~n1556 ;
  assign n1701 = n1554 & n4718 ;
  assign n1702 = n1700 & n1701 ;
  assign n1703 = n1700 | n1701 ;
  assign n4719 = ~n1702 ;
  assign n1704 = n4719 & n1703 ;
  assign n1705 = n1661 & n1704 ;
  assign n1706 = n1661 | n1704 ;
  assign n4720 = ~n1705 ;
  assign n1707 = n4720 & n1706 ;
  assign n4721 = ~n1584 ;
  assign n1708 = n1581 & n4721 ;
  assign n1709 = n1596 & n1598 ;
  assign n1710 = n602 | n1709 ;
  assign n4722 = ~n1571 ;
  assign n1711 = n1568 & n4722 ;
  assign n608 = x0 & x49 ;
  assign n609 = x2 & x47 ;
  assign n1712 = n608 | n609 ;
  assign n610 = x2 & x49 ;
  assign n1713 = n160 & n610 ;
  assign n4723 = ~n1713 ;
  assign n1714 = n1712 & n4723 ;
  assign n1715 = n189 & n1714 ;
  assign n1716 = n189 | n1714 ;
  assign n4724 = ~n1715 ;
  assign n1717 = n4724 & n1716 ;
  assign n1718 = n1711 | n1717 ;
  assign n1719 = n1711 & n1717 ;
  assign n4725 = ~n1719 ;
  assign n1721 = n1718 & n4725 ;
  assign n1723 = n1710 & n1721 ;
  assign n1724 = n1710 | n1721 ;
  assign n4726 = ~n1723 ;
  assign n1725 = n4726 & n1724 ;
  assign n1726 = n1602 & n1725 ;
  assign n1727 = n1602 | n1725 ;
  assign n4727 = ~n1726 ;
  assign n1728 = n4727 & n1727 ;
  assign n1729 = n1708 & n1728 ;
  assign n1730 = n1708 | n1728 ;
  assign n4728 = ~n1729 ;
  assign n1731 = n4728 & n1730 ;
  assign n1732 = n1590 | n1592 ;
  assign n1733 = n1731 | n1732 ;
  assign n1734 = n1731 & n1732 ;
  assign n4729 = ~n1734 ;
  assign n1735 = n1733 & n4729 ;
  assign n4730 = ~n1707 ;
  assign n1736 = n4730 & n1735 ;
  assign n4731 = ~n1735 ;
  assign n1737 = n1707 & n4731 ;
  assign n1738 = n1736 | n1737 ;
  assign n4732 = ~n1613 ;
  assign n1739 = n1611 & n4732 ;
  assign n1740 = n1606 & n1739 ;
  assign n1741 = n1606 | n1739 ;
  assign n4733 = ~n1740 ;
  assign n1742 = n4733 & n1741 ;
  assign n4734 = ~n1738 ;
  assign n1743 = n4734 & n1742 ;
  assign n4735 = ~n1742 ;
  assign n1744 = n1738 & n4735 ;
  assign n1745 = n1743 | n1744 ;
  assign n4736 = ~n1634 ;
  assign n1746 = n4736 & n1745 ;
  assign n4737 = ~n1745 ;
  assign n1747 = n1634 & n4737 ;
  assign n1748 = n1746 | n1747 ;
  assign n1749 = n1632 | n1748 ;
  assign n1750 = n1632 & n1748 ;
  assign n4738 = ~n1750 ;
  assign n82 = n1749 & n4738 ;
  assign n1752 = n1634 | n1745 ;
  assign n4739 = ~n1632 ;
  assign n1753 = n4739 & n1748 ;
  assign n4740 = ~n1753 ;
  assign n1754 = n1752 & n4740 ;
  assign n4741 = ~n195 ;
  assign n1755 = n4741 & n1643 ;
  assign n4742 = ~n1755 ;
  assign n1756 = n1642 & n4742 ;
  assign n205 = x4 & x46 ;
  assign n206 = x5 & x45 ;
  assign n207 = x6 & x44 ;
  assign n611 = n206 & n207 ;
  assign n1757 = n206 | n207 ;
  assign n4743 = ~n611 ;
  assign n1758 = n4743 & n1757 ;
  assign n1759 = n205 & n1758 ;
  assign n1760 = n205 | n1758 ;
  assign n4744 = ~n1759 ;
  assign n1761 = n4744 & n1760 ;
  assign n210 = x9 & x41 ;
  assign n208 = x8 & x42 ;
  assign n209 = x7 & x43 ;
  assign n612 = n208 & n209 ;
  assign n1762 = n208 | n209 ;
  assign n4745 = ~n612 ;
  assign n1763 = n4745 & n1762 ;
  assign n4746 = ~n1763 ;
  assign n1764 = n210 & n4746 ;
  assign n4747 = ~n210 ;
  assign n1765 = n4747 & n1763 ;
  assign n1766 = n1764 | n1765 ;
  assign n1767 = n1761 | n1766 ;
  assign n1768 = n1761 & n1766 ;
  assign n4748 = ~n1768 ;
  assign n1769 = n1767 & n4748 ;
  assign n1770 = n1756 & n1769 ;
  assign n1771 = n1756 | n1769 ;
  assign n4749 = ~n1770 ;
  assign n1772 = n4749 & n1771 ;
  assign n1773 = n1641 | n1646 ;
  assign n4750 = ~n1650 ;
  assign n1774 = n4750 & n1773 ;
  assign n1775 = n1681 & n1690 ;
  assign n1776 = n1689 | n1775 ;
  assign n4751 = ~n1776 ;
  assign n1777 = n1774 & n4751 ;
  assign n4752 = ~n1774 ;
  assign n1778 = n4752 & n1776 ;
  assign n1779 = n1777 | n1778 ;
  assign n1780 = n1772 & n1779 ;
  assign n1782 = n1772 | n1779 ;
  assign n4753 = ~n1780 ;
  assign n1783 = n4753 & n1782 ;
  assign n211 = x17 & x33 ;
  assign n212 = x18 & x32 ;
  assign n213 = x15 & x35 ;
  assign n613 = n212 & n213 ;
  assign n1784 = n212 | n213 ;
  assign n4754 = ~n613 ;
  assign n1785 = n4754 & n1784 ;
  assign n1786 = n211 & n1785 ;
  assign n1787 = n211 | n1785 ;
  assign n4755 = ~n1786 ;
  assign n1788 = n4755 & n1787 ;
  assign n4756 = ~n196 ;
  assign n1789 = n4756 & n1663 ;
  assign n4757 = ~n1789 ;
  assign n1790 = n1662 & n4757 ;
  assign n216 = x13 & x37 ;
  assign n214 = x14 & x36 ;
  assign n215 = x16 & x34 ;
  assign n614 = n214 & n215 ;
  assign n1791 = n214 | n215 ;
  assign n4758 = ~n614 ;
  assign n1792 = n4758 & n1791 ;
  assign n1793 = n216 & n1792 ;
  assign n1794 = n216 | n1792 ;
  assign n4759 = ~n1793 ;
  assign n1795 = n4759 & n1794 ;
  assign n4760 = ~n1795 ;
  assign n1796 = n1790 & n4760 ;
  assign n4761 = ~n1790 ;
  assign n1797 = n4761 & n1795 ;
  assign n1798 = n1796 | n1797 ;
  assign n1799 = n1788 & n1798 ;
  assign n1800 = n1788 | n1798 ;
  assign n4762 = ~n1799 ;
  assign n1801 = n4762 & n1800 ;
  assign n4763 = ~n199 ;
  assign n1671 = n4763 & n1669 ;
  assign n4764 = ~n1671 ;
  assign n1802 = n1668 & n4764 ;
  assign n4765 = ~n1686 ;
  assign n1803 = n1683 & n4765 ;
  assign n219 = x10 & x40 ;
  assign n217 = x11 & x39 ;
  assign n218 = x12 & x38 ;
  assign n615 = n217 & n218 ;
  assign n1804 = n217 | n218 ;
  assign n4766 = ~n615 ;
  assign n1805 = n4766 & n1804 ;
  assign n4767 = ~n1805 ;
  assign n1806 = n219 & n4767 ;
  assign n4768 = ~n219 ;
  assign n1807 = n4768 & n1805 ;
  assign n1808 = n1806 | n1807 ;
  assign n1809 = n1803 | n1808 ;
  assign n1810 = n1803 & n1808 ;
  assign n4769 = ~n1810 ;
  assign n1811 = n1809 & n4769 ;
  assign n1812 = n1802 & n1811 ;
  assign n1813 = n1802 | n1811 ;
  assign n4770 = ~n1812 ;
  assign n1814 = n4770 & n1813 ;
  assign n4771 = ~n1666 ;
  assign n1815 = n4771 & n1676 ;
  assign n4772 = ~n1815 ;
  assign n1816 = n1674 & n4772 ;
  assign n1817 = n1814 & n1816 ;
  assign n1818 = n1814 | n1816 ;
  assign n4773 = ~n1817 ;
  assign n1819 = n4773 & n1818 ;
  assign n4774 = ~n1801 ;
  assign n1820 = n4774 & n1819 ;
  assign n4775 = ~n1819 ;
  assign n1821 = n1801 & n4775 ;
  assign n1822 = n1820 | n1821 ;
  assign n1823 = n1696 | n1698 ;
  assign n4776 = ~n1823 ;
  assign n1824 = n1822 & n4776 ;
  assign n4777 = ~n1822 ;
  assign n1825 = n4777 & n1823 ;
  assign n1826 = n1824 | n1825 ;
  assign n4778 = ~n1783 ;
  assign n1827 = n4778 & n1826 ;
  assign n4779 = ~n1826 ;
  assign n1829 = n1783 & n4779 ;
  assign n1830 = n1827 | n1829 ;
  assign n4780 = ~n1661 ;
  assign n1831 = n4780 & n1704 ;
  assign n4781 = ~n1831 ;
  assign n1832 = n1703 & n4781 ;
  assign n1833 = n1713 | n1715 ;
  assign n4782 = ~n190 ;
  assign n1638 = n4782 & n1636 ;
  assign n4783 = ~n1638 ;
  assign n1834 = n1635 & n4783 ;
  assign n4784 = ~n1833 ;
  assign n1835 = n4784 & n1834 ;
  assign n4785 = ~n1834 ;
  assign n1836 = n1833 & n4785 ;
  assign n1837 = n1835 | n1836 ;
  assign n222 = x1 & x49 ;
  assign n220 = x2 & x48 ;
  assign n221 = x3 & x47 ;
  assign n616 = n220 & n221 ;
  assign n1838 = n220 | n221 ;
  assign n4786 = ~n616 ;
  assign n1839 = n4786 & n1838 ;
  assign n1840 = n222 & n1839 ;
  assign n1841 = n222 | n1839 ;
  assign n4787 = ~n1840 ;
  assign n1842 = n4787 & n1841 ;
  assign n4788 = ~n1842 ;
  assign n1843 = n1837 & n4788 ;
  assign n4789 = ~n1837 ;
  assign n1844 = n4789 & n1842 ;
  assign n1845 = n1843 | n1844 ;
  assign n223 = x0 & x50 ;
  assign n1720 = n602 | n1719 ;
  assign n1846 = n1718 & n1720 ;
  assign n1847 = n223 & n1846 ;
  assign n1848 = n223 | n1846 ;
  assign n4790 = ~n1847 ;
  assign n1849 = n4790 & n1848 ;
  assign n1850 = n1845 & n1849 ;
  assign n1852 = n1845 | n1849 ;
  assign n4791 = ~n1850 ;
  assign n1853 = n4791 & n1852 ;
  assign n1722 = n1709 & n1721 ;
  assign n1854 = n1652 & n1658 ;
  assign n1855 = n1657 | n1854 ;
  assign n1856 = n1722 & n1855 ;
  assign n1857 = n1722 | n1855 ;
  assign n4792 = ~n1856 ;
  assign n1858 = n4792 & n1857 ;
  assign n4793 = ~n1853 ;
  assign n1859 = n4793 & n1858 ;
  assign n4794 = ~n1858 ;
  assign n1860 = n1853 & n4794 ;
  assign n1861 = n1859 | n1860 ;
  assign n1862 = n1832 | n1861 ;
  assign n1863 = n1832 & n1861 ;
  assign n4795 = ~n1863 ;
  assign n1864 = n1862 & n4795 ;
  assign n1865 = n1830 & n1864 ;
  assign n1866 = n1830 | n1864 ;
  assign n4796 = ~n1865 ;
  assign n1867 = n4796 & n1866 ;
  assign n1868 = n1707 & n1735 ;
  assign n1869 = n1734 | n1868 ;
  assign n1870 = n1726 | n1729 ;
  assign n1871 = n1869 | n1870 ;
  assign n1872 = n1869 & n1870 ;
  assign n4797 = ~n1872 ;
  assign n1873 = n1871 & n4797 ;
  assign n1874 = n1867 & n1873 ;
  assign n1875 = n1867 | n1873 ;
  assign n4798 = ~n1874 ;
  assign n1876 = n4798 & n1875 ;
  assign n4799 = ~n1743 ;
  assign n1877 = n1741 & n4799 ;
  assign n1878 = n1876 & n1877 ;
  assign n1879 = n1876 | n1877 ;
  assign n4800 = ~n1878 ;
  assign n1880 = n4800 & n1879 ;
  assign n1881 = n1754 & n1880 ;
  assign n1882 = n1754 | n1880 ;
  assign n4801 = ~n1881 ;
  assign n83 = n4801 & n1882 ;
  assign n4802 = ~n1754 ;
  assign n1884 = n4802 & n1880 ;
  assign n4803 = ~n1884 ;
  assign n1885 = n1879 & n4803 ;
  assign n4804 = ~n1772 ;
  assign n1781 = n4804 & n1779 ;
  assign n1886 = n1774 | n1776 ;
  assign n4805 = ~n1781 ;
  assign n1887 = n4805 & n1886 ;
  assign n1888 = n1833 & n1834 ;
  assign n1889 = n1837 & n1842 ;
  assign n1890 = n1888 | n1889 ;
  assign n4806 = ~n222 ;
  assign n1891 = n4806 & n1839 ;
  assign n4807 = ~n1891 ;
  assign n1892 = n1838 & n4807 ;
  assign n4808 = ~n205 ;
  assign n1893 = n4808 & n1758 ;
  assign n4809 = ~n1893 ;
  assign n1894 = n1757 & n4809 ;
  assign n224 = x3 & x48 ;
  assign n225 = x4 & x47 ;
  assign n617 = n224 & n225 ;
  assign n1895 = n224 | n225 ;
  assign n4810 = ~n617 ;
  assign n1896 = n4810 & n1895 ;
  assign n4811 = ~n610 ;
  assign n1897 = n4811 & n1896 ;
  assign n4812 = ~n1896 ;
  assign n1898 = n610 & n4812 ;
  assign n1899 = n1897 | n1898 ;
  assign n1900 = n1894 | n1899 ;
  assign n1901 = n1894 & n1899 ;
  assign n4813 = ~n1901 ;
  assign n1902 = n1900 & n4813 ;
  assign n1903 = n1892 & n1902 ;
  assign n1904 = n1892 | n1902 ;
  assign n4814 = ~n1903 ;
  assign n1905 = n4814 & n1904 ;
  assign n226 = x0 & x51 ;
  assign n227 = x1 & x50 ;
  assign n618 = n226 & n227 ;
  assign n1906 = n226 | n227 ;
  assign n4815 = ~n618 ;
  assign n1907 = n4815 & n1906 ;
  assign n1908 = n1905 & n1907 ;
  assign n1909 = n1905 | n1907 ;
  assign n4816 = ~n1908 ;
  assign n1910 = n4816 & n1909 ;
  assign n1911 = n1890 & n1910 ;
  assign n1912 = n1890 | n1910 ;
  assign n4817 = ~n1911 ;
  assign n1913 = n4817 & n1912 ;
  assign n4818 = ~n1845 ;
  assign n1851 = n4818 & n1849 ;
  assign n4819 = ~n1851 ;
  assign n1914 = n1848 & n4819 ;
  assign n1915 = n1913 & n1914 ;
  assign n1916 = n1913 | n1914 ;
  assign n4820 = ~n1915 ;
  assign n1917 = n4820 & n1916 ;
  assign n1918 = n1887 & n1917 ;
  assign n1919 = n1887 | n1917 ;
  assign n4821 = ~n1918 ;
  assign n1920 = n4821 & n1919 ;
  assign n228 = x8 & x43 ;
  assign n229 = x10 & x41 ;
  assign n230 = x9 & x42 ;
  assign n619 = n229 & n230 ;
  assign n1921 = n229 | n230 ;
  assign n4822 = ~n619 ;
  assign n1922 = n4822 & n1921 ;
  assign n1923 = n228 & n1922 ;
  assign n1925 = n228 | n1922 ;
  assign n4823 = ~n1923 ;
  assign n1926 = n4823 & n1925 ;
  assign n4824 = ~n1765 ;
  assign n1927 = n1762 & n4824 ;
  assign n233 = x5 & x46 ;
  assign n231 = x6 & x45 ;
  assign n232 = x7 & x44 ;
  assign n620 = n231 & n232 ;
  assign n1928 = n231 | n232 ;
  assign n4825 = ~n620 ;
  assign n1929 = n4825 & n1928 ;
  assign n1930 = n233 & n1929 ;
  assign n1931 = n233 | n1929 ;
  assign n4826 = ~n1930 ;
  assign n1932 = n4826 & n1931 ;
  assign n4827 = ~n1932 ;
  assign n1933 = n1927 & n4827 ;
  assign n4828 = ~n1927 ;
  assign n1934 = n4828 & n1932 ;
  assign n1935 = n1933 | n1934 ;
  assign n4829 = ~n1926 ;
  assign n1936 = n4829 & n1935 ;
  assign n4830 = ~n1935 ;
  assign n1937 = n1926 & n4830 ;
  assign n1938 = n1936 | n1937 ;
  assign n1939 = n1768 | n1770 ;
  assign n1940 = n1810 | n1812 ;
  assign n1941 = n1939 | n1940 ;
  assign n1942 = n1939 & n1940 ;
  assign n4831 = ~n1942 ;
  assign n1943 = n1941 & n4831 ;
  assign n4832 = ~n1938 ;
  assign n1944 = n4832 & n1943 ;
  assign n4833 = ~n1943 ;
  assign n1945 = n1938 & n4833 ;
  assign n1946 = n1944 | n1945 ;
  assign n1947 = n1790 | n1795 ;
  assign n4834 = ~n1788 ;
  assign n1948 = n4834 & n1798 ;
  assign n4835 = ~n1948 ;
  assign n1949 = n1947 & n4835 ;
  assign n4836 = ~n1807 ;
  assign n1950 = n1804 & n4836 ;
  assign n4837 = ~n216 ;
  assign n1951 = n4837 & n1792 ;
  assign n4838 = ~n1951 ;
  assign n1952 = n1791 & n4838 ;
  assign n4839 = ~n1950 ;
  assign n1953 = n4839 & n1952 ;
  assign n4840 = ~n1952 ;
  assign n1954 = n1950 & n4840 ;
  assign n1955 = n1953 | n1954 ;
  assign n621 = x12 & x39 ;
  assign n234 = x11 & x40 ;
  assign n235 = x13 & x38 ;
  assign n622 = n234 & n235 ;
  assign n1956 = n234 | n235 ;
  assign n4841 = ~n622 ;
  assign n1957 = n4841 & n1956 ;
  assign n4842 = ~n621 ;
  assign n1958 = n4842 & n1957 ;
  assign n4843 = ~n1957 ;
  assign n1959 = n621 & n4843 ;
  assign n1960 = n1958 | n1959 ;
  assign n1961 = n1955 | n1960 ;
  assign n1962 = n1955 & n1960 ;
  assign n4844 = ~n1962 ;
  assign n1963 = n1961 & n4844 ;
  assign n4845 = ~n211 ;
  assign n1964 = n4845 & n1785 ;
  assign n4846 = ~n1964 ;
  assign n1965 = n1784 & n4846 ;
  assign n236 = x15 & x36 ;
  assign n237 = x17 & x34 ;
  assign n238 = x14 & x37 ;
  assign n623 = n237 & n238 ;
  assign n1966 = n237 | n238 ;
  assign n4847 = ~n623 ;
  assign n1967 = n4847 & n1966 ;
  assign n1968 = n236 & n1967 ;
  assign n1969 = n236 | n1967 ;
  assign n4848 = ~n1968 ;
  assign n1970 = n4848 & n1969 ;
  assign n241 = x19 & x32 ;
  assign n239 = x16 & x35 ;
  assign n240 = x18 & x33 ;
  assign n624 = n239 & n240 ;
  assign n1971 = n239 | n240 ;
  assign n4849 = ~n624 ;
  assign n1972 = n4849 & n1971 ;
  assign n4850 = ~n1972 ;
  assign n1973 = n241 & n4850 ;
  assign n4851 = ~n241 ;
  assign n1974 = n4851 & n1972 ;
  assign n1975 = n1973 | n1974 ;
  assign n1976 = n1970 | n1975 ;
  assign n1977 = n1970 & n1975 ;
  assign n4852 = ~n1977 ;
  assign n1978 = n1976 & n4852 ;
  assign n1979 = n1965 & n1978 ;
  assign n1980 = n1965 | n1978 ;
  assign n4853 = ~n1979 ;
  assign n1981 = n4853 & n1980 ;
  assign n1982 = n1963 & n1981 ;
  assign n1983 = n1963 | n1981 ;
  assign n4854 = ~n1982 ;
  assign n1984 = n4854 & n1983 ;
  assign n4855 = ~n1949 ;
  assign n1985 = n4855 & n1984 ;
  assign n4856 = ~n1984 ;
  assign n1986 = n1949 & n4856 ;
  assign n1987 = n1985 | n1986 ;
  assign n1988 = n1801 & n1819 ;
  assign n1989 = n1817 | n1988 ;
  assign n1990 = n1987 | n1989 ;
  assign n1991 = n1987 & n1989 ;
  assign n4857 = ~n1991 ;
  assign n1992 = n1990 & n4857 ;
  assign n4858 = ~n1946 ;
  assign n1993 = n4858 & n1992 ;
  assign n4859 = ~n1992 ;
  assign n1994 = n1946 & n4859 ;
  assign n1995 = n1993 | n1994 ;
  assign n1828 = n1783 & n1826 ;
  assign n1996 = n1822 & n1823 ;
  assign n1997 = n1828 | n1996 ;
  assign n1998 = n1995 | n1997 ;
  assign n1999 = n1995 & n1997 ;
  assign n4860 = ~n1999 ;
  assign n2000 = n1998 & n4860 ;
  assign n2001 = n1920 & n2000 ;
  assign n2002 = n1920 | n2000 ;
  assign n4861 = ~n2001 ;
  assign n2003 = n4861 & n2002 ;
  assign n2004 = n1863 | n1865 ;
  assign n4862 = ~n1859 ;
  assign n2005 = n1857 & n4862 ;
  assign n2006 = n2004 & n2005 ;
  assign n2007 = n2004 | n2005 ;
  assign n4863 = ~n2006 ;
  assign n2008 = n4863 & n2007 ;
  assign n4864 = ~n2003 ;
  assign n2009 = n4864 & n2008 ;
  assign n4865 = ~n2008 ;
  assign n2010 = n2003 & n4865 ;
  assign n2011 = n2009 | n2010 ;
  assign n2012 = n1872 | n1874 ;
  assign n4866 = ~n2012 ;
  assign n2013 = n2011 & n4866 ;
  assign n4867 = ~n2011 ;
  assign n2014 = n4867 & n2012 ;
  assign n2015 = n2013 | n2014 ;
  assign n2016 = n1885 | n2015 ;
  assign n2017 = n1885 & n2015 ;
  assign n4868 = ~n2017 ;
  assign n84 = n2016 & n4868 ;
  assign n2019 = n2011 | n2012 ;
  assign n4869 = ~n1885 ;
  assign n2020 = n4869 & n2015 ;
  assign n4870 = ~n2020 ;
  assign n2021 = n2019 & n4870 ;
  assign n4871 = ~n1920 ;
  assign n2022 = n4871 & n2000 ;
  assign n4872 = ~n2022 ;
  assign n2023 = n1998 & n4872 ;
  assign n242 = x7 & x45 ;
  assign n243 = x8 & x44 ;
  assign n244 = x6 & x46 ;
  assign n625 = n243 & n244 ;
  assign n2024 = n243 | n244 ;
  assign n4873 = ~n625 ;
  assign n2025 = n4873 & n2024 ;
  assign n2026 = n242 & n2025 ;
  assign n2027 = n242 | n2025 ;
  assign n4874 = ~n2026 ;
  assign n2028 = n4874 & n2027 ;
  assign n4875 = ~n228 ;
  assign n1924 = n4875 & n1922 ;
  assign n4876 = ~n1924 ;
  assign n2029 = n1921 & n4876 ;
  assign n247 = x9 & x43 ;
  assign n245 = x10 & x42 ;
  assign n246 = x11 & x41 ;
  assign n626 = n245 & n246 ;
  assign n2030 = n245 | n246 ;
  assign n4877 = ~n626 ;
  assign n2031 = n4877 & n2030 ;
  assign n2032 = n247 & n2031 ;
  assign n2033 = n247 | n2031 ;
  assign n4878 = ~n2032 ;
  assign n2034 = n4878 & n2033 ;
  assign n4879 = ~n2034 ;
  assign n2035 = n2029 & n4879 ;
  assign n4880 = ~n2029 ;
  assign n2036 = n4880 & n2034 ;
  assign n2037 = n2035 | n2036 ;
  assign n2038 = n2028 & n2037 ;
  assign n2039 = n2028 | n2037 ;
  assign n4881 = ~n2038 ;
  assign n2040 = n4881 & n2039 ;
  assign n2041 = n1950 & n1952 ;
  assign n2042 = n1962 | n2041 ;
  assign n2043 = n1927 | n1932 ;
  assign n4882 = ~n1936 ;
  assign n2044 = n4882 & n2043 ;
  assign n2045 = n2042 & n2044 ;
  assign n2046 = n2042 | n2044 ;
  assign n4883 = ~n2045 ;
  assign n2047 = n4883 & n2046 ;
  assign n2048 = n2040 & n2047 ;
  assign n2049 = n2040 | n2047 ;
  assign n4884 = ~n2048 ;
  assign n2050 = n4884 & n2049 ;
  assign n2051 = n1977 | n1979 ;
  assign n4885 = ~n236 ;
  assign n2052 = n4885 & n1967 ;
  assign n4886 = ~n2052 ;
  assign n2053 = n1966 & n4886 ;
  assign n4887 = ~n1958 ;
  assign n2054 = n1956 & n4887 ;
  assign n4888 = ~n2053 ;
  assign n2055 = n4888 & n2054 ;
  assign n4889 = ~n2054 ;
  assign n2056 = n2053 & n4889 ;
  assign n2057 = n2055 | n2056 ;
  assign n250 = x12 & x40 ;
  assign n248 = x13 & x39 ;
  assign n249 = x14 & x38 ;
  assign n627 = n248 & n249 ;
  assign n2058 = n248 | n249 ;
  assign n4890 = ~n627 ;
  assign n2059 = n4890 & n2058 ;
  assign n2060 = n250 & n2059 ;
  assign n2061 = n250 | n2059 ;
  assign n4891 = ~n2060 ;
  assign n2062 = n4891 & n2061 ;
  assign n4892 = ~n2062 ;
  assign n2063 = n2057 & n4892 ;
  assign n4893 = ~n2057 ;
  assign n2064 = n4893 & n2062 ;
  assign n2065 = n2063 | n2064 ;
  assign n4894 = ~n1974 ;
  assign n2066 = n1971 & n4894 ;
  assign n251 = x16 & x36 ;
  assign n252 = x18 & x34 ;
  assign n253 = x15 & x37 ;
  assign n628 = n252 & n253 ;
  assign n2067 = n252 | n253 ;
  assign n4895 = ~n628 ;
  assign n2068 = n4895 & n2067 ;
  assign n2069 = n251 & n2068 ;
  assign n2070 = n251 | n2068 ;
  assign n4896 = ~n2069 ;
  assign n2071 = n4896 & n2070 ;
  assign n256 = x17 & x35 ;
  assign n254 = x19 & x33 ;
  assign n255 = x20 & x32 ;
  assign n629 = n254 & n255 ;
  assign n2072 = n254 | n255 ;
  assign n4897 = ~n629 ;
  assign n2073 = n4897 & n2072 ;
  assign n4898 = ~n2073 ;
  assign n2074 = n256 & n4898 ;
  assign n4899 = ~n256 ;
  assign n2075 = n4899 & n2073 ;
  assign n2076 = n2074 | n2075 ;
  assign n2077 = n2071 | n2076 ;
  assign n2078 = n2071 & n2076 ;
  assign n4900 = ~n2078 ;
  assign n2079 = n2077 & n4900 ;
  assign n2080 = n2066 & n2079 ;
  assign n2081 = n2066 | n2079 ;
  assign n4901 = ~n2080 ;
  assign n2082 = n4901 & n2081 ;
  assign n2083 = n2065 & n2082 ;
  assign n2084 = n2065 | n2082 ;
  assign n4902 = ~n2083 ;
  assign n2085 = n4902 & n2084 ;
  assign n4903 = ~n2051 ;
  assign n2086 = n4903 & n2085 ;
  assign n4904 = ~n2085 ;
  assign n2087 = n2051 & n4904 ;
  assign n2088 = n2086 | n2087 ;
  assign n4905 = ~n1985 ;
  assign n2089 = n1983 & n4905 ;
  assign n2090 = n2088 & n2089 ;
  assign n2091 = n2088 | n2089 ;
  assign n4906 = ~n2090 ;
  assign n2092 = n4906 & n2091 ;
  assign n4907 = ~n2050 ;
  assign n2093 = n4907 & n2092 ;
  assign n4908 = ~n2092 ;
  assign n2094 = n2050 & n4908 ;
  assign n2095 = n2093 | n2094 ;
  assign n2096 = n1938 & n1943 ;
  assign n2097 = n1942 | n2096 ;
  assign n4909 = ~n1897 ;
  assign n2098 = n1895 & n4909 ;
  assign n4910 = ~n233 ;
  assign n2099 = n4910 & n1929 ;
  assign n4911 = ~n2099 ;
  assign n2100 = n1928 & n4911 ;
  assign n630 = x4 & x48 ;
  assign n257 = x3 & x49 ;
  assign n258 = x5 & x47 ;
  assign n631 = n257 & n258 ;
  assign n2101 = n257 | n258 ;
  assign n4912 = ~n631 ;
  assign n2102 = n4912 & n2101 ;
  assign n4913 = ~n630 ;
  assign n2103 = n4913 & n2102 ;
  assign n4914 = ~n2102 ;
  assign n2104 = n630 & n4914 ;
  assign n2105 = n2103 | n2104 ;
  assign n4915 = ~n2105 ;
  assign n2106 = n2100 & n4915 ;
  assign n4916 = ~n2100 ;
  assign n2107 = n4916 & n2105 ;
  assign n2108 = n2106 | n2107 ;
  assign n2109 = n2098 & n2108 ;
  assign n2110 = n2098 | n2108 ;
  assign n4917 = ~n2109 ;
  assign n2111 = n4917 & n2110 ;
  assign n2112 = n1901 | n1903 ;
  assign n4918 = ~n2112 ;
  assign n2113 = n2111 & n4918 ;
  assign n4919 = ~n2111 ;
  assign n2114 = n4919 & n2112 ;
  assign n2115 = n2113 | n2114 ;
  assign n261 = x1 & x51 ;
  assign n259 = x0 & x52 ;
  assign n260 = x2 & x50 ;
  assign n2116 = n259 | n260 ;
  assign n2117 = n261 & n2116 ;
  assign n2118 = n1907 & n2117 ;
  assign n262 = x2 & x52 ;
  assign n4920 = ~n262 ;
  assign n2119 = n4920 & n2116 ;
  assign n4921 = ~n2119 ;
  assign n2120 = n223 & n4921 ;
  assign n2121 = n261 | n2116 ;
  assign n4922 = ~n2120 ;
  assign n2122 = n4922 & n2121 ;
  assign n4923 = ~n2118 ;
  assign n2123 = n4923 & n2122 ;
  assign n4924 = ~n2115 ;
  assign n2124 = n4924 & n2123 ;
  assign n4925 = ~n2123 ;
  assign n2125 = n2115 & n4925 ;
  assign n2126 = n2124 | n2125 ;
  assign n2127 = n1908 | n1911 ;
  assign n2128 = n2126 | n2127 ;
  assign n2129 = n2126 & n2127 ;
  assign n4926 = ~n2129 ;
  assign n2130 = n2128 & n4926 ;
  assign n4927 = ~n2097 ;
  assign n2131 = n4927 & n2130 ;
  assign n4928 = ~n2130 ;
  assign n2132 = n2097 & n4928 ;
  assign n2133 = n2131 | n2132 ;
  assign n4929 = ~n1993 ;
  assign n2134 = n1990 & n4929 ;
  assign n4930 = ~n2133 ;
  assign n2135 = n4930 & n2134 ;
  assign n4931 = ~n2134 ;
  assign n2136 = n2133 & n4931 ;
  assign n2137 = n2135 | n2136 ;
  assign n4932 = ~n2095 ;
  assign n2138 = n4932 & n2137 ;
  assign n4933 = ~n2137 ;
  assign n2139 = n2095 & n4933 ;
  assign n2140 = n2138 | n2139 ;
  assign n2141 = n1915 | n1918 ;
  assign n2142 = n2140 | n2141 ;
  assign n2143 = n2140 & n2141 ;
  assign n4934 = ~n2143 ;
  assign n2144 = n2142 & n4934 ;
  assign n2145 = n2023 & n2144 ;
  assign n2146 = n2023 | n2144 ;
  assign n4935 = ~n2145 ;
  assign n2147 = n4935 & n2146 ;
  assign n2148 = n2003 & n2008 ;
  assign n2149 = n2006 | n2148 ;
  assign n2150 = n2147 | n2149 ;
  assign n2151 = n2147 & n2149 ;
  assign n4936 = ~n2151 ;
  assign n2152 = n2150 & n4936 ;
  assign n2153 = n2021 & n2152 ;
  assign n2154 = n2021 | n2152 ;
  assign n4937 = ~n2153 ;
  assign n85 = n4937 & n2154 ;
  assign n2156 = n2133 | n2134 ;
  assign n4938 = ~n2138 ;
  assign n2157 = n4938 & n2156 ;
  assign n2158 = n2111 | n2112 ;
  assign n4939 = ~n2125 ;
  assign n2159 = n4939 & n2158 ;
  assign n263 = x2 & x51 ;
  assign n264 = x3 & x50 ;
  assign n265 = x1 & x52 ;
  assign n632 = n264 & n265 ;
  assign n2160 = n264 | n265 ;
  assign n4940 = ~n632 ;
  assign n2161 = n4940 & n2160 ;
  assign n2162 = n263 & n2161 ;
  assign n2164 = n263 | n2161 ;
  assign n4941 = ~n2162 ;
  assign n2165 = n4941 & n2164 ;
  assign n266 = x0 & x53 ;
  assign n633 = n259 & n260 ;
  assign n2166 = n633 | n2117 ;
  assign n4942 = ~n2166 ;
  assign n2167 = n266 & n4942 ;
  assign n4943 = ~n266 ;
  assign n2168 = n4943 & n2166 ;
  assign n2169 = n2167 | n2168 ;
  assign n4944 = ~n2165 ;
  assign n2170 = n4944 & n2169 ;
  assign n4945 = ~n2169 ;
  assign n2172 = n2165 & n4945 ;
  assign n2173 = n2170 | n2172 ;
  assign n4946 = ~n242 ;
  assign n2174 = n4946 & n2025 ;
  assign n4947 = ~n2174 ;
  assign n2175 = n2024 & n4947 ;
  assign n4948 = ~n2103 ;
  assign n2176 = n2101 & n4948 ;
  assign n269 = x4 & x49 ;
  assign n267 = x6 & x47 ;
  assign n268 = x5 & x48 ;
  assign n634 = n267 & n268 ;
  assign n2177 = n267 | n268 ;
  assign n4949 = ~n634 ;
  assign n2178 = n4949 & n2177 ;
  assign n4950 = ~n2178 ;
  assign n2179 = n269 & n4950 ;
  assign n4951 = ~n269 ;
  assign n2180 = n4951 & n2178 ;
  assign n2181 = n2179 | n2180 ;
  assign n4952 = ~n2181 ;
  assign n2182 = n2176 & n4952 ;
  assign n4953 = ~n2176 ;
  assign n2183 = n4953 & n2181 ;
  assign n2184 = n2182 | n2183 ;
  assign n2185 = n2175 & n2184 ;
  assign n2186 = n2175 | n2184 ;
  assign n4954 = ~n2185 ;
  assign n2187 = n4954 & n2186 ;
  assign n2188 = n2100 & n2105 ;
  assign n2189 = n2109 | n2188 ;
  assign n4955 = ~n2189 ;
  assign n2190 = n2187 & n4955 ;
  assign n4956 = ~n2187 ;
  assign n2191 = n4956 & n2189 ;
  assign n2192 = n2190 | n2191 ;
  assign n2193 = n2173 & n2192 ;
  assign n2195 = n2173 | n2192 ;
  assign n4957 = ~n2193 ;
  assign n2196 = n4957 & n2195 ;
  assign n2197 = n2045 | n2048 ;
  assign n2198 = n2196 | n2197 ;
  assign n2199 = n2196 & n2197 ;
  assign n4958 = ~n2199 ;
  assign n2200 = n2198 & n4958 ;
  assign n2201 = n2159 | n2200 ;
  assign n2202 = n2159 & n2200 ;
  assign n4959 = ~n2202 ;
  assign n2203 = n2201 & n4959 ;
  assign n270 = x18 & x35 ;
  assign n271 = x20 & x33 ;
  assign n272 = x21 & x32 ;
  assign n635 = n271 & n272 ;
  assign n2204 = n271 | n272 ;
  assign n4960 = ~n635 ;
  assign n2205 = n4960 & n2204 ;
  assign n2206 = n270 & n2205 ;
  assign n2208 = n270 | n2205 ;
  assign n4961 = ~n2206 ;
  assign n2209 = n4961 & n2208 ;
  assign n4962 = ~n2075 ;
  assign n2210 = n2072 & n4962 ;
  assign n275 = x17 & x36 ;
  assign n273 = x16 & x37 ;
  assign n274 = x19 & x34 ;
  assign n636 = n273 & n274 ;
  assign n2211 = n273 | n274 ;
  assign n4963 = ~n636 ;
  assign n2212 = n4963 & n2211 ;
  assign n2213 = n275 & n2212 ;
  assign n2214 = n275 | n2212 ;
  assign n4964 = ~n2213 ;
  assign n2215 = n4964 & n2214 ;
  assign n2216 = n2210 | n2215 ;
  assign n2217 = n2210 & n2215 ;
  assign n4965 = ~n2217 ;
  assign n2218 = n2216 & n4965 ;
  assign n4966 = ~n2209 ;
  assign n2219 = n4966 & n2218 ;
  assign n4967 = ~n2218 ;
  assign n2220 = n2209 & n4967 ;
  assign n2221 = n2219 | n2220 ;
  assign n4968 = ~n250 ;
  assign n2222 = n4968 & n2059 ;
  assign n4969 = ~n2222 ;
  assign n2223 = n2058 & n4969 ;
  assign n4970 = ~n251 ;
  assign n2224 = n4970 & n2068 ;
  assign n4971 = ~n2224 ;
  assign n2225 = n2067 & n4971 ;
  assign n637 = x13 & x40 ;
  assign n276 = x14 & x39 ;
  assign n277 = x15 & x38 ;
  assign n638 = n276 & n277 ;
  assign n2226 = n276 | n277 ;
  assign n4972 = ~n638 ;
  assign n2227 = n4972 & n2226 ;
  assign n4973 = ~n637 ;
  assign n2228 = n4973 & n2227 ;
  assign n4974 = ~n2227 ;
  assign n2229 = n637 & n4974 ;
  assign n2230 = n2228 | n2229 ;
  assign n2231 = n2225 | n2230 ;
  assign n2232 = n2225 & n2230 ;
  assign n4975 = ~n2232 ;
  assign n2233 = n2231 & n4975 ;
  assign n2234 = n2223 & n2233 ;
  assign n2235 = n2223 | n2233 ;
  assign n4976 = ~n2234 ;
  assign n2236 = n4976 & n2235 ;
  assign n2237 = n2078 | n2080 ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = n2236 & n2237 ;
  assign n4977 = ~n2239 ;
  assign n2240 = n2238 & n4977 ;
  assign n4978 = ~n2221 ;
  assign n2241 = n4978 & n2240 ;
  assign n4979 = ~n2240 ;
  assign n2243 = n2221 & n4979 ;
  assign n2244 = n2241 | n2243 ;
  assign n2245 = n2029 | n2034 ;
  assign n4980 = ~n2028 ;
  assign n2246 = n4980 & n2037 ;
  assign n4981 = ~n2246 ;
  assign n2247 = n2245 & n4981 ;
  assign n278 = x9 & x44 ;
  assign n279 = x8 & x45 ;
  assign n280 = x7 & x46 ;
  assign n639 = n279 & n280 ;
  assign n2248 = n279 | n280 ;
  assign n4982 = ~n639 ;
  assign n2249 = n4982 & n2248 ;
  assign n2250 = n278 & n2249 ;
  assign n2252 = n278 | n2249 ;
  assign n4983 = ~n2250 ;
  assign n2253 = n4983 & n2252 ;
  assign n4984 = ~n247 ;
  assign n2254 = n4984 & n2031 ;
  assign n4985 = ~n2254 ;
  assign n2255 = n2030 & n4985 ;
  assign n283 = x10 & x43 ;
  assign n281 = x11 & x42 ;
  assign n282 = x12 & x41 ;
  assign n640 = n281 & n282 ;
  assign n2256 = n281 | n282 ;
  assign n4986 = ~n640 ;
  assign n2257 = n4986 & n2256 ;
  assign n4987 = ~n2257 ;
  assign n2258 = n283 & n4987 ;
  assign n4988 = ~n283 ;
  assign n2259 = n4988 & n2257 ;
  assign n2260 = n2258 | n2259 ;
  assign n2261 = n2255 | n2260 ;
  assign n2262 = n2255 & n2260 ;
  assign n4989 = ~n2262 ;
  assign n2263 = n2261 & n4989 ;
  assign n4990 = ~n2253 ;
  assign n2264 = n4990 & n2263 ;
  assign n4991 = ~n2263 ;
  assign n2266 = n2253 & n4991 ;
  assign n2267 = n2264 | n2266 ;
  assign n2268 = n2053 & n2054 ;
  assign n2269 = n2057 & n2062 ;
  assign n2270 = n2268 | n2269 ;
  assign n4992 = ~n2270 ;
  assign n2271 = n2267 & n4992 ;
  assign n4993 = ~n2267 ;
  assign n2272 = n4993 & n2270 ;
  assign n2273 = n2271 | n2272 ;
  assign n2274 = n2247 & n2273 ;
  assign n2276 = n2247 | n2273 ;
  assign n4994 = ~n2274 ;
  assign n2277 = n4994 & n2276 ;
  assign n2278 = n2051 & n2085 ;
  assign n2279 = n2083 | n2278 ;
  assign n2280 = n2277 | n2279 ;
  assign n2281 = n2277 & n2279 ;
  assign n4995 = ~n2281 ;
  assign n2282 = n2280 & n4995 ;
  assign n2283 = n2244 & n2282 ;
  assign n2284 = n2244 | n2282 ;
  assign n4996 = ~n2283 ;
  assign n2285 = n4996 & n2284 ;
  assign n4997 = ~n2093 ;
  assign n2286 = n2091 & n4997 ;
  assign n2287 = n2285 & n2286 ;
  assign n2288 = n2285 | n2286 ;
  assign n4998 = ~n2287 ;
  assign n2289 = n4998 & n2288 ;
  assign n4999 = ~n2203 ;
  assign n2290 = n4999 & n2289 ;
  assign n5000 = ~n2289 ;
  assign n2291 = n2203 & n5000 ;
  assign n2292 = n2290 | n2291 ;
  assign n2293 = n261 & n2120 ;
  assign n5001 = ~n2292 ;
  assign n2294 = n5001 & n2293 ;
  assign n5002 = ~n2293 ;
  assign n2295 = n2292 & n5002 ;
  assign n2296 = n2294 | n2295 ;
  assign n5003 = ~n2131 ;
  assign n2297 = n2128 & n5003 ;
  assign n2298 = n2296 & n2297 ;
  assign n2299 = n2296 | n2297 ;
  assign n5004 = ~n2298 ;
  assign n2300 = n5004 & n2299 ;
  assign n2301 = n2157 & n2300 ;
  assign n2302 = n2157 | n2300 ;
  assign n5005 = ~n2301 ;
  assign n2303 = n5005 & n2302 ;
  assign n2304 = n2143 | n2145 ;
  assign n5006 = ~n2304 ;
  assign n2305 = n2303 & n5006 ;
  assign n5007 = ~n2303 ;
  assign n2306 = n5007 & n2304 ;
  assign n2307 = n2305 | n2306 ;
  assign n2308 = n2021 | n2151 ;
  assign n2309 = n2150 & n2308 ;
  assign n2310 = n2307 | n2309 ;
  assign n2311 = n2307 & n2309 ;
  assign n5008 = ~n2311 ;
  assign n86 = n2310 & n5008 ;
  assign n2313 = n2303 & n2304 ;
  assign n2314 = n2311 | n2313 ;
  assign n5009 = ~n2180 ;
  assign n2315 = n2177 & n5009 ;
  assign n5010 = ~n278 ;
  assign n2251 = n5010 & n2249 ;
  assign n5011 = ~n2251 ;
  assign n2316 = n2248 & n5011 ;
  assign n2317 = n2315 & n2316 ;
  assign n2318 = n2315 | n2316 ;
  assign n5012 = ~n2317 ;
  assign n2319 = n5012 & n2318 ;
  assign n284 = x5 & x49 ;
  assign n285 = x6 & x48 ;
  assign n286 = x7 & x47 ;
  assign n641 = n285 & n286 ;
  assign n2320 = n285 | n286 ;
  assign n5013 = ~n641 ;
  assign n2321 = n5013 & n2320 ;
  assign n2322 = n284 & n2321 ;
  assign n2324 = n284 | n2321 ;
  assign n5014 = ~n2322 ;
  assign n2325 = n5014 & n2324 ;
  assign n5015 = ~n2325 ;
  assign n2326 = n2319 & n5015 ;
  assign n5016 = ~n2319 ;
  assign n2327 = n5016 & n2325 ;
  assign n2328 = n2326 | n2327 ;
  assign n5017 = ~n263 ;
  assign n2163 = n5017 & n2161 ;
  assign n5018 = ~n2163 ;
  assign n2329 = n2160 & n5018 ;
  assign n287 = x3 & x51 ;
  assign n288 = x4 & x50 ;
  assign n642 = n287 & n288 ;
  assign n2330 = n287 | n288 ;
  assign n5019 = ~n642 ;
  assign n2331 = n5019 & n2330 ;
  assign n2332 = n262 & n2331 ;
  assign n2334 = n262 | n2331 ;
  assign n5020 = ~n2332 ;
  assign n2335 = n5020 & n2334 ;
  assign n5021 = ~n2335 ;
  assign n2336 = n2329 & n5021 ;
  assign n5022 = ~n2329 ;
  assign n2337 = n5022 & n2335 ;
  assign n2338 = n2336 | n2337 ;
  assign n289 = x0 & x54 ;
  assign n290 = x1 & x53 ;
  assign n643 = n289 & n290 ;
  assign n2339 = n289 | n290 ;
  assign n5023 = ~n643 ;
  assign n2340 = n5023 & n2339 ;
  assign n5024 = ~n2338 ;
  assign n2341 = n5024 & n2340 ;
  assign n5025 = ~n2340 ;
  assign n2342 = n2338 & n5025 ;
  assign n2343 = n2341 | n2342 ;
  assign n2344 = n2176 & n2181 ;
  assign n2345 = n2185 | n2344 ;
  assign n5026 = ~n2345 ;
  assign n2346 = n2343 & n5026 ;
  assign n5027 = ~n2343 ;
  assign n2347 = n5027 & n2345 ;
  assign n2348 = n2346 | n2347 ;
  assign n2349 = n2328 & n2348 ;
  assign n2350 = n2328 | n2348 ;
  assign n5028 = ~n2349 ;
  assign n2351 = n5028 & n2350 ;
  assign n5029 = ~n2173 ;
  assign n2194 = n5029 & n2192 ;
  assign n2352 = n2187 | n2189 ;
  assign n5030 = ~n2194 ;
  assign n2353 = n5030 & n2352 ;
  assign n5031 = ~n2247 ;
  assign n2275 = n5031 & n2273 ;
  assign n2354 = n2267 | n2270 ;
  assign n5032 = ~n2275 ;
  assign n2355 = n5032 & n2354 ;
  assign n2356 = n2353 & n2355 ;
  assign n2357 = n2353 | n2355 ;
  assign n5033 = ~n2356 ;
  assign n2358 = n5033 & n2357 ;
  assign n5034 = ~n2351 ;
  assign n2359 = n5034 & n2358 ;
  assign n5035 = ~n2358 ;
  assign n2360 = n2351 & n5035 ;
  assign n2361 = n2359 | n2360 ;
  assign n291 = x8 & x46 ;
  assign n292 = x10 & x44 ;
  assign n293 = x9 & x45 ;
  assign n644 = n292 & n293 ;
  assign n2362 = n292 | n293 ;
  assign n5036 = ~n644 ;
  assign n2363 = n5036 & n2362 ;
  assign n2364 = n291 & n2363 ;
  assign n2365 = n291 | n2363 ;
  assign n5037 = ~n2364 ;
  assign n2366 = n5037 & n2365 ;
  assign n5038 = ~n2259 ;
  assign n2367 = n2256 & n5038 ;
  assign n294 = x12 & x42 ;
  assign n295 = x11 & x43 ;
  assign n296 = x13 & x41 ;
  assign n645 = n295 & n296 ;
  assign n2368 = n295 | n296 ;
  assign n5039 = ~n645 ;
  assign n2369 = n5039 & n2368 ;
  assign n2370 = n294 & n2369 ;
  assign n2371 = n294 | n2369 ;
  assign n5040 = ~n2370 ;
  assign n2372 = n5040 & n2371 ;
  assign n5041 = ~n2372 ;
  assign n2373 = n2367 & n5041 ;
  assign n5042 = ~n2367 ;
  assign n2374 = n5042 & n2372 ;
  assign n2375 = n2373 | n2374 ;
  assign n2376 = n2366 & n2375 ;
  assign n2377 = n2366 | n2375 ;
  assign n5043 = ~n2376 ;
  assign n2378 = n5043 & n2377 ;
  assign n2265 = n2253 & n2263 ;
  assign n2379 = n2262 | n2265 ;
  assign n2380 = n2232 | n2234 ;
  assign n2381 = n2379 | n2380 ;
  assign n2382 = n2379 & n2380 ;
  assign n5044 = ~n2382 ;
  assign n2383 = n2381 & n5044 ;
  assign n2384 = n2378 & n2383 ;
  assign n2385 = n2378 | n2383 ;
  assign n5045 = ~n2384 ;
  assign n2386 = n5045 & n2385 ;
  assign n5046 = ~n2219 ;
  assign n2387 = n2216 & n5046 ;
  assign n5047 = ~n270 ;
  assign n2207 = n5047 & n2205 ;
  assign n5048 = ~n2207 ;
  assign n2388 = n2204 & n5048 ;
  assign n297 = x19 & x35 ;
  assign n298 = x21 & x33 ;
  assign n299 = x22 & x32 ;
  assign n646 = n298 & n299 ;
  assign n2389 = n298 | n299 ;
  assign n5049 = ~n646 ;
  assign n2390 = n5049 & n2389 ;
  assign n2391 = n297 & n2390 ;
  assign n2392 = n297 | n2390 ;
  assign n5050 = ~n2391 ;
  assign n2393 = n5050 & n2392 ;
  assign n647 = x17 & x37 ;
  assign n300 = x18 & x36 ;
  assign n301 = x20 & x34 ;
  assign n648 = n300 & n301 ;
  assign n2394 = n300 | n301 ;
  assign n5051 = ~n648 ;
  assign n2395 = n5051 & n2394 ;
  assign n5052 = ~n647 ;
  assign n2396 = n5052 & n2395 ;
  assign n5053 = ~n2395 ;
  assign n2397 = n647 & n5053 ;
  assign n2398 = n2396 | n2397 ;
  assign n2399 = n2393 | n2398 ;
  assign n2400 = n2393 & n2398 ;
  assign n5054 = ~n2400 ;
  assign n2401 = n2399 & n5054 ;
  assign n2402 = n2388 & n2401 ;
  assign n2403 = n2388 | n2401 ;
  assign n5055 = ~n2402 ;
  assign n2404 = n5055 & n2403 ;
  assign n5056 = ~n2228 ;
  assign n2405 = n2226 & n5056 ;
  assign n5057 = ~n275 ;
  assign n2406 = n5057 & n2212 ;
  assign n5058 = ~n2406 ;
  assign n2407 = n2211 & n5058 ;
  assign n304 = x14 & x40 ;
  assign n302 = x15 & x39 ;
  assign n303 = x16 & x38 ;
  assign n649 = n302 & n303 ;
  assign n2408 = n302 | n303 ;
  assign n5059 = ~n649 ;
  assign n2409 = n5059 & n2408 ;
  assign n5060 = ~n2409 ;
  assign n2410 = n304 & n5060 ;
  assign n5061 = ~n304 ;
  assign n2411 = n5061 & n2409 ;
  assign n2412 = n2410 | n2411 ;
  assign n5062 = ~n2412 ;
  assign n2413 = n2407 & n5062 ;
  assign n5063 = ~n2407 ;
  assign n2414 = n5063 & n2412 ;
  assign n2415 = n2413 | n2414 ;
  assign n2416 = n2405 & n2415 ;
  assign n2417 = n2405 | n2415 ;
  assign n5064 = ~n2416 ;
  assign n2418 = n5064 & n2417 ;
  assign n2419 = n2404 & n2418 ;
  assign n2420 = n2404 | n2418 ;
  assign n5065 = ~n2419 ;
  assign n2421 = n5065 & n2420 ;
  assign n5066 = ~n2387 ;
  assign n2422 = n5066 & n2421 ;
  assign n5067 = ~n2421 ;
  assign n2423 = n2387 & n5067 ;
  assign n2424 = n2422 | n2423 ;
  assign n2242 = n2221 & n2240 ;
  assign n2425 = n2239 | n2242 ;
  assign n2426 = n2424 | n2425 ;
  assign n2427 = n2424 & n2425 ;
  assign n5068 = ~n2427 ;
  assign n2428 = n2426 & n5068 ;
  assign n5069 = ~n2386 ;
  assign n2429 = n5069 & n2428 ;
  assign n5070 = ~n2428 ;
  assign n2430 = n2386 & n5070 ;
  assign n2431 = n2429 | n2430 ;
  assign n5071 = ~n2244 ;
  assign n2432 = n5071 & n2282 ;
  assign n5072 = ~n2432 ;
  assign n2433 = n2280 & n5072 ;
  assign n5073 = ~n2431 ;
  assign n2434 = n5073 & n2433 ;
  assign n5074 = ~n2433 ;
  assign n2435 = n2431 & n5074 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = n2361 & n2436 ;
  assign n2438 = n2361 | n2436 ;
  assign n5075 = ~n2437 ;
  assign n2439 = n5075 & n2438 ;
  assign n2440 = n2199 | n2202 ;
  assign n2171 = n2165 & n2169 ;
  assign n2441 = n266 & n2166 ;
  assign n2442 = n2171 | n2441 ;
  assign n5076 = ~n2442 ;
  assign n2443 = n2440 & n5076 ;
  assign n5077 = ~n2440 ;
  assign n2444 = n5077 & n2442 ;
  assign n2445 = n2443 | n2444 ;
  assign n5078 = ~n2290 ;
  assign n2446 = n2288 & n5078 ;
  assign n2447 = n2445 & n2446 ;
  assign n2448 = n2445 | n2446 ;
  assign n5079 = ~n2447 ;
  assign n2449 = n5079 & n2448 ;
  assign n2450 = n2439 & n2449 ;
  assign n2451 = n2439 | n2449 ;
  assign n5080 = ~n2450 ;
  assign n2452 = n5080 & n2451 ;
  assign n2453 = n2292 & n2293 ;
  assign n2454 = n2301 & n2453 ;
  assign n2455 = n2301 | n2453 ;
  assign n5081 = ~n2454 ;
  assign n2456 = n5081 & n2455 ;
  assign n2457 = n2298 | n2456 ;
  assign n5082 = ~n2457 ;
  assign n2458 = n2452 & n5082 ;
  assign n5083 = ~n2452 ;
  assign n2459 = n5083 & n2457 ;
  assign n2460 = n2458 | n2459 ;
  assign n5084 = ~n2460 ;
  assign n2461 = n2314 & n5084 ;
  assign n5085 = ~n2314 ;
  assign n2462 = n5085 & n2460 ;
  assign n87 = n2461 | n2462 ;
  assign n2464 = n2314 & n2460 ;
  assign n2465 = n2351 & n2358 ;
  assign n2466 = n2356 | n2465 ;
  assign n2467 = n2338 & n2340 ;
  assign n2468 = n2329 & n2335 ;
  assign n2469 = n5023 & n2468 ;
  assign n5086 = ~n2468 ;
  assign n2470 = n643 & n5086 ;
  assign n2471 = n2469 | n2470 ;
  assign n2472 = n2467 | n2471 ;
  assign n2473 = n2466 | n2472 ;
  assign n2474 = n2466 & n2472 ;
  assign n5087 = ~n2474 ;
  assign n2475 = n2473 & n5087 ;
  assign n2476 = n2387 & n2421 ;
  assign n2477 = n2419 | n2476 ;
  assign n305 = x14 & x41 ;
  assign n306 = x13 & x42 ;
  assign n307 = x12 & x43 ;
  assign n650 = n306 & n307 ;
  assign n2478 = n306 | n307 ;
  assign n5088 = ~n650 ;
  assign n2479 = n5088 & n2478 ;
  assign n2480 = n305 & n2479 ;
  assign n2482 = n305 | n2479 ;
  assign n5089 = ~n2480 ;
  assign n2483 = n5089 & n2482 ;
  assign n5090 = ~n294 ;
  assign n2484 = n5090 & n2369 ;
  assign n5091 = ~n2484 ;
  assign n2485 = n2368 & n5091 ;
  assign n310 = x9 & x46 ;
  assign n308 = x10 & x45 ;
  assign n309 = x11 & x44 ;
  assign n651 = n308 & n309 ;
  assign n2486 = n308 | n309 ;
  assign n5092 = ~n651 ;
  assign n2487 = n5092 & n2486 ;
  assign n2488 = n310 & n2487 ;
  assign n2489 = n310 | n2487 ;
  assign n5093 = ~n2488 ;
  assign n2490 = n5093 & n2489 ;
  assign n5094 = ~n2490 ;
  assign n2491 = n2485 & n5094 ;
  assign n5095 = ~n2485 ;
  assign n2492 = n5095 & n2490 ;
  assign n2493 = n2491 | n2492 ;
  assign n5096 = ~n2483 ;
  assign n2494 = n5096 & n2493 ;
  assign n5097 = ~n2493 ;
  assign n2495 = n2483 & n5097 ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = n2407 & n2412 ;
  assign n2498 = n2416 | n2497 ;
  assign n2499 = n2367 | n2372 ;
  assign n5098 = ~n2366 ;
  assign n2500 = n5098 & n2375 ;
  assign n5099 = ~n2500 ;
  assign n2501 = n2499 & n5099 ;
  assign n5100 = ~n2498 ;
  assign n2502 = n5100 & n2501 ;
  assign n5101 = ~n2501 ;
  assign n2503 = n2498 & n5101 ;
  assign n2504 = n2502 | n2503 ;
  assign n5102 = ~n2496 ;
  assign n2505 = n5102 & n2504 ;
  assign n5103 = ~n2504 ;
  assign n2507 = n2496 & n5103 ;
  assign n2508 = n2505 | n2507 ;
  assign n311 = x20 & x35 ;
  assign n312 = x22 & x33 ;
  assign n313 = x23 & x32 ;
  assign n652 = n312 & n313 ;
  assign n2509 = n312 | n313 ;
  assign n5104 = ~n652 ;
  assign n2510 = n5104 & n2509 ;
  assign n2511 = n311 & n2510 ;
  assign n2513 = n311 | n2510 ;
  assign n5105 = ~n2511 ;
  assign n2514 = n5105 & n2513 ;
  assign n5106 = ~n297 ;
  assign n2515 = n5106 & n2390 ;
  assign n5107 = ~n2515 ;
  assign n2516 = n2389 & n5107 ;
  assign n316 = x19 & x36 ;
  assign n314 = x18 & x37 ;
  assign n315 = x21 & x34 ;
  assign n653 = n314 & n315 ;
  assign n2517 = n314 | n315 ;
  assign n5108 = ~n653 ;
  assign n2518 = n5108 & n2517 ;
  assign n2519 = n316 & n2518 ;
  assign n2520 = n316 | n2518 ;
  assign n5109 = ~n2519 ;
  assign n2521 = n5109 & n2520 ;
  assign n5110 = ~n2521 ;
  assign n2522 = n2516 & n5110 ;
  assign n5111 = ~n2516 ;
  assign n2523 = n5111 & n2521 ;
  assign n2524 = n2522 | n2523 ;
  assign n5112 = ~n2514 ;
  assign n2525 = n5112 & n2524 ;
  assign n5113 = ~n2524 ;
  assign n2526 = n2514 & n5113 ;
  assign n2527 = n2525 | n2526 ;
  assign n5114 = ~n2396 ;
  assign n2528 = n2394 & n5114 ;
  assign n5115 = ~n2411 ;
  assign n2529 = n2408 & n5115 ;
  assign n319 = x15 & x40 ;
  assign n317 = x16 & x39 ;
  assign n318 = x17 & x38 ;
  assign n654 = n317 & n318 ;
  assign n2530 = n317 | n318 ;
  assign n5116 = ~n654 ;
  assign n2531 = n5116 & n2530 ;
  assign n5117 = ~n2531 ;
  assign n2532 = n319 & n5117 ;
  assign n5118 = ~n319 ;
  assign n2533 = n5118 & n2531 ;
  assign n2534 = n2532 | n2533 ;
  assign n5119 = ~n2534 ;
  assign n2535 = n2529 & n5119 ;
  assign n5120 = ~n2529 ;
  assign n2536 = n5120 & n2534 ;
  assign n2537 = n2535 | n2536 ;
  assign n5121 = ~n2528 ;
  assign n2538 = n5121 & n2537 ;
  assign n5122 = ~n2537 ;
  assign n2539 = n2528 & n5122 ;
  assign n2540 = n2538 | n2539 ;
  assign n2541 = n2400 | n2402 ;
  assign n2542 = n2540 | n2541 ;
  assign n2543 = n2540 & n2541 ;
  assign n5123 = ~n2543 ;
  assign n2544 = n2542 & n5123 ;
  assign n5124 = ~n2527 ;
  assign n2545 = n5124 & n2544 ;
  assign n5125 = ~n2544 ;
  assign n2547 = n2527 & n5125 ;
  assign n2548 = n2545 | n2547 ;
  assign n2549 = n2508 & n2548 ;
  assign n2550 = n2508 | n2548 ;
  assign n5126 = ~n2549 ;
  assign n2551 = n5126 & n2550 ;
  assign n5127 = ~n2477 ;
  assign n2552 = n5127 & n2551 ;
  assign n5128 = ~n2551 ;
  assign n2553 = n2477 & n5128 ;
  assign n2554 = n2552 | n2553 ;
  assign n2555 = n2343 | n2345 ;
  assign n5129 = ~n2328 ;
  assign n2556 = n5129 & n2348 ;
  assign n5130 = ~n2556 ;
  assign n2557 = n2555 & n5130 ;
  assign n5131 = ~n291 ;
  assign n2558 = n5131 & n2363 ;
  assign n5132 = ~n2558 ;
  assign n2559 = n2362 & n5132 ;
  assign n5133 = ~n284 ;
  assign n2323 = n5133 & n2321 ;
  assign n5134 = ~n2323 ;
  assign n2560 = n2320 & n5134 ;
  assign n2561 = n2559 & n2560 ;
  assign n2562 = n2559 | n2560 ;
  assign n5135 = ~n2561 ;
  assign n2563 = n5135 & n2562 ;
  assign n320 = x7 & x48 ;
  assign n321 = x6 & x49 ;
  assign n322 = x8 & x47 ;
  assign n655 = n321 & n322 ;
  assign n2564 = n321 | n322 ;
  assign n5136 = ~n655 ;
  assign n2565 = n5136 & n2564 ;
  assign n2566 = n320 & n2565 ;
  assign n2568 = n320 | n2565 ;
  assign n5137 = ~n2566 ;
  assign n2569 = n5137 & n2568 ;
  assign n5138 = ~n2569 ;
  assign n2570 = n2563 & n5138 ;
  assign n5139 = ~n2563 ;
  assign n2571 = n5139 & n2569 ;
  assign n2572 = n2570 | n2571 ;
  assign n2333 = n4920 & n2331 ;
  assign n5140 = ~n2333 ;
  assign n2573 = n2330 & n5140 ;
  assign n323 = x1 & x54 ;
  assign n324 = x2 & x53 ;
  assign n325 = x0 & x55 ;
  assign n656 = n324 & n325 ;
  assign n2574 = n324 | n325 ;
  assign n5141 = ~n656 ;
  assign n2575 = n5141 & n2574 ;
  assign n2576 = n323 & n2575 ;
  assign n2578 = n323 | n2575 ;
  assign n5142 = ~n2576 ;
  assign n2579 = n5142 & n2578 ;
  assign n657 = x3 & x52 ;
  assign n326 = x4 & x51 ;
  assign n327 = x5 & x50 ;
  assign n658 = n326 & n327 ;
  assign n2580 = n326 | n327 ;
  assign n5143 = ~n658 ;
  assign n2581 = n5143 & n2580 ;
  assign n5144 = ~n657 ;
  assign n2582 = n5144 & n2581 ;
  assign n5145 = ~n2581 ;
  assign n2583 = n657 & n5145 ;
  assign n2584 = n2582 | n2583 ;
  assign n2585 = n2579 | n2584 ;
  assign n2586 = n2579 & n2584 ;
  assign n5146 = ~n2586 ;
  assign n2587 = n2585 & n5146 ;
  assign n2588 = n2573 & n2587 ;
  assign n2589 = n2573 | n2587 ;
  assign n5147 = ~n2588 ;
  assign n2590 = n5147 & n2589 ;
  assign n2591 = n2319 & n2325 ;
  assign n2592 = n2317 | n2591 ;
  assign n5148 = ~n2592 ;
  assign n2593 = n2590 & n5148 ;
  assign n5149 = ~n2590 ;
  assign n2594 = n5149 & n2592 ;
  assign n2595 = n2593 | n2594 ;
  assign n2596 = n2572 & n2595 ;
  assign n2598 = n2572 | n2595 ;
  assign n5150 = ~n2596 ;
  assign n2599 = n5150 & n2598 ;
  assign n2600 = n2382 | n2384 ;
  assign n2601 = n2599 | n2600 ;
  assign n2602 = n2599 & n2600 ;
  assign n5151 = ~n2602 ;
  assign n2603 = n2601 & n5151 ;
  assign n2604 = n2557 & n2603 ;
  assign n2605 = n2557 | n2603 ;
  assign n5152 = ~n2604 ;
  assign n2606 = n5152 & n2605 ;
  assign n5153 = ~n2429 ;
  assign n2607 = n2426 & n5153 ;
  assign n2608 = n2606 & n2607 ;
  assign n2609 = n2606 | n2607 ;
  assign n5154 = ~n2608 ;
  assign n2610 = n5154 & n2609 ;
  assign n2611 = n2554 & n2610 ;
  assign n2613 = n2554 | n2610 ;
  assign n5155 = ~n2611 ;
  assign n2614 = n5155 & n2613 ;
  assign n2615 = n2431 & n2433 ;
  assign n2616 = n2437 | n2615 ;
  assign n2617 = n2614 | n2616 ;
  assign n2618 = n2614 & n2616 ;
  assign n5156 = ~n2618 ;
  assign n2619 = n2617 & n5156 ;
  assign n2620 = n2475 & n2619 ;
  assign n2621 = n2475 | n2619 ;
  assign n5157 = ~n2620 ;
  assign n2622 = n5157 & n2621 ;
  assign n2623 = n2440 & n2442 ;
  assign n5158 = ~n2439 ;
  assign n2624 = n5158 & n2449 ;
  assign n5159 = ~n2624 ;
  assign n2625 = n2448 & n5159 ;
  assign n2626 = n2623 & n2625 ;
  assign n2627 = n2623 | n2625 ;
  assign n5160 = ~n2626 ;
  assign n2628 = n5160 & n2627 ;
  assign n2629 = n2622 & n2628 ;
  assign n2630 = n2622 | n2628 ;
  assign n5161 = ~n2629 ;
  assign n2631 = n5161 & n2630 ;
  assign n2632 = n2452 & n2457 ;
  assign n2633 = n2454 | n2632 ;
  assign n5162 = ~n2633 ;
  assign n2634 = n2631 & n5162 ;
  assign n5163 = ~n2631 ;
  assign n2635 = n5163 & n2633 ;
  assign n2636 = n2634 | n2635 ;
  assign n2637 = n2464 | n2636 ;
  assign n2638 = n2464 & n2636 ;
  assign n5164 = ~n2638 ;
  assign n88 = n2637 & n5164 ;
  assign n5165 = ~n2554 ;
  assign n2612 = n5165 & n2610 ;
  assign n5166 = ~n2612 ;
  assign n2640 = n2609 & n5166 ;
  assign n2641 = n2602 | n2604 ;
  assign n2642 = n643 & n2468 ;
  assign n2643 = n2586 | n2588 ;
  assign n328 = x0 & x56 ;
  assign n5167 = ~n323 ;
  assign n2577 = n5167 & n2575 ;
  assign n5168 = ~n2577 ;
  assign n2644 = n2574 & n5168 ;
  assign n2645 = n328 & n2644 ;
  assign n2646 = n328 | n2644 ;
  assign n5169 = ~n2645 ;
  assign n2647 = n5169 & n2646 ;
  assign n2648 = n2643 & n2647 ;
  assign n2649 = n2643 | n2647 ;
  assign n5170 = ~n2648 ;
  assign n2650 = n5170 & n2649 ;
  assign n5171 = ~n2650 ;
  assign n2651 = n2642 & n5171 ;
  assign n5172 = ~n2642 ;
  assign n2652 = n5172 & n2650 ;
  assign n2653 = n2651 | n2652 ;
  assign n5173 = ~n2641 ;
  assign n2654 = n5173 & n2653 ;
  assign n5174 = ~n2653 ;
  assign n2655 = n2641 & n5174 ;
  assign n2656 = n2654 | n2655 ;
  assign n2657 = n2640 & n2656 ;
  assign n2658 = n2640 | n2656 ;
  assign n5175 = ~n2657 ;
  assign n2659 = n5175 & n2658 ;
  assign n5176 = ~n305 ;
  assign n2481 = n5176 & n2479 ;
  assign n5177 = ~n2481 ;
  assign n2660 = n2478 & n5177 ;
  assign n329 = x11 & x45 ;
  assign n330 = x12 & x44 ;
  assign n331 = x10 & x46 ;
  assign n659 = n330 & n331 ;
  assign n2661 = n330 | n331 ;
  assign n5178 = ~n659 ;
  assign n2662 = n5178 & n2661 ;
  assign n2663 = n329 & n2662 ;
  assign n2664 = n329 | n2662 ;
  assign n5179 = ~n2663 ;
  assign n2665 = n5179 & n2664 ;
  assign n660 = x13 & x43 ;
  assign n332 = x14 & x42 ;
  assign n333 = x15 & x41 ;
  assign n661 = n332 & n333 ;
  assign n2666 = n332 | n333 ;
  assign n5180 = ~n661 ;
  assign n2667 = n5180 & n2666 ;
  assign n5181 = ~n660 ;
  assign n2668 = n5181 & n2667 ;
  assign n5182 = ~n2667 ;
  assign n2669 = n660 & n5182 ;
  assign n2670 = n2668 | n2669 ;
  assign n2671 = n2665 | n2670 ;
  assign n2672 = n2665 & n2670 ;
  assign n5183 = ~n2672 ;
  assign n2673 = n2671 & n5183 ;
  assign n2674 = n2660 & n2673 ;
  assign n2675 = n2660 | n2673 ;
  assign n5184 = ~n2674 ;
  assign n2676 = n5184 & n2675 ;
  assign n2677 = n2529 & n2534 ;
  assign n2678 = n2528 & n2537 ;
  assign n2679 = n2677 | n2678 ;
  assign n2680 = n2485 | n2490 ;
  assign n5185 = ~n2494 ;
  assign n2681 = n5185 & n2680 ;
  assign n5186 = ~n2679 ;
  assign n2682 = n5186 & n2681 ;
  assign n5187 = ~n2681 ;
  assign n2683 = n2679 & n5187 ;
  assign n2684 = n2682 | n2683 ;
  assign n2685 = n2676 & n2684 ;
  assign n2687 = n2676 | n2684 ;
  assign n5188 = ~n2685 ;
  assign n2688 = n5188 & n2687 ;
  assign n334 = x23 & x33 ;
  assign n335 = x24 & x32 ;
  assign n336 = x21 & x35 ;
  assign n662 = n335 & n336 ;
  assign n2689 = n335 | n336 ;
  assign n5189 = ~n662 ;
  assign n2690 = n5189 & n2689 ;
  assign n2691 = n334 & n2690 ;
  assign n2692 = n334 | n2690 ;
  assign n5190 = ~n2691 ;
  assign n2693 = n5190 & n2692 ;
  assign n5191 = ~n311 ;
  assign n2512 = n5191 & n2510 ;
  assign n5192 = ~n2512 ;
  assign n2694 = n2509 & n5192 ;
  assign n663 = x20 & x36 ;
  assign n337 = x19 & x37 ;
  assign n338 = x22 & x34 ;
  assign n664 = n337 & n338 ;
  assign n2695 = n337 | n338 ;
  assign n5193 = ~n664 ;
  assign n2696 = n5193 & n2695 ;
  assign n5194 = ~n663 ;
  assign n2697 = n5194 & n2696 ;
  assign n5195 = ~n2696 ;
  assign n2698 = n663 & n5195 ;
  assign n2699 = n2697 | n2698 ;
  assign n5196 = ~n2699 ;
  assign n2700 = n2694 & n5196 ;
  assign n5197 = ~n2694 ;
  assign n2701 = n5197 & n2699 ;
  assign n2702 = n2700 | n2701 ;
  assign n5198 = ~n2693 ;
  assign n2703 = n5198 & n2702 ;
  assign n5199 = ~n2702 ;
  assign n2705 = n2693 & n5199 ;
  assign n2706 = n2703 | n2705 ;
  assign n5200 = ~n2533 ;
  assign n2707 = n2530 & n5200 ;
  assign n5201 = ~n316 ;
  assign n2708 = n5201 & n2518 ;
  assign n5202 = ~n2708 ;
  assign n2709 = n2517 & n5202 ;
  assign n2710 = n2707 & n2709 ;
  assign n2711 = n2707 | n2709 ;
  assign n5203 = ~n2710 ;
  assign n2712 = n5203 & n2711 ;
  assign n341 = x18 & x38 ;
  assign n339 = x17 & x39 ;
  assign n340 = x16 & x40 ;
  assign n665 = n339 & n340 ;
  assign n2713 = n339 | n340 ;
  assign n5204 = ~n665 ;
  assign n2714 = n5204 & n2713 ;
  assign n2715 = n341 & n2714 ;
  assign n2716 = n341 | n2714 ;
  assign n5205 = ~n2715 ;
  assign n2717 = n5205 & n2716 ;
  assign n5206 = ~n2717 ;
  assign n2718 = n2712 & n5206 ;
  assign n5207 = ~n2712 ;
  assign n2719 = n5207 & n2717 ;
  assign n2720 = n2718 | n2719 ;
  assign n2721 = n2516 | n2521 ;
  assign n5208 = ~n2525 ;
  assign n2722 = n5208 & n2721 ;
  assign n2723 = n2720 & n2722 ;
  assign n2724 = n2720 | n2722 ;
  assign n5209 = ~n2723 ;
  assign n2725 = n5209 & n2724 ;
  assign n5210 = ~n2706 ;
  assign n2726 = n5210 & n2725 ;
  assign n5211 = ~n2725 ;
  assign n2727 = n2706 & n5211 ;
  assign n2728 = n2726 | n2727 ;
  assign n2546 = n2527 & n2544 ;
  assign n2729 = n2543 | n2546 ;
  assign n2730 = n2728 | n2729 ;
  assign n2731 = n2728 & n2729 ;
  assign n5212 = ~n2731 ;
  assign n2732 = n2730 & n5212 ;
  assign n5213 = ~n2688 ;
  assign n2733 = n5213 & n2732 ;
  assign n5214 = ~n2732 ;
  assign n2734 = n2688 & n5214 ;
  assign n2735 = n2733 | n2734 ;
  assign n2736 = n2477 & n2551 ;
  assign n2737 = n2549 | n2736 ;
  assign n342 = x5 & x51 ;
  assign n343 = x6 & x50 ;
  assign n344 = x4 & x52 ;
  assign n666 = n343 & n344 ;
  assign n2738 = n343 | n344 ;
  assign n5215 = ~n666 ;
  assign n2739 = n5215 & n2738 ;
  assign n2740 = n342 & n2739 ;
  assign n2741 = n342 | n2739 ;
  assign n5216 = ~n2740 ;
  assign n2742 = n5216 & n2741 ;
  assign n5217 = ~n2582 ;
  assign n2743 = n2580 & n5217 ;
  assign n347 = x3 & x53 ;
  assign n345 = x1 & x55 ;
  assign n346 = x2 & x54 ;
  assign n667 = n345 & n346 ;
  assign n2744 = n345 | n346 ;
  assign n5218 = ~n667 ;
  assign n2745 = n5218 & n2744 ;
  assign n2746 = n347 & n2745 ;
  assign n2747 = n347 | n2745 ;
  assign n5219 = ~n2746 ;
  assign n2748 = n5219 & n2747 ;
  assign n5220 = ~n2748 ;
  assign n2749 = n2743 & n5220 ;
  assign n5221 = ~n2743 ;
  assign n2750 = n5221 & n2748 ;
  assign n2751 = n2749 | n2750 ;
  assign n5222 = ~n2742 ;
  assign n2752 = n5222 & n2751 ;
  assign n5223 = ~n2751 ;
  assign n2753 = n2742 & n5223 ;
  assign n2754 = n2752 | n2753 ;
  assign n5224 = ~n310 ;
  assign n2755 = n5224 & n2487 ;
  assign n5225 = ~n2755 ;
  assign n2756 = n2486 & n5225 ;
  assign n5226 = ~n320 ;
  assign n2567 = n5226 & n2565 ;
  assign n5227 = ~n2567 ;
  assign n2757 = n2564 & n5227 ;
  assign n2758 = n2756 & n2757 ;
  assign n2759 = n2756 | n2757 ;
  assign n5228 = ~n2758 ;
  assign n2760 = n5228 & n2759 ;
  assign n350 = x8 & x48 ;
  assign n348 = x7 & x49 ;
  assign n349 = x9 & x47 ;
  assign n668 = n348 & n349 ;
  assign n2761 = n348 | n349 ;
  assign n5229 = ~n668 ;
  assign n2762 = n5229 & n2761 ;
  assign n2763 = n350 & n2762 ;
  assign n2764 = n350 | n2762 ;
  assign n5230 = ~n2763 ;
  assign n2765 = n5230 & n2764 ;
  assign n5231 = ~n2765 ;
  assign n2766 = n2760 & n5231 ;
  assign n5232 = ~n2760 ;
  assign n2767 = n5232 & n2765 ;
  assign n2768 = n2766 | n2767 ;
  assign n2769 = n2563 & n2569 ;
  assign n2770 = n2561 | n2769 ;
  assign n5233 = ~n2770 ;
  assign n2771 = n2768 & n5233 ;
  assign n5234 = ~n2768 ;
  assign n2772 = n5234 & n2770 ;
  assign n2773 = n2771 | n2772 ;
  assign n5235 = ~n2754 ;
  assign n2774 = n5235 & n2773 ;
  assign n5236 = ~n2773 ;
  assign n2776 = n2754 & n5236 ;
  assign n2777 = n2774 | n2776 ;
  assign n5237 = ~n2572 ;
  assign n2597 = n5237 & n2595 ;
  assign n2778 = n2590 | n2592 ;
  assign n5238 = ~n2597 ;
  assign n2779 = n5238 & n2778 ;
  assign n2506 = n2496 & n2504 ;
  assign n2780 = n2498 & n2501 ;
  assign n2781 = n2506 | n2780 ;
  assign n5239 = ~n2781 ;
  assign n2782 = n2779 & n5239 ;
  assign n5240 = ~n2779 ;
  assign n2783 = n5240 & n2781 ;
  assign n2784 = n2782 | n2783 ;
  assign n2785 = n2777 & n2784 ;
  assign n2787 = n2777 | n2784 ;
  assign n5241 = ~n2785 ;
  assign n2788 = n5241 & n2787 ;
  assign n2789 = n2737 | n2788 ;
  assign n2790 = n2737 & n2788 ;
  assign n5242 = ~n2790 ;
  assign n2791 = n2789 & n5242 ;
  assign n5243 = ~n2735 ;
  assign n2792 = n5243 & n2791 ;
  assign n5244 = ~n2791 ;
  assign n2793 = n2735 & n5244 ;
  assign n2794 = n2792 | n2793 ;
  assign n2795 = n2659 | n2794 ;
  assign n2796 = n2659 & n2794 ;
  assign n5245 = ~n2796 ;
  assign n2797 = n2795 & n5245 ;
  assign n2798 = n2474 & n5156 ;
  assign n5246 = ~n2475 ;
  assign n2799 = n5246 & n2619 ;
  assign n5247 = ~n2799 ;
  assign n2800 = n2617 & n5247 ;
  assign n2801 = n5087 & n2800 ;
  assign n2802 = n2798 | n2801 ;
  assign n2803 = n2797 & n2802 ;
  assign n2805 = n2797 | n2802 ;
  assign n5248 = ~n2803 ;
  assign n2806 = n5248 & n2805 ;
  assign n2807 = n2626 | n2629 ;
  assign n2808 = n2806 | n2807 ;
  assign n2809 = n2806 & n2807 ;
  assign n5249 = ~n2809 ;
  assign n2810 = n2808 & n5249 ;
  assign n2811 = n2631 & n2633 ;
  assign n2812 = n2638 | n2811 ;
  assign n2813 = n2810 & n2812 ;
  assign n2814 = n2810 | n2812 ;
  assign n5250 = ~n2813 ;
  assign n89 = n5250 & n2814 ;
  assign n2816 = n2809 | n2813 ;
  assign n2817 = n2641 | n2653 ;
  assign n5251 = ~n2640 ;
  assign n2818 = n5251 & n2656 ;
  assign n5252 = ~n2818 ;
  assign n2819 = n2817 & n5252 ;
  assign n2775 = n2754 & n2773 ;
  assign n2820 = n2768 & n2770 ;
  assign n2821 = n2775 | n2820 ;
  assign n351 = x6 & x51 ;
  assign n352 = x7 & x50 ;
  assign n353 = x5 & x52 ;
  assign n669 = n352 & n353 ;
  assign n2822 = n352 | n353 ;
  assign n5253 = ~n669 ;
  assign n2823 = n5253 & n2822 ;
  assign n2824 = n351 & n2823 ;
  assign n2826 = n351 | n2823 ;
  assign n5254 = ~n2824 ;
  assign n2827 = n5254 & n2826 ;
  assign n5255 = ~n342 ;
  assign n2828 = n5255 & n2739 ;
  assign n5256 = ~n2828 ;
  assign n2829 = n2738 & n5256 ;
  assign n354 = x2 & x55 ;
  assign n355 = x3 & x54 ;
  assign n356 = x4 & x53 ;
  assign n670 = n355 & n356 ;
  assign n2830 = n355 | n356 ;
  assign n5257 = ~n670 ;
  assign n2831 = n5257 & n2830 ;
  assign n2832 = n354 & n2831 ;
  assign n2834 = n354 | n2831 ;
  assign n5258 = ~n2832 ;
  assign n2835 = n5258 & n2834 ;
  assign n5259 = ~n2835 ;
  assign n2836 = n2829 & n5259 ;
  assign n5260 = ~n2829 ;
  assign n2837 = n5260 & n2835 ;
  assign n2838 = n2836 | n2837 ;
  assign n5261 = ~n2827 ;
  assign n2839 = n5261 & n2838 ;
  assign n5262 = ~n2838 ;
  assign n2840 = n2827 & n5262 ;
  assign n2841 = n2839 | n2840 ;
  assign n5263 = ~n350 ;
  assign n2842 = n5263 & n2762 ;
  assign n5264 = ~n2842 ;
  assign n2843 = n2761 & n5264 ;
  assign n5265 = ~n329 ;
  assign n2844 = n5265 & n2662 ;
  assign n5266 = ~n2844 ;
  assign n2845 = n2661 & n5266 ;
  assign n671 = x8 & x49 ;
  assign n357 = x9 & x48 ;
  assign n358 = x10 & x47 ;
  assign n672 = n357 & n358 ;
  assign n2846 = n357 | n358 ;
  assign n5267 = ~n672 ;
  assign n2847 = n5267 & n2846 ;
  assign n5268 = ~n671 ;
  assign n2848 = n5268 & n2847 ;
  assign n5269 = ~n2847 ;
  assign n2849 = n671 & n5269 ;
  assign n2850 = n2848 | n2849 ;
  assign n2851 = n2845 | n2850 ;
  assign n2852 = n2845 & n2850 ;
  assign n5270 = ~n2852 ;
  assign n2853 = n2851 & n5270 ;
  assign n2854 = n2843 & n2853 ;
  assign n2855 = n2843 | n2853 ;
  assign n5271 = ~n2854 ;
  assign n2856 = n5271 & n2855 ;
  assign n2857 = n2760 & n2765 ;
  assign n2858 = n2758 | n2857 ;
  assign n5272 = ~n2858 ;
  assign n2859 = n2856 & n5272 ;
  assign n5273 = ~n2856 ;
  assign n2860 = n5273 & n2858 ;
  assign n2861 = n2859 | n2860 ;
  assign n5274 = ~n2841 ;
  assign n2862 = n5274 & n2861 ;
  assign n5275 = ~n2861 ;
  assign n2864 = n2841 & n5275 ;
  assign n2865 = n2862 | n2864 ;
  assign n5276 = ~n2676 ;
  assign n2686 = n5276 & n2684 ;
  assign n2866 = n2679 | n2681 ;
  assign n5277 = ~n2686 ;
  assign n2867 = n5277 & n2866 ;
  assign n2868 = n2865 & n2867 ;
  assign n2869 = n2865 | n2867 ;
  assign n5278 = ~n2868 ;
  assign n2870 = n5278 & n2869 ;
  assign n5279 = ~n2821 ;
  assign n2871 = n5279 & n2870 ;
  assign n5280 = ~n2870 ;
  assign n2872 = n2821 & n5280 ;
  assign n2873 = n2871 | n2872 ;
  assign n359 = x24 & x33 ;
  assign n360 = x25 & x32 ;
  assign n361 = x22 & x35 ;
  assign n673 = n360 & n361 ;
  assign n2874 = n360 | n361 ;
  assign n5281 = ~n673 ;
  assign n2875 = n5281 & n2874 ;
  assign n2876 = n359 & n2875 ;
  assign n2877 = n359 | n2875 ;
  assign n5282 = ~n2876 ;
  assign n2878 = n5282 & n2877 ;
  assign n5283 = ~n334 ;
  assign n2879 = n5283 & n2690 ;
  assign n5284 = ~n2879 ;
  assign n2880 = n2689 & n5284 ;
  assign n364 = x21 & x36 ;
  assign n362 = x20 & x37 ;
  assign n363 = x23 & x34 ;
  assign n674 = n362 & n363 ;
  assign n2881 = n362 | n363 ;
  assign n5285 = ~n674 ;
  assign n2882 = n5285 & n2881 ;
  assign n2883 = n364 & n2882 ;
  assign n2884 = n364 | n2882 ;
  assign n5286 = ~n2883 ;
  assign n2885 = n5286 & n2884 ;
  assign n5287 = ~n2885 ;
  assign n2886 = n2880 & n5287 ;
  assign n5288 = ~n2880 ;
  assign n2887 = n5288 & n2885 ;
  assign n2888 = n2886 | n2887 ;
  assign n5289 = ~n2878 ;
  assign n2889 = n5289 & n2888 ;
  assign n5290 = ~n2888 ;
  assign n2890 = n2878 & n5290 ;
  assign n2891 = n2889 | n2890 ;
  assign n5291 = ~n2697 ;
  assign n2892 = n2695 & n5291 ;
  assign n5292 = ~n341 ;
  assign n2893 = n5292 & n2714 ;
  assign n5293 = ~n2893 ;
  assign n2894 = n2713 & n5293 ;
  assign n2895 = n2892 & n2894 ;
  assign n2896 = n2892 | n2894 ;
  assign n5294 = ~n2895 ;
  assign n2897 = n5294 & n2896 ;
  assign n365 = x17 & x40 ;
  assign n366 = x18 & x39 ;
  assign n367 = x19 & x38 ;
  assign n675 = n366 & n367 ;
  assign n2898 = n366 | n367 ;
  assign n5295 = ~n675 ;
  assign n2899 = n5295 & n2898 ;
  assign n2900 = n365 & n2899 ;
  assign n2902 = n365 | n2899 ;
  assign n5296 = ~n2900 ;
  assign n2903 = n5296 & n2902 ;
  assign n5297 = ~n2903 ;
  assign n2904 = n2897 & n5297 ;
  assign n5298 = ~n2897 ;
  assign n2905 = n5298 & n2903 ;
  assign n2906 = n2904 | n2905 ;
  assign n2704 = n2693 & n2702 ;
  assign n2907 = n2694 & n2699 ;
  assign n2908 = n2704 | n2907 ;
  assign n2909 = n2906 | n2908 ;
  assign n2910 = n2906 & n2908 ;
  assign n5299 = ~n2910 ;
  assign n2911 = n2909 & n5299 ;
  assign n2912 = n2891 & n2911 ;
  assign n2913 = n2891 | n2911 ;
  assign n5300 = ~n2912 ;
  assign n2914 = n5300 & n2913 ;
  assign n2915 = n2672 | n2674 ;
  assign n368 = x12 & x45 ;
  assign n369 = x13 & x44 ;
  assign n370 = x11 & x46 ;
  assign n676 = n369 & n370 ;
  assign n2916 = n369 | n370 ;
  assign n5301 = ~n676 ;
  assign n2917 = n5301 & n2916 ;
  assign n2918 = n368 & n2917 ;
  assign n2920 = n368 | n2917 ;
  assign n5302 = ~n2918 ;
  assign n2921 = n5302 & n2920 ;
  assign n5303 = ~n2668 ;
  assign n2922 = n2666 & n5303 ;
  assign n373 = x14 & x43 ;
  assign n371 = x15 & x42 ;
  assign n372 = x16 & x41 ;
  assign n677 = n371 & n372 ;
  assign n2923 = n371 | n372 ;
  assign n5304 = ~n677 ;
  assign n2924 = n5304 & n2923 ;
  assign n5305 = ~n2924 ;
  assign n2925 = n373 & n5305 ;
  assign n5306 = ~n373 ;
  assign n2926 = n5306 & n2924 ;
  assign n2927 = n2925 | n2926 ;
  assign n2928 = n2922 | n2927 ;
  assign n2929 = n2922 & n2927 ;
  assign n5307 = ~n2929 ;
  assign n2930 = n2928 & n5307 ;
  assign n5308 = ~n2921 ;
  assign n2931 = n5308 & n2930 ;
  assign n5309 = ~n2930 ;
  assign n2932 = n2921 & n5309 ;
  assign n2933 = n2931 | n2932 ;
  assign n2934 = n2712 & n2717 ;
  assign n2935 = n2710 | n2934 ;
  assign n2936 = n2933 | n2935 ;
  assign n2937 = n2933 & n2935 ;
  assign n5310 = ~n2937 ;
  assign n2938 = n2936 & n5310 ;
  assign n5311 = ~n2915 ;
  assign n2939 = n5311 & n2938 ;
  assign n5312 = ~n2938 ;
  assign n2941 = n2915 & n5312 ;
  assign n2942 = n2939 | n2941 ;
  assign n5313 = ~n2726 ;
  assign n2943 = n2724 & n5313 ;
  assign n2944 = n2942 & n2943 ;
  assign n2945 = n2942 | n2943 ;
  assign n5314 = ~n2944 ;
  assign n2946 = n5314 & n2945 ;
  assign n2947 = n2914 & n2946 ;
  assign n2948 = n2914 | n2946 ;
  assign n5315 = ~n2947 ;
  assign n2949 = n5315 & n2948 ;
  assign n5316 = ~n2733 ;
  assign n2950 = n2730 & n5316 ;
  assign n2951 = n2949 & n2950 ;
  assign n2952 = n2949 | n2950 ;
  assign n5317 = ~n2951 ;
  assign n2953 = n5317 & n2952 ;
  assign n2954 = n2873 & n2953 ;
  assign n2955 = n2873 | n2953 ;
  assign n5318 = ~n2954 ;
  assign n2956 = n5318 & n2955 ;
  assign n5319 = ~n2777 ;
  assign n2786 = n5319 & n2784 ;
  assign n2957 = n2779 | n2781 ;
  assign n5320 = ~n2786 ;
  assign n2958 = n5320 & n2957 ;
  assign n2959 = n2642 & n2650 ;
  assign n5321 = ~n347 ;
  assign n2960 = n5321 & n2745 ;
  assign n5322 = ~n2960 ;
  assign n2961 = n2744 & n5322 ;
  assign n374 = x0 & x57 ;
  assign n375 = x1 & x56 ;
  assign n678 = n374 & n375 ;
  assign n2962 = n374 | n375 ;
  assign n5323 = ~n678 ;
  assign n2963 = n5323 & n2962 ;
  assign n2964 = n2961 & n2963 ;
  assign n2965 = n2961 | n2963 ;
  assign n5324 = ~n2964 ;
  assign n2966 = n5324 & n2965 ;
  assign n2967 = n2743 | n2748 ;
  assign n5325 = ~n2752 ;
  assign n2968 = n5325 & n2967 ;
  assign n2969 = n2966 & n2968 ;
  assign n2970 = n2966 | n2968 ;
  assign n5326 = ~n2969 ;
  assign n2971 = n5326 & n2970 ;
  assign n2973 = n2645 | n2648 ;
  assign n5327 = ~n2973 ;
  assign n2974 = n2971 & n5327 ;
  assign n5328 = ~n2971 ;
  assign n2975 = n5328 & n2973 ;
  assign n2976 = n2974 | n2975 ;
  assign n5329 = ~n2976 ;
  assign n2977 = n2959 & n5329 ;
  assign n5330 = ~n2959 ;
  assign n2978 = n5330 & n2976 ;
  assign n2979 = n2977 | n2978 ;
  assign n2980 = n2958 & n2979 ;
  assign n2981 = n2958 | n2979 ;
  assign n5331 = ~n2980 ;
  assign n2982 = n5331 & n2981 ;
  assign n5332 = ~n2792 ;
  assign n2983 = n2789 & n5332 ;
  assign n2984 = n2982 & n2983 ;
  assign n2985 = n2982 | n2983 ;
  assign n5333 = ~n2984 ;
  assign n2986 = n5333 & n2985 ;
  assign n2987 = n2956 & n2986 ;
  assign n2988 = n2956 | n2986 ;
  assign n5334 = ~n2987 ;
  assign n2989 = n5334 & n2988 ;
  assign n2990 = n2819 & n2989 ;
  assign n2991 = n2819 | n2989 ;
  assign n5335 = ~n2990 ;
  assign n2992 = n5335 & n2991 ;
  assign n2993 = n2796 & n2992 ;
  assign n2995 = n2796 | n2992 ;
  assign n5336 = ~n2993 ;
  assign n2996 = n5336 & n2995 ;
  assign n5337 = ~n2797 ;
  assign n2804 = n5337 & n2802 ;
  assign n2997 = n2474 | n2800 ;
  assign n5338 = ~n2804 ;
  assign n2998 = n5338 & n2997 ;
  assign n5339 = ~n2996 ;
  assign n2999 = n5339 & n2998 ;
  assign n5340 = ~n2998 ;
  assign n3000 = n2996 & n5340 ;
  assign n3001 = n2999 | n3000 ;
  assign n3002 = n2816 | n3001 ;
  assign n3003 = n2816 & n3001 ;
  assign n5341 = ~n3003 ;
  assign n90 = n3002 & n5341 ;
  assign n3005 = n2996 & n2998 ;
  assign n3006 = n3003 | n3005 ;
  assign n2994 = n5245 & n2992 ;
  assign n5342 = ~n2994 ;
  assign n3007 = n2991 & n5342 ;
  assign n376 = x4 & x54 ;
  assign n377 = x5 & x53 ;
  assign n378 = x3 & x55 ;
  assign n679 = n377 & n378 ;
  assign n3008 = n377 | n378 ;
  assign n5343 = ~n679 ;
  assign n3009 = n5343 & n3008 ;
  assign n3010 = n376 & n3009 ;
  assign n3012 = n376 | n3009 ;
  assign n5344 = ~n3010 ;
  assign n3013 = n5344 & n3012 ;
  assign n5345 = ~n351 ;
  assign n2825 = n5345 & n2823 ;
  assign n5346 = ~n2825 ;
  assign n3014 = n2822 & n5346 ;
  assign n379 = x6 & x52 ;
  assign n380 = x7 & x51 ;
  assign n381 = x8 & x50 ;
  assign n680 = n380 & n381 ;
  assign n3015 = n380 | n381 ;
  assign n5347 = ~n680 ;
  assign n3016 = n5347 & n3015 ;
  assign n3017 = n379 & n3016 ;
  assign n3019 = n379 | n3016 ;
  assign n5348 = ~n3017 ;
  assign n3020 = n5348 & n3019 ;
  assign n5349 = ~n3020 ;
  assign n3021 = n3014 & n5349 ;
  assign n5350 = ~n3014 ;
  assign n3022 = n5350 & n3020 ;
  assign n3023 = n3021 | n3022 ;
  assign n5351 = ~n3013 ;
  assign n3024 = n5351 & n3023 ;
  assign n5352 = ~n3023 ;
  assign n3025 = n3013 & n5352 ;
  assign n3026 = n3024 | n3025 ;
  assign n5353 = ~n368 ;
  assign n2919 = n5353 & n2917 ;
  assign n5354 = ~n2919 ;
  assign n3027 = n2916 & n5354 ;
  assign n5355 = ~n2848 ;
  assign n3028 = n2846 & n5355 ;
  assign n384 = x11 & x47 ;
  assign n382 = x9 & x49 ;
  assign n383 = x10 & x48 ;
  assign n681 = n382 & n383 ;
  assign n3029 = n382 | n383 ;
  assign n5356 = ~n681 ;
  assign n3030 = n5356 & n3029 ;
  assign n5357 = ~n3030 ;
  assign n3031 = n384 & n5357 ;
  assign n5358 = ~n384 ;
  assign n3032 = n5358 & n3030 ;
  assign n3033 = n3031 | n3032 ;
  assign n3034 = n3028 | n3033 ;
  assign n3035 = n3028 & n3033 ;
  assign n5359 = ~n3035 ;
  assign n3036 = n3034 & n5359 ;
  assign n3037 = n3027 & n3036 ;
  assign n3038 = n3027 | n3036 ;
  assign n5360 = ~n3037 ;
  assign n3039 = n5360 & n3038 ;
  assign n3040 = n2852 | n2854 ;
  assign n5361 = ~n3040 ;
  assign n3041 = n3039 & n5361 ;
  assign n5362 = ~n3039 ;
  assign n3042 = n5362 & n3040 ;
  assign n3043 = n3041 | n3042 ;
  assign n5363 = ~n3026 ;
  assign n3044 = n5363 & n3043 ;
  assign n5364 = ~n3043 ;
  assign n3046 = n3026 & n5364 ;
  assign n3047 = n3044 | n3046 ;
  assign n2940 = n2915 & n2938 ;
  assign n3048 = n2937 | n2940 ;
  assign n2863 = n2841 & n2861 ;
  assign n3049 = n2856 & n2858 ;
  assign n3050 = n2863 | n3049 ;
  assign n3051 = n3048 | n3050 ;
  assign n3052 = n3048 & n3050 ;
  assign n5365 = ~n3052 ;
  assign n3053 = n3051 & n5365 ;
  assign n3054 = n3047 & n3053 ;
  assign n3055 = n3047 | n3053 ;
  assign n5366 = ~n3054 ;
  assign n3056 = n5366 & n3055 ;
  assign n385 = x23 & x35 ;
  assign n386 = x26 & x32 ;
  assign n387 = x25 & x33 ;
  assign n682 = n386 & n387 ;
  assign n3057 = n386 | n387 ;
  assign n5367 = ~n682 ;
  assign n3058 = n5367 & n3057 ;
  assign n3059 = n385 & n3058 ;
  assign n3060 = n385 | n3058 ;
  assign n5368 = ~n3059 ;
  assign n3061 = n5368 & n3060 ;
  assign n5369 = ~n359 ;
  assign n3062 = n5369 & n2875 ;
  assign n5370 = ~n3062 ;
  assign n3063 = n2874 & n5370 ;
  assign n390 = x22 & x36 ;
  assign n388 = x21 & x37 ;
  assign n389 = x24 & x34 ;
  assign n683 = n388 & n389 ;
  assign n3064 = n388 | n389 ;
  assign n5371 = ~n683 ;
  assign n3065 = n5371 & n3064 ;
  assign n5372 = ~n3065 ;
  assign n3066 = n390 & n5372 ;
  assign n5373 = ~n390 ;
  assign n3067 = n5373 & n3065 ;
  assign n3068 = n3066 | n3067 ;
  assign n3069 = n3063 | n3068 ;
  assign n3070 = n3063 & n3068 ;
  assign n5374 = ~n3070 ;
  assign n3071 = n3069 & n5374 ;
  assign n5375 = ~n3061 ;
  assign n3072 = n5375 & n3071 ;
  assign n5376 = ~n3071 ;
  assign n3074 = n3061 & n5376 ;
  assign n3075 = n3072 | n3074 ;
  assign n5377 = ~n364 ;
  assign n3076 = n5377 & n2882 ;
  assign n5378 = ~n3076 ;
  assign n3077 = n2881 & n5378 ;
  assign n5379 = ~n365 ;
  assign n2901 = n5379 & n2899 ;
  assign n5380 = ~n2901 ;
  assign n3078 = n2898 & n5380 ;
  assign n3079 = n3077 & n3078 ;
  assign n3080 = n3077 | n3078 ;
  assign n5381 = ~n3079 ;
  assign n3081 = n5381 & n3080 ;
  assign n393 = x18 & x40 ;
  assign n391 = x19 & x39 ;
  assign n392 = x20 & x38 ;
  assign n684 = n391 & n392 ;
  assign n3082 = n391 | n392 ;
  assign n5382 = ~n684 ;
  assign n3083 = n5382 & n3082 ;
  assign n3084 = n393 & n3083 ;
  assign n3085 = n393 | n3083 ;
  assign n5383 = ~n3084 ;
  assign n3086 = n5383 & n3085 ;
  assign n5384 = ~n3086 ;
  assign n3087 = n3081 & n5384 ;
  assign n5385 = ~n3081 ;
  assign n3088 = n5385 & n3086 ;
  assign n3089 = n3087 | n3088 ;
  assign n3090 = n2880 | n2885 ;
  assign n5386 = ~n2889 ;
  assign n3091 = n5386 & n3090 ;
  assign n3092 = n3089 & n3091 ;
  assign n3093 = n3089 | n3091 ;
  assign n5387 = ~n3092 ;
  assign n3094 = n5387 & n3093 ;
  assign n3095 = n3075 & n3094 ;
  assign n3097 = n3075 | n3094 ;
  assign n5388 = ~n3095 ;
  assign n3098 = n5388 & n3097 ;
  assign n3099 = n2897 & n2903 ;
  assign n3100 = n2895 | n3099 ;
  assign n394 = x13 & x45 ;
  assign n395 = x12 & x46 ;
  assign n396 = x14 & x44 ;
  assign n685 = n395 & n396 ;
  assign n3101 = n395 | n396 ;
  assign n5389 = ~n685 ;
  assign n3102 = n5389 & n3101 ;
  assign n3103 = n394 & n3102 ;
  assign n3105 = n394 | n3102 ;
  assign n5390 = ~n3103 ;
  assign n3106 = n5390 & n3105 ;
  assign n5391 = ~n2926 ;
  assign n3107 = n2923 & n5391 ;
  assign n686 = x16 & x42 ;
  assign n397 = x15 & x43 ;
  assign n398 = x17 & x41 ;
  assign n687 = n397 & n398 ;
  assign n3108 = n397 | n398 ;
  assign n5392 = ~n687 ;
  assign n3109 = n5392 & n3108 ;
  assign n5393 = ~n686 ;
  assign n3110 = n5393 & n3109 ;
  assign n5394 = ~n3109 ;
  assign n3111 = n686 & n5394 ;
  assign n3112 = n3110 | n3111 ;
  assign n5395 = ~n3112 ;
  assign n3113 = n3107 & n5395 ;
  assign n5396 = ~n3107 ;
  assign n3114 = n5396 & n3112 ;
  assign n3115 = n3113 | n3114 ;
  assign n5397 = ~n3106 ;
  assign n3116 = n5397 & n3115 ;
  assign n5398 = ~n3115 ;
  assign n3118 = n3106 & n5398 ;
  assign n3119 = n3116 | n3118 ;
  assign n3120 = n2921 & n2930 ;
  assign n3121 = n2929 | n3120 ;
  assign n3122 = n3119 | n3121 ;
  assign n3123 = n3119 & n3121 ;
  assign n5399 = ~n3123 ;
  assign n3124 = n3122 & n5399 ;
  assign n5400 = ~n3100 ;
  assign n3125 = n5400 & n3124 ;
  assign n5401 = ~n3124 ;
  assign n3126 = n3100 & n5401 ;
  assign n3127 = n3125 | n3126 ;
  assign n3128 = n2910 | n2912 ;
  assign n3129 = n3127 | n3128 ;
  assign n3130 = n3127 & n3128 ;
  assign n5402 = ~n3130 ;
  assign n3131 = n3129 & n5402 ;
  assign n5403 = ~n3098 ;
  assign n3132 = n5403 & n3131 ;
  assign n5404 = ~n3131 ;
  assign n3133 = n3098 & n5404 ;
  assign n3134 = n3132 | n3133 ;
  assign n5405 = ~n2914 ;
  assign n3135 = n5405 & n2946 ;
  assign n5406 = ~n3135 ;
  assign n3136 = n2945 & n5406 ;
  assign n3137 = n3134 & n3136 ;
  assign n3138 = n3134 | n3136 ;
  assign n5407 = ~n3137 ;
  assign n3139 = n5407 & n3138 ;
  assign n5408 = ~n3056 ;
  assign n3140 = n5408 & n3139 ;
  assign n5409 = ~n3139 ;
  assign n3141 = n3056 & n5409 ;
  assign n3142 = n3140 | n3141 ;
  assign n3143 = n2821 & n2870 ;
  assign n3144 = n2868 | n3143 ;
  assign n2972 = n2648 & n2971 ;
  assign n5410 = ~n354 ;
  assign n2833 = n5410 & n2831 ;
  assign n5411 = ~n2833 ;
  assign n3145 = n2830 & n5411 ;
  assign n401 = x1 & x57 ;
  assign n399 = x0 & x58 ;
  assign n400 = x2 & x56 ;
  assign n3146 = n399 | n400 ;
  assign n3147 = n401 & n3146 ;
  assign n3148 = n2963 & n3147 ;
  assign n402 = x2 & x58 ;
  assign n5412 = ~n402 ;
  assign n3149 = n5412 & n3146 ;
  assign n5413 = ~n3149 ;
  assign n3150 = n328 & n5413 ;
  assign n3152 = n401 | n3146 ;
  assign n5414 = ~n3150 ;
  assign n3153 = n5414 & n3152 ;
  assign n5415 = ~n3148 ;
  assign n3154 = n5415 & n3153 ;
  assign n3155 = n3145 & n3154 ;
  assign n3156 = n3145 | n3154 ;
  assign n5416 = ~n3155 ;
  assign n3157 = n5416 & n3156 ;
  assign n3158 = n2829 | n2835 ;
  assign n5417 = ~n2839 ;
  assign n3159 = n5417 & n3158 ;
  assign n3160 = n2964 & n3159 ;
  assign n3161 = n2964 | n3159 ;
  assign n5418 = ~n3160 ;
  assign n3162 = n5418 & n3161 ;
  assign n3163 = n3157 & n3162 ;
  assign n3164 = n3157 | n3162 ;
  assign n5419 = ~n3163 ;
  assign n3165 = n5419 & n3164 ;
  assign n3166 = n2645 | n2969 ;
  assign n3167 = n2970 & n3166 ;
  assign n3168 = n3165 | n3167 ;
  assign n3169 = n3165 & n3167 ;
  assign n5420 = ~n3169 ;
  assign n3170 = n3168 & n5420 ;
  assign n3171 = n2972 & n3170 ;
  assign n3172 = n2972 | n3170 ;
  assign n5421 = ~n3171 ;
  assign n3173 = n5421 & n3172 ;
  assign n5422 = ~n3144 ;
  assign n3174 = n5422 & n3173 ;
  assign n5423 = ~n3173 ;
  assign n3175 = n3144 & n5423 ;
  assign n3176 = n3174 | n3175 ;
  assign n5424 = ~n2873 ;
  assign n3177 = n5424 & n2953 ;
  assign n5425 = ~n3177 ;
  assign n3178 = n2952 & n5425 ;
  assign n5426 = ~n3176 ;
  assign n3179 = n5426 & n3178 ;
  assign n5427 = ~n3178 ;
  assign n3180 = n3176 & n5427 ;
  assign n3181 = n3179 | n3180 ;
  assign n5428 = ~n3142 ;
  assign n3182 = n5428 & n3181 ;
  assign n5429 = ~n3181 ;
  assign n3183 = n3142 & n5429 ;
  assign n3184 = n3182 | n3183 ;
  assign n3185 = n2984 | n2987 ;
  assign n3186 = n2959 & n2976 ;
  assign n3187 = n2980 | n3186 ;
  assign n3188 = n3185 | n3187 ;
  assign n3189 = n3185 & n3187 ;
  assign n5430 = ~n3189 ;
  assign n3190 = n3188 & n5430 ;
  assign n5431 = ~n3184 ;
  assign n3191 = n5431 & n3190 ;
  assign n5432 = ~n3190 ;
  assign n3192 = n3184 & n5432 ;
  assign n3193 = n3191 | n3192 ;
  assign n5433 = ~n3193 ;
  assign n3194 = n3007 & n5433 ;
  assign n5434 = ~n3007 ;
  assign n3195 = n5434 & n3193 ;
  assign n3196 = n3194 | n3195 ;
  assign n3197 = n3006 & n3196 ;
  assign n3198 = n3006 | n3196 ;
  assign n5435 = ~n3197 ;
  assign n91 = n5435 & n3198 ;
  assign n3200 = n3007 & n3193 ;
  assign n3201 = n3197 | n3200 ;
  assign n403 = x4 & x55 ;
  assign n404 = x6 & x53 ;
  assign n405 = x5 & x54 ;
  assign n688 = n404 & n405 ;
  assign n3202 = n404 | n405 ;
  assign n5436 = ~n688 ;
  assign n3203 = n5436 & n3202 ;
  assign n3204 = n403 & n3203 ;
  assign n3205 = n403 | n3203 ;
  assign n5437 = ~n3204 ;
  assign n3206 = n5437 & n3205 ;
  assign n5438 = ~n379 ;
  assign n3018 = n5438 & n3016 ;
  assign n5439 = ~n3018 ;
  assign n3207 = n3015 & n5439 ;
  assign n406 = x7 & x52 ;
  assign n407 = x8 & x51 ;
  assign n408 = x9 & x50 ;
  assign n689 = n407 & n408 ;
  assign n3208 = n407 | n408 ;
  assign n5440 = ~n689 ;
  assign n3209 = n5440 & n3208 ;
  assign n3210 = n406 & n3209 ;
  assign n3212 = n406 | n3209 ;
  assign n5441 = ~n3210 ;
  assign n3213 = n5441 & n3212 ;
  assign n5442 = ~n3213 ;
  assign n3214 = n3207 & n5442 ;
  assign n5443 = ~n3207 ;
  assign n3215 = n5443 & n3213 ;
  assign n3216 = n3214 | n3215 ;
  assign n5444 = ~n3206 ;
  assign n3217 = n5444 & n3216 ;
  assign n5445 = ~n3216 ;
  assign n3218 = n3206 & n5445 ;
  assign n3219 = n3217 | n3218 ;
  assign n5446 = ~n394 ;
  assign n3104 = n5446 & n3102 ;
  assign n5447 = ~n3104 ;
  assign n3220 = n3101 & n5447 ;
  assign n5448 = ~n3032 ;
  assign n3221 = n3029 & n5448 ;
  assign n690 = x10 & x49 ;
  assign n409 = x11 & x48 ;
  assign n410 = x12 & x47 ;
  assign n691 = n409 & n410 ;
  assign n3222 = n409 | n410 ;
  assign n5449 = ~n691 ;
  assign n3223 = n5449 & n3222 ;
  assign n5450 = ~n690 ;
  assign n3224 = n5450 & n3223 ;
  assign n5451 = ~n3223 ;
  assign n3225 = n690 & n5451 ;
  assign n3226 = n3224 | n3225 ;
  assign n3227 = n3221 | n3226 ;
  assign n3228 = n3221 & n3226 ;
  assign n5452 = ~n3228 ;
  assign n3229 = n3227 & n5452 ;
  assign n3230 = n3220 & n3229 ;
  assign n3231 = n3220 | n3229 ;
  assign n5453 = ~n3230 ;
  assign n3232 = n5453 & n3231 ;
  assign n3233 = n3035 | n3037 ;
  assign n5454 = ~n3233 ;
  assign n3234 = n3232 & n5454 ;
  assign n5455 = ~n3232 ;
  assign n3235 = n5455 & n3233 ;
  assign n3236 = n3234 | n3235 ;
  assign n5456 = ~n3219 ;
  assign n3237 = n5456 & n3236 ;
  assign n5457 = ~n3236 ;
  assign n3239 = n3219 & n5457 ;
  assign n3240 = n3237 | n3239 ;
  assign n3045 = n3026 & n3043 ;
  assign n3241 = n3039 & n3040 ;
  assign n3242 = n3045 | n3241 ;
  assign n5458 = ~n3125 ;
  assign n3243 = n3122 & n5458 ;
  assign n5459 = ~n3242 ;
  assign n3244 = n5459 & n3243 ;
  assign n5460 = ~n3243 ;
  assign n3245 = n3242 & n5460 ;
  assign n3246 = n3244 | n3245 ;
  assign n3247 = n3240 & n3246 ;
  assign n3248 = n3240 | n3246 ;
  assign n5461 = ~n3247 ;
  assign n3249 = n5461 & n3248 ;
  assign n3250 = n3098 & n3131 ;
  assign n3251 = n3130 | n3250 ;
  assign n5462 = ~n3075 ;
  assign n3096 = n5462 & n3094 ;
  assign n5463 = ~n3096 ;
  assign n3252 = n3093 & n5463 ;
  assign n5464 = ~n3110 ;
  assign n3253 = n3108 & n5464 ;
  assign n411 = x14 & x45 ;
  assign n412 = x13 & x46 ;
  assign n413 = x15 & x44 ;
  assign n692 = n412 & n413 ;
  assign n3254 = n412 | n413 ;
  assign n5465 = ~n692 ;
  assign n3255 = n5465 & n3254 ;
  assign n3256 = n411 & n3255 ;
  assign n3258 = n411 | n3255 ;
  assign n5466 = ~n3256 ;
  assign n3259 = n5466 & n3258 ;
  assign n416 = x16 & x43 ;
  assign n414 = x17 & x42 ;
  assign n415 = x18 & x41 ;
  assign n693 = n414 & n415 ;
  assign n3260 = n414 | n415 ;
  assign n5467 = ~n693 ;
  assign n3261 = n5467 & n3260 ;
  assign n5468 = ~n3261 ;
  assign n3262 = n416 & n5468 ;
  assign n5469 = ~n416 ;
  assign n3263 = n5469 & n3261 ;
  assign n3264 = n3262 | n3263 ;
  assign n3265 = n3259 | n3264 ;
  assign n3266 = n3259 & n3264 ;
  assign n5470 = ~n3266 ;
  assign n3267 = n3265 & n5470 ;
  assign n3268 = n3253 & n3267 ;
  assign n3269 = n3253 | n3267 ;
  assign n5471 = ~n3268 ;
  assign n3270 = n5471 & n3269 ;
  assign n3117 = n3106 & n3115 ;
  assign n3271 = n3107 & n3112 ;
  assign n3272 = n3117 | n3271 ;
  assign n3273 = n3081 & n3086 ;
  assign n3274 = n3079 | n3273 ;
  assign n3275 = n3272 | n3274 ;
  assign n3276 = n3272 & n3274 ;
  assign n5472 = ~n3276 ;
  assign n3277 = n3275 & n5472 ;
  assign n5473 = ~n3270 ;
  assign n3278 = n5473 & n3277 ;
  assign n5474 = ~n3277 ;
  assign n3279 = n3270 & n5474 ;
  assign n3280 = n3278 | n3279 ;
  assign n3073 = n3061 & n3071 ;
  assign n3281 = n3070 | n3073 ;
  assign n5475 = ~n3067 ;
  assign n3282 = n3064 & n5475 ;
  assign n5476 = ~n393 ;
  assign n3283 = n5476 & n3083 ;
  assign n5477 = ~n3283 ;
  assign n3284 = n3082 & n5477 ;
  assign n3285 = n3282 & n3284 ;
  assign n3286 = n3282 | n3284 ;
  assign n5478 = ~n3285 ;
  assign n3287 = n5478 & n3286 ;
  assign n419 = x19 & x40 ;
  assign n417 = x20 & x39 ;
  assign n418 = x21 & x38 ;
  assign n694 = n417 & n418 ;
  assign n3288 = n417 | n418 ;
  assign n5479 = ~n694 ;
  assign n3289 = n5479 & n3288 ;
  assign n3290 = n419 & n3289 ;
  assign n3291 = n419 | n3289 ;
  assign n5480 = ~n3290 ;
  assign n3292 = n5480 & n3291 ;
  assign n5481 = ~n3292 ;
  assign n3293 = n3287 & n5481 ;
  assign n5482 = ~n3287 ;
  assign n3294 = n5482 & n3292 ;
  assign n3295 = n3293 | n3294 ;
  assign n420 = x23 & x36 ;
  assign n421 = x22 & x37 ;
  assign n422 = x25 & x34 ;
  assign n695 = n421 & n422 ;
  assign n3296 = n421 | n422 ;
  assign n5483 = ~n695 ;
  assign n3297 = n5483 & n3296 ;
  assign n3298 = n420 & n3297 ;
  assign n3299 = n420 | n3297 ;
  assign n5484 = ~n3298 ;
  assign n3300 = n5484 & n3299 ;
  assign n5485 = ~n385 ;
  assign n3301 = n5485 & n3058 ;
  assign n5486 = ~n3301 ;
  assign n3302 = n3057 & n5486 ;
  assign n696 = x24 & x35 ;
  assign n423 = x26 & x33 ;
  assign n424 = x27 & x32 ;
  assign n697 = n423 & n424 ;
  assign n3303 = n423 | n424 ;
  assign n5487 = ~n697 ;
  assign n3304 = n5487 & n3303 ;
  assign n5488 = ~n696 ;
  assign n3305 = n5488 & n3304 ;
  assign n5489 = ~n3304 ;
  assign n3306 = n696 & n5489 ;
  assign n3307 = n3305 | n3306 ;
  assign n3308 = n3302 | n3307 ;
  assign n3309 = n3302 & n3307 ;
  assign n5490 = ~n3309 ;
  assign n3310 = n3308 & n5490 ;
  assign n3311 = n3300 & n3310 ;
  assign n3312 = n3300 | n3310 ;
  assign n5491 = ~n3311 ;
  assign n3313 = n5491 & n3312 ;
  assign n3314 = n3295 & n3313 ;
  assign n3315 = n3295 | n3313 ;
  assign n5492 = ~n3314 ;
  assign n3316 = n5492 & n3315 ;
  assign n5493 = ~n3281 ;
  assign n3317 = n5493 & n3316 ;
  assign n5494 = ~n3316 ;
  assign n3318 = n3281 & n5494 ;
  assign n3319 = n3317 | n3318 ;
  assign n3320 = n3280 | n3319 ;
  assign n3321 = n3280 & n3319 ;
  assign n5495 = ~n3321 ;
  assign n3322 = n3320 & n5495 ;
  assign n3323 = n3252 & n3322 ;
  assign n3324 = n3252 | n3322 ;
  assign n5496 = ~n3323 ;
  assign n3325 = n5496 & n3324 ;
  assign n3326 = n3251 & n3325 ;
  assign n3327 = n3251 | n3325 ;
  assign n5497 = ~n3326 ;
  assign n3328 = n5497 & n3327 ;
  assign n3329 = n3249 & n3328 ;
  assign n3330 = n3249 | n3328 ;
  assign n5498 = ~n3329 ;
  assign n3331 = n5498 & n3330 ;
  assign n5499 = ~n3047 ;
  assign n3332 = n5499 & n3053 ;
  assign n5500 = ~n3332 ;
  assign n3333 = n3051 & n5500 ;
  assign n3334 = n3014 | n3020 ;
  assign n5501 = ~n3024 ;
  assign n3335 = n5501 & n3334 ;
  assign n3151 = n401 & n3150 ;
  assign n3336 = n3151 | n3155 ;
  assign n698 = n399 & n400 ;
  assign n3337 = n698 | n3147 ;
  assign n5502 = ~n376 ;
  assign n3011 = n5502 & n3009 ;
  assign n5503 = ~n3011 ;
  assign n3338 = n3008 & n5503 ;
  assign n427 = x2 & x57 ;
  assign n425 = x1 & x58 ;
  assign n426 = x3 & x56 ;
  assign n699 = n425 & n426 ;
  assign n3339 = n425 | n426 ;
  assign n5504 = ~n699 ;
  assign n3340 = n5504 & n3339 ;
  assign n5505 = ~n3340 ;
  assign n3341 = n427 & n5505 ;
  assign n5506 = ~n427 ;
  assign n3342 = n5506 & n3340 ;
  assign n3343 = n3341 | n3342 ;
  assign n5507 = ~n3343 ;
  assign n3344 = n3338 & n5507 ;
  assign n5508 = ~n3338 ;
  assign n3345 = n5508 & n3343 ;
  assign n3346 = n3344 | n3345 ;
  assign n5509 = ~n3337 ;
  assign n3347 = n5509 & n3346 ;
  assign n5510 = ~n3346 ;
  assign n3348 = n3337 & n5510 ;
  assign n3349 = n3347 | n3348 ;
  assign n5511 = ~n3336 ;
  assign n3350 = n5511 & n3349 ;
  assign n5512 = ~n3349 ;
  assign n3351 = n3336 & n5512 ;
  assign n3352 = n3350 | n3351 ;
  assign n3353 = n3335 & n3352 ;
  assign n3354 = n3335 | n3352 ;
  assign n5513 = ~n3353 ;
  assign n3355 = n5513 & n3354 ;
  assign n428 = x0 & x59 ;
  assign n5514 = ~n3157 ;
  assign n3356 = n5514 & n3162 ;
  assign n5515 = ~n3356 ;
  assign n3357 = n3161 & n5515 ;
  assign n3358 = n428 & n3357 ;
  assign n3359 = n428 | n3357 ;
  assign n5516 = ~n3358 ;
  assign n3360 = n5516 & n3359 ;
  assign n3361 = n3355 & n3360 ;
  assign n3362 = n3355 | n3360 ;
  assign n5517 = ~n3361 ;
  assign n3363 = n5517 & n3362 ;
  assign n3364 = n3169 & n3363 ;
  assign n3365 = n3169 | n3363 ;
  assign n5518 = ~n3364 ;
  assign n3366 = n5518 & n3365 ;
  assign n5519 = ~n3333 ;
  assign n3367 = n5519 & n3366 ;
  assign n5520 = ~n3366 ;
  assign n3368 = n3333 & n5520 ;
  assign n3369 = n3367 | n3368 ;
  assign n3370 = n3056 & n3139 ;
  assign n3371 = n3137 | n3370 ;
  assign n3372 = n3369 | n3371 ;
  assign n3373 = n3369 & n3371 ;
  assign n5521 = ~n3373 ;
  assign n3374 = n3372 & n5521 ;
  assign n3375 = n3331 & n3374 ;
  assign n3376 = n3331 | n3374 ;
  assign n5522 = ~n3375 ;
  assign n3377 = n5522 & n3376 ;
  assign n3378 = n3176 & n3178 ;
  assign n3379 = n3142 & n3181 ;
  assign n3380 = n3378 | n3379 ;
  assign n5523 = ~n3174 ;
  assign n3381 = n3172 & n5523 ;
  assign n3382 = n3380 & n3381 ;
  assign n3383 = n3380 | n3381 ;
  assign n5524 = ~n3382 ;
  assign n3384 = n5524 & n3383 ;
  assign n3385 = n3377 & n3384 ;
  assign n3386 = n3377 | n3384 ;
  assign n5525 = ~n3385 ;
  assign n3387 = n5525 & n3386 ;
  assign n5526 = ~n3191 ;
  assign n3388 = n3188 & n5526 ;
  assign n3389 = n3387 & n3388 ;
  assign n3390 = n3387 | n3388 ;
  assign n5527 = ~n3389 ;
  assign n3391 = n5527 & n3390 ;
  assign n5528 = ~n3201 ;
  assign n3392 = n5528 & n3391 ;
  assign n5529 = ~n3391 ;
  assign n3393 = n3201 & n5529 ;
  assign n92 = n3392 | n3393 ;
  assign n5530 = ~n3392 ;
  assign n3395 = n3390 & n5530 ;
  assign n3238 = n3219 & n3236 ;
  assign n3396 = n3232 & n3233 ;
  assign n3397 = n3238 | n3396 ;
  assign n429 = x10 & x50 ;
  assign n430 = x9 & x51 ;
  assign n431 = x8 & x52 ;
  assign n700 = n430 & n431 ;
  assign n3398 = n430 | n431 ;
  assign n5531 = ~n700 ;
  assign n3399 = n5531 & n3398 ;
  assign n3400 = n429 & n3399 ;
  assign n3402 = n429 | n3399 ;
  assign n5532 = ~n3400 ;
  assign n3403 = n5532 & n3402 ;
  assign n5533 = ~n406 ;
  assign n3211 = n5533 & n3209 ;
  assign n5534 = ~n3211 ;
  assign n3404 = n3208 & n5534 ;
  assign n432 = x6 & x54 ;
  assign n433 = x5 & x55 ;
  assign n434 = x7 & x53 ;
  assign n701 = n433 & n434 ;
  assign n3405 = n433 | n434 ;
  assign n5535 = ~n701 ;
  assign n3406 = n5535 & n3405 ;
  assign n3407 = n432 & n3406 ;
  assign n3408 = n432 | n3406 ;
  assign n5536 = ~n3407 ;
  assign n3409 = n5536 & n3408 ;
  assign n5537 = ~n3409 ;
  assign n3410 = n3404 & n5537 ;
  assign n5538 = ~n3404 ;
  assign n3411 = n5538 & n3409 ;
  assign n3412 = n3410 | n3411 ;
  assign n5539 = ~n3403 ;
  assign n3413 = n5539 & n3412 ;
  assign n5540 = ~n3412 ;
  assign n3414 = n3403 & n5540 ;
  assign n3415 = n3413 | n3414 ;
  assign n5541 = ~n3224 ;
  assign n3416 = n3222 & n5541 ;
  assign n5542 = ~n411 ;
  assign n3257 = n5542 & n3255 ;
  assign n5543 = ~n3257 ;
  assign n3417 = n3254 & n5543 ;
  assign n702 = x12 & x48 ;
  assign n435 = x11 & x49 ;
  assign n436 = x13 & x47 ;
  assign n703 = n435 & n436 ;
  assign n3418 = n435 | n436 ;
  assign n5544 = ~n703 ;
  assign n3419 = n5544 & n3418 ;
  assign n5545 = ~n702 ;
  assign n3420 = n5545 & n3419 ;
  assign n5546 = ~n3419 ;
  assign n3421 = n702 & n5546 ;
  assign n3422 = n3420 | n3421 ;
  assign n5547 = ~n3422 ;
  assign n3423 = n3417 & n5547 ;
  assign n5548 = ~n3417 ;
  assign n3424 = n5548 & n3422 ;
  assign n3425 = n3423 | n3424 ;
  assign n3426 = n3416 & n3425 ;
  assign n3427 = n3416 | n3425 ;
  assign n5549 = ~n3426 ;
  assign n3428 = n5549 & n3427 ;
  assign n3429 = n3228 | n3230 ;
  assign n5550 = ~n3429 ;
  assign n3430 = n3428 & n5550 ;
  assign n5551 = ~n3428 ;
  assign n3431 = n5551 & n3429 ;
  assign n3432 = n3430 | n3431 ;
  assign n5552 = ~n3415 ;
  assign n3433 = n5552 & n3432 ;
  assign n5553 = ~n3432 ;
  assign n3435 = n3415 & n5553 ;
  assign n3436 = n3433 | n3435 ;
  assign n5554 = ~n3278 ;
  assign n3437 = n3275 & n5554 ;
  assign n3438 = n3436 & n3437 ;
  assign n3439 = n3436 | n3437 ;
  assign n5555 = ~n3438 ;
  assign n3440 = n5555 & n3439 ;
  assign n5556 = ~n3397 ;
  assign n3441 = n5556 & n3440 ;
  assign n5557 = ~n3440 ;
  assign n3442 = n3397 & n5557 ;
  assign n3443 = n3441 | n3442 ;
  assign n5558 = ~n3317 ;
  assign n3444 = n3315 & n5558 ;
  assign n437 = x14 & x46 ;
  assign n438 = x16 & x44 ;
  assign n439 = x15 & x45 ;
  assign n704 = n438 & n439 ;
  assign n3445 = n438 | n439 ;
  assign n5559 = ~n704 ;
  assign n3446 = n5559 & n3445 ;
  assign n3447 = n437 & n3446 ;
  assign n3448 = n437 | n3446 ;
  assign n5560 = ~n3447 ;
  assign n3449 = n5560 & n3448 ;
  assign n5561 = ~n3263 ;
  assign n3450 = n3260 & n5561 ;
  assign n705 = x17 & x43 ;
  assign n440 = x18 & x42 ;
  assign n441 = x19 & x41 ;
  assign n706 = n440 & n441 ;
  assign n3451 = n440 | n441 ;
  assign n5562 = ~n706 ;
  assign n3452 = n5562 & n3451 ;
  assign n5563 = ~n705 ;
  assign n3453 = n5563 & n3452 ;
  assign n5564 = ~n3452 ;
  assign n3454 = n705 & n5564 ;
  assign n3455 = n3453 | n3454 ;
  assign n3456 = n3450 | n3455 ;
  assign n3457 = n3450 & n3455 ;
  assign n5565 = ~n3457 ;
  assign n3458 = n3456 & n5565 ;
  assign n5566 = ~n3449 ;
  assign n3459 = n5566 & n3458 ;
  assign n5567 = ~n3458 ;
  assign n3460 = n3449 & n5567 ;
  assign n3461 = n3459 | n3460 ;
  assign n3462 = n3266 | n3268 ;
  assign n3463 = n3287 & n3292 ;
  assign n3464 = n3285 | n3463 ;
  assign n3465 = n3462 | n3464 ;
  assign n3466 = n3462 & n3464 ;
  assign n5568 = ~n3466 ;
  assign n3467 = n3465 & n5568 ;
  assign n5569 = ~n3461 ;
  assign n3468 = n5569 & n3467 ;
  assign n5570 = ~n3467 ;
  assign n3469 = n3461 & n5570 ;
  assign n3470 = n3468 | n3469 ;
  assign n5571 = ~n419 ;
  assign n3471 = n5571 & n3289 ;
  assign n5572 = ~n3471 ;
  assign n3472 = n3288 & n5572 ;
  assign n5573 = ~n420 ;
  assign n3473 = n5573 & n3297 ;
  assign n5574 = ~n3473 ;
  assign n3474 = n3296 & n5574 ;
  assign n3475 = n3472 & n3474 ;
  assign n3476 = n3472 | n3474 ;
  assign n5575 = ~n3475 ;
  assign n3477 = n5575 & n3476 ;
  assign n444 = x20 & x40 ;
  assign n442 = x21 & x39 ;
  assign n443 = x22 & x38 ;
  assign n707 = n442 & n443 ;
  assign n3478 = n442 | n443 ;
  assign n5576 = ~n707 ;
  assign n3479 = n5576 & n3478 ;
  assign n3480 = n444 & n3479 ;
  assign n3481 = n444 | n3479 ;
  assign n5577 = ~n3480 ;
  assign n3482 = n5577 & n3481 ;
  assign n5578 = ~n3482 ;
  assign n3483 = n3477 & n5578 ;
  assign n5579 = ~n3477 ;
  assign n3484 = n5579 & n3482 ;
  assign n3485 = n3483 | n3484 ;
  assign n708 = x25 & x35 ;
  assign n445 = x27 & x33 ;
  assign n446 = x28 & x32 ;
  assign n709 = n445 & n446 ;
  assign n3486 = n445 | n446 ;
  assign n5580 = ~n709 ;
  assign n3487 = n5580 & n3486 ;
  assign n5581 = ~n708 ;
  assign n3488 = n5581 & n3487 ;
  assign n5582 = ~n3487 ;
  assign n3489 = n708 & n5582 ;
  assign n3490 = n3488 | n3489 ;
  assign n5583 = ~n3305 ;
  assign n3491 = n3303 & n5583 ;
  assign n710 = x23 & x37 ;
  assign n447 = x24 & x36 ;
  assign n448 = x26 & x34 ;
  assign n711 = n447 & n448 ;
  assign n3492 = n447 | n448 ;
  assign n5584 = ~n711 ;
  assign n3493 = n5584 & n3492 ;
  assign n5585 = ~n710 ;
  assign n3494 = n5585 & n3493 ;
  assign n5586 = ~n3493 ;
  assign n3495 = n710 & n5586 ;
  assign n3496 = n3494 | n3495 ;
  assign n5587 = ~n3496 ;
  assign n3497 = n3491 & n5587 ;
  assign n5588 = ~n3491 ;
  assign n3498 = n5588 & n3496 ;
  assign n3499 = n3497 | n3498 ;
  assign n5589 = ~n3490 ;
  assign n3500 = n5589 & n3499 ;
  assign n5590 = ~n3499 ;
  assign n3502 = n3490 & n5590 ;
  assign n3503 = n3500 | n3502 ;
  assign n3504 = n3309 | n3311 ;
  assign n3505 = n3503 | n3504 ;
  assign n3506 = n3503 & n3504 ;
  assign n5591 = ~n3506 ;
  assign n3507 = n3505 & n5591 ;
  assign n5592 = ~n3485 ;
  assign n3508 = n5592 & n3507 ;
  assign n5593 = ~n3507 ;
  assign n3509 = n3485 & n5593 ;
  assign n3510 = n3508 | n3509 ;
  assign n3511 = n3470 | n3510 ;
  assign n3512 = n3470 & n3510 ;
  assign n5594 = ~n3512 ;
  assign n3513 = n3511 & n5594 ;
  assign n5595 = ~n3444 ;
  assign n3514 = n5595 & n3513 ;
  assign n5596 = ~n3513 ;
  assign n3515 = n3444 & n5596 ;
  assign n3516 = n3514 | n3515 ;
  assign n3517 = n3321 | n3323 ;
  assign n3518 = n3516 | n3517 ;
  assign n3519 = n3516 & n3517 ;
  assign n5597 = ~n3519 ;
  assign n3520 = n3518 & n5597 ;
  assign n5598 = ~n3443 ;
  assign n3521 = n5598 & n3520 ;
  assign n5599 = ~n3520 ;
  assign n3522 = n3443 & n5599 ;
  assign n3523 = n3521 | n3522 ;
  assign n3524 = n3242 | n3243 ;
  assign n5600 = ~n3240 ;
  assign n3525 = n5600 & n3246 ;
  assign n5601 = ~n3525 ;
  assign n3526 = n3524 & n5601 ;
  assign n3527 = n3336 | n3349 ;
  assign n5602 = ~n3335 ;
  assign n3528 = n5602 & n3352 ;
  assign n5603 = ~n3528 ;
  assign n3529 = n3527 & n5603 ;
  assign n3530 = n3207 | n3213 ;
  assign n5604 = ~n3217 ;
  assign n3531 = n5604 & n3530 ;
  assign n5605 = ~n3342 ;
  assign n3532 = n3339 & n5605 ;
  assign n5606 = ~n403 ;
  assign n3533 = n5606 & n3203 ;
  assign n5607 = ~n3533 ;
  assign n3534 = n3202 & n5607 ;
  assign n449 = x3 & x57 ;
  assign n450 = x4 & x56 ;
  assign n712 = n449 & n450 ;
  assign n3535 = n449 | n450 ;
  assign n5608 = ~n712 ;
  assign n3536 = n5608 & n3535 ;
  assign n3537 = n5412 & n3536 ;
  assign n5609 = ~n3536 ;
  assign n3538 = n402 & n5609 ;
  assign n3539 = n3537 | n3538 ;
  assign n3540 = n3534 | n3539 ;
  assign n3541 = n3534 & n3539 ;
  assign n5610 = ~n3541 ;
  assign n3542 = n3540 & n5610 ;
  assign n3543 = n3532 & n3542 ;
  assign n3544 = n3532 | n3542 ;
  assign n5611 = ~n3543 ;
  assign n3545 = n5611 & n3544 ;
  assign n3546 = n3338 & n3343 ;
  assign n3547 = n3337 & n3346 ;
  assign n3548 = n3546 | n3547 ;
  assign n5612 = ~n3548 ;
  assign n3549 = n3545 & n5612 ;
  assign n5613 = ~n3545 ;
  assign n3550 = n5613 & n3548 ;
  assign n3551 = n3549 | n3550 ;
  assign n3552 = n3531 & n3551 ;
  assign n3553 = n3531 | n3551 ;
  assign n5614 = ~n3552 ;
  assign n3554 = n5614 & n3553 ;
  assign n451 = x1 & x60 ;
  assign n452 = n428 & n451 ;
  assign n713 = x1 & x59 ;
  assign n714 = x0 & x60 ;
  assign n3555 = n713 | n714 ;
  assign n5615 = ~n452 ;
  assign n3556 = n5615 & n3555 ;
  assign n3557 = n3554 & n3556 ;
  assign n3558 = n3554 | n3556 ;
  assign n5616 = ~n3557 ;
  assign n3559 = n5616 & n3558 ;
  assign n5617 = ~n3529 ;
  assign n3560 = n5617 & n3559 ;
  assign n5618 = ~n3559 ;
  assign n3561 = n3529 & n5618 ;
  assign n3562 = n3560 | n3561 ;
  assign n3563 = n3358 | n3361 ;
  assign n3564 = n3562 | n3563 ;
  assign n3565 = n3562 & n3563 ;
  assign n5619 = ~n3565 ;
  assign n3566 = n3564 & n5619 ;
  assign n3567 = n3526 & n3566 ;
  assign n3568 = n3526 | n3566 ;
  assign n5620 = ~n3567 ;
  assign n3569 = n5620 & n3568 ;
  assign n3570 = n3326 | n3329 ;
  assign n3571 = n3569 | n3570 ;
  assign n3572 = n3569 & n3570 ;
  assign n5621 = ~n3572 ;
  assign n3573 = n3571 & n5621 ;
  assign n5622 = ~n3523 ;
  assign n3574 = n5622 & n3573 ;
  assign n5623 = ~n3573 ;
  assign n3575 = n3523 & n5623 ;
  assign n3576 = n3574 | n3575 ;
  assign n5624 = ~n3331 ;
  assign n3577 = n5624 & n3374 ;
  assign n5625 = ~n3577 ;
  assign n3578 = n3372 & n5625 ;
  assign n5626 = ~n3367 ;
  assign n3579 = n3365 & n5626 ;
  assign n3580 = n3578 & n3579 ;
  assign n3581 = n3578 | n3579 ;
  assign n5627 = ~n3580 ;
  assign n3582 = n5627 & n3581 ;
  assign n5628 = ~n3576 ;
  assign n3583 = n5628 & n3582 ;
  assign n5629 = ~n3582 ;
  assign n3584 = n3576 & n5629 ;
  assign n3585 = n3583 | n3584 ;
  assign n3586 = n3382 | n3385 ;
  assign n3587 = n3585 | n3586 ;
  assign n3588 = n3585 & n3586 ;
  assign n5630 = ~n3588 ;
  assign n3589 = n3587 & n5630 ;
  assign n3590 = n3395 & n3589 ;
  assign n3591 = n3395 | n3589 ;
  assign n5631 = ~n3590 ;
  assign n93 = n5631 & n3591 ;
  assign n3593 = n3588 | n3590 ;
  assign n453 = x26 & x35 ;
  assign n454 = x28 & x33 ;
  assign n455 = x29 & x32 ;
  assign n715 = n454 & n455 ;
  assign n3594 = n454 | n455 ;
  assign n5632 = ~n715 ;
  assign n3595 = n5632 & n3594 ;
  assign n3596 = n453 & n3595 ;
  assign n3597 = n453 | n3595 ;
  assign n5633 = ~n3596 ;
  assign n3598 = n5633 & n3597 ;
  assign n5634 = ~n3488 ;
  assign n3599 = n3486 & n5634 ;
  assign n5635 = ~n3598 ;
  assign n3600 = n5635 & n3599 ;
  assign n5636 = ~n3599 ;
  assign n3601 = n3598 & n5636 ;
  assign n3602 = n3600 | n3601 ;
  assign n458 = x25 & x36 ;
  assign n456 = x24 & x37 ;
  assign n457 = x27 & x34 ;
  assign n716 = n456 & n457 ;
  assign n3603 = n456 | n457 ;
  assign n5637 = ~n716 ;
  assign n3604 = n5637 & n3603 ;
  assign n5638 = ~n3604 ;
  assign n3605 = n458 & n5638 ;
  assign n5639 = ~n458 ;
  assign n3606 = n5639 & n3604 ;
  assign n3607 = n3605 | n3606 ;
  assign n5640 = ~n3607 ;
  assign n3608 = n3602 & n5640 ;
  assign n5641 = ~n3602 ;
  assign n3609 = n5641 & n3607 ;
  assign n3610 = n3608 | n3609 ;
  assign n5642 = ~n3494 ;
  assign n3611 = n3492 & n5642 ;
  assign n5643 = ~n444 ;
  assign n3612 = n5643 & n3479 ;
  assign n5644 = ~n3612 ;
  assign n3613 = n3478 & n5644 ;
  assign n461 = x21 & x40 ;
  assign n459 = x22 & x39 ;
  assign n460 = x23 & x38 ;
  assign n717 = n459 & n460 ;
  assign n3614 = n459 | n460 ;
  assign n5645 = ~n717 ;
  assign n3615 = n5645 & n3614 ;
  assign n5646 = ~n3615 ;
  assign n3616 = n461 & n5646 ;
  assign n5647 = ~n461 ;
  assign n3617 = n5647 & n3615 ;
  assign n3618 = n3616 | n3617 ;
  assign n3619 = n3613 | n3618 ;
  assign n3620 = n3613 & n3618 ;
  assign n5648 = ~n3620 ;
  assign n3621 = n3619 & n5648 ;
  assign n5649 = ~n3611 ;
  assign n3622 = n5649 & n3621 ;
  assign n5650 = ~n3621 ;
  assign n3623 = n3611 & n5650 ;
  assign n3624 = n3622 | n3623 ;
  assign n3501 = n3490 & n3499 ;
  assign n3625 = n3491 & n3496 ;
  assign n3626 = n3501 | n3625 ;
  assign n3627 = n3624 | n3626 ;
  assign n3628 = n3624 & n3626 ;
  assign n5651 = ~n3628 ;
  assign n3629 = n3627 & n5651 ;
  assign n3630 = n3610 & n3629 ;
  assign n3631 = n3610 | n3629 ;
  assign n5652 = ~n3630 ;
  assign n3632 = n5652 & n3631 ;
  assign n5653 = ~n3453 ;
  assign n3633 = n3451 & n5653 ;
  assign n462 = x18 & x43 ;
  assign n463 = x19 & x42 ;
  assign n464 = x20 & x41 ;
  assign n718 = n463 & n464 ;
  assign n3634 = n463 | n464 ;
  assign n5654 = ~n718 ;
  assign n3635 = n5654 & n3634 ;
  assign n3636 = n462 & n3635 ;
  assign n3637 = n462 | n3635 ;
  assign n5655 = ~n3636 ;
  assign n3638 = n5655 & n3637 ;
  assign n719 = x16 & x45 ;
  assign n465 = x15 & x46 ;
  assign n466 = x17 & x44 ;
  assign n720 = n465 & n466 ;
  assign n3639 = n465 | n466 ;
  assign n5656 = ~n720 ;
  assign n3640 = n5656 & n3639 ;
  assign n5657 = ~n719 ;
  assign n3641 = n5657 & n3640 ;
  assign n5658 = ~n3640 ;
  assign n3642 = n719 & n5658 ;
  assign n3643 = n3641 | n3642 ;
  assign n3644 = n3638 | n3643 ;
  assign n3645 = n3638 & n3643 ;
  assign n5659 = ~n3645 ;
  assign n3646 = n3644 & n5659 ;
  assign n3647 = n3633 & n3646 ;
  assign n3648 = n3633 | n3646 ;
  assign n5660 = ~n3647 ;
  assign n3649 = n5660 & n3648 ;
  assign n3650 = n3449 & n3458 ;
  assign n3651 = n3457 | n3650 ;
  assign n3652 = n3477 & n3482 ;
  assign n3653 = n3475 | n3652 ;
  assign n3654 = n3651 | n3653 ;
  assign n3655 = n3651 & n3653 ;
  assign n5661 = ~n3655 ;
  assign n3656 = n3654 & n5661 ;
  assign n3657 = n3649 & n3656 ;
  assign n3658 = n3649 | n3656 ;
  assign n5662 = ~n3657 ;
  assign n3659 = n5662 & n3658 ;
  assign n5663 = ~n3508 ;
  assign n3660 = n3505 & n5663 ;
  assign n3661 = n3659 & n3660 ;
  assign n3662 = n3659 | n3660 ;
  assign n5664 = ~n3661 ;
  assign n3663 = n5664 & n3662 ;
  assign n5665 = ~n3632 ;
  assign n3664 = n5665 & n3663 ;
  assign n5666 = ~n3663 ;
  assign n3665 = n3632 & n5666 ;
  assign n3666 = n3664 | n3665 ;
  assign n3434 = n3415 & n3432 ;
  assign n3667 = n3428 & n3429 ;
  assign n3668 = n3434 | n3667 ;
  assign n5667 = ~n429 ;
  assign n3401 = n5667 & n3399 ;
  assign n5668 = ~n3401 ;
  assign n3669 = n3398 & n5668 ;
  assign n721 = x10 & x51 ;
  assign n467 = x9 & x52 ;
  assign n468 = x11 & x50 ;
  assign n722 = n467 & n468 ;
  assign n3670 = n467 | n468 ;
  assign n5669 = ~n722 ;
  assign n3671 = n5669 & n3670 ;
  assign n5670 = ~n721 ;
  assign n3672 = n5670 & n3671 ;
  assign n5671 = ~n3671 ;
  assign n3673 = n721 & n5671 ;
  assign n3674 = n3672 | n3673 ;
  assign n471 = x8 & x53 ;
  assign n469 = x6 & x55 ;
  assign n470 = x7 & x54 ;
  assign n723 = n469 & n470 ;
  assign n3675 = n469 | n470 ;
  assign n5672 = ~n723 ;
  assign n3676 = n5672 & n3675 ;
  assign n5673 = ~n3676 ;
  assign n3677 = n471 & n5673 ;
  assign n5674 = ~n471 ;
  assign n3678 = n5674 & n3676 ;
  assign n3679 = n3677 | n3678 ;
  assign n3680 = n3674 | n3679 ;
  assign n3681 = n3674 & n3679 ;
  assign n5675 = ~n3681 ;
  assign n3682 = n3680 & n5675 ;
  assign n3683 = n3669 & n3682 ;
  assign n3684 = n3669 | n3682 ;
  assign n5676 = ~n3683 ;
  assign n3685 = n5676 & n3684 ;
  assign n5677 = ~n3420 ;
  assign n3686 = n3418 & n5677 ;
  assign n5678 = ~n437 ;
  assign n3687 = n5678 & n3446 ;
  assign n5679 = ~n3687 ;
  assign n3688 = n3445 & n5679 ;
  assign n474 = x13 & x48 ;
  assign n472 = x14 & x47 ;
  assign n473 = x12 & x49 ;
  assign n724 = n472 & n473 ;
  assign n3689 = n472 | n473 ;
  assign n5680 = ~n724 ;
  assign n3690 = n5680 & n3689 ;
  assign n5681 = ~n3690 ;
  assign n3691 = n474 & n5681 ;
  assign n5682 = ~n474 ;
  assign n3692 = n5682 & n3690 ;
  assign n3693 = n3691 | n3692 ;
  assign n5683 = ~n3693 ;
  assign n3694 = n3688 & n5683 ;
  assign n5684 = ~n3688 ;
  assign n3695 = n5684 & n3693 ;
  assign n3696 = n3694 | n3695 ;
  assign n5685 = ~n3686 ;
  assign n3697 = n5685 & n3696 ;
  assign n5686 = ~n3696 ;
  assign n3698 = n3686 & n5686 ;
  assign n3699 = n3697 | n3698 ;
  assign n3700 = n3417 & n3422 ;
  assign n3701 = n3426 | n3700 ;
  assign n3702 = n3699 | n3701 ;
  assign n3703 = n3699 & n3701 ;
  assign n5687 = ~n3703 ;
  assign n3704 = n3702 & n5687 ;
  assign n3705 = n3685 & n3704 ;
  assign n3706 = n3685 | n3704 ;
  assign n5688 = ~n3705 ;
  assign n3707 = n5688 & n3706 ;
  assign n5689 = ~n3468 ;
  assign n3708 = n3465 & n5689 ;
  assign n3709 = n3707 & n3708 ;
  assign n3710 = n3707 | n3708 ;
  assign n5690 = ~n3709 ;
  assign n3711 = n5690 & n3710 ;
  assign n5691 = ~n3668 ;
  assign n3712 = n5691 & n3711 ;
  assign n5692 = ~n3711 ;
  assign n3713 = n3668 & n5692 ;
  assign n3714 = n3712 | n3713 ;
  assign n5693 = ~n3514 ;
  assign n3715 = n3511 & n5693 ;
  assign n5694 = ~n3714 ;
  assign n3716 = n5694 & n3715 ;
  assign n5695 = ~n3715 ;
  assign n3717 = n3714 & n5695 ;
  assign n3718 = n3716 | n3717 ;
  assign n5696 = ~n3666 ;
  assign n3719 = n5696 & n3718 ;
  assign n5697 = ~n3718 ;
  assign n3720 = n3666 & n5697 ;
  assign n3721 = n3719 | n3720 ;
  assign n3722 = n3404 | n3409 ;
  assign n5698 = ~n3413 ;
  assign n3723 = n5698 & n3722 ;
  assign n5699 = ~n432 ;
  assign n3724 = n5699 & n3406 ;
  assign n5700 = ~n3724 ;
  assign n3725 = n3405 & n5700 ;
  assign n5701 = ~n3537 ;
  assign n3726 = n3535 & n5701 ;
  assign n725 = x3 & x58 ;
  assign n475 = x4 & x57 ;
  assign n476 = x5 & x56 ;
  assign n726 = n475 & n476 ;
  assign n3727 = n475 | n476 ;
  assign n5702 = ~n726 ;
  assign n3728 = n5702 & n3727 ;
  assign n5703 = ~n725 ;
  assign n3729 = n5703 & n3728 ;
  assign n5704 = ~n3728 ;
  assign n3730 = n725 & n5704 ;
  assign n3731 = n3729 | n3730 ;
  assign n3732 = n3726 | n3731 ;
  assign n3733 = n3726 & n3731 ;
  assign n5705 = ~n3733 ;
  assign n3734 = n3732 & n5705 ;
  assign n5706 = ~n3725 ;
  assign n3735 = n5706 & n3734 ;
  assign n5707 = ~n3734 ;
  assign n3736 = n3725 & n5707 ;
  assign n3737 = n3735 | n3736 ;
  assign n3738 = n3541 | n3543 ;
  assign n3739 = n3737 | n3738 ;
  assign n3740 = n3737 & n3738 ;
  assign n5708 = ~n3740 ;
  assign n3741 = n3739 & n5708 ;
  assign n3742 = n3723 & n3741 ;
  assign n3743 = n3723 | n3741 ;
  assign n5709 = ~n3742 ;
  assign n3744 = n5709 & n3743 ;
  assign n3745 = n3545 | n3548 ;
  assign n5710 = ~n3531 ;
  assign n3746 = n5710 & n3551 ;
  assign n5711 = ~n3746 ;
  assign n3747 = n3745 & n5711 ;
  assign n477 = x2 & x61 ;
  assign n3748 = x2 | x61 ;
  assign n5712 = ~n477 ;
  assign n3749 = n5712 & n3748 ;
  assign n3750 = n428 & n3749 ;
  assign n727 = x0 & x61 ;
  assign n728 = x2 & x59 ;
  assign n3751 = n727 | n728 ;
  assign n3752 = n451 | n3751 ;
  assign n3753 = n451 & n3751 ;
  assign n3754 = n428 | n3753 ;
  assign n5713 = ~n3754 ;
  assign n3755 = n3752 & n5713 ;
  assign n3756 = n3750 | n3755 ;
  assign n5714 = ~n3756 ;
  assign n3757 = n3747 & n5714 ;
  assign n5715 = ~n3747 ;
  assign n3758 = n5715 & n3756 ;
  assign n3759 = n3757 | n3758 ;
  assign n3760 = n3744 & n3759 ;
  assign n3762 = n3744 | n3759 ;
  assign n5716 = ~n3760 ;
  assign n3763 = n5716 & n3762 ;
  assign n5717 = ~n3441 ;
  assign n3764 = n3439 & n5717 ;
  assign n5718 = ~n3560 ;
  assign n3765 = n3558 & n5718 ;
  assign n3766 = n3764 & n3765 ;
  assign n3767 = n3764 | n3765 ;
  assign n5719 = ~n3766 ;
  assign n3768 = n5719 & n3767 ;
  assign n5720 = ~n3763 ;
  assign n3769 = n5720 & n3768 ;
  assign n5721 = ~n3768 ;
  assign n3770 = n3763 & n5721 ;
  assign n3771 = n3769 | n3770 ;
  assign n3772 = n3443 & n3520 ;
  assign n3773 = n3519 | n3772 ;
  assign n3774 = n3771 | n3773 ;
  assign n3775 = n3771 & n3773 ;
  assign n5722 = ~n3775 ;
  assign n3776 = n3774 & n5722 ;
  assign n5723 = ~n3721 ;
  assign n3777 = n5723 & n3776 ;
  assign n5724 = ~n3776 ;
  assign n3778 = n3721 & n5724 ;
  assign n3779 = n3777 | n3778 ;
  assign n3780 = n3523 & n3573 ;
  assign n3781 = n3572 | n3780 ;
  assign n5725 = ~n3526 ;
  assign n3782 = n5725 & n3566 ;
  assign n5726 = ~n3782 ;
  assign n3783 = n3564 & n5726 ;
  assign n5727 = ~n3781 ;
  assign n3784 = n5727 & n3783 ;
  assign n5728 = ~n3783 ;
  assign n3785 = n3781 & n5728 ;
  assign n3786 = n3784 | n3785 ;
  assign n5729 = ~n3779 ;
  assign n3787 = n5729 & n3786 ;
  assign n5730 = ~n3786 ;
  assign n3789 = n3779 & n5730 ;
  assign n3790 = n3787 | n3789 ;
  assign n5731 = ~n3583 ;
  assign n3791 = n3581 & n5731 ;
  assign n3792 = n3790 & n3791 ;
  assign n3793 = n3790 | n3791 ;
  assign n5732 = ~n3792 ;
  assign n3794 = n5732 & n3793 ;
  assign n5733 = ~n3593 ;
  assign n3795 = n5733 & n3794 ;
  assign n5734 = ~n3794 ;
  assign n3796 = n3593 & n5734 ;
  assign n94 = n3795 | n3796 ;
  assign n5735 = ~n3795 ;
  assign n3798 = n3793 & n5735 ;
  assign n5736 = ~n3777 ;
  assign n3799 = n3774 & n5736 ;
  assign n3800 = n3714 | n3715 ;
  assign n5737 = ~n3719 ;
  assign n3801 = n5737 & n3800 ;
  assign n478 = x8 & x54 ;
  assign n479 = x7 & x55 ;
  assign n480 = x9 & x53 ;
  assign n729 = n479 & n480 ;
  assign n3802 = n479 | n480 ;
  assign n5738 = ~n729 ;
  assign n3803 = n5738 & n3802 ;
  assign n3804 = n478 & n3803 ;
  assign n3805 = n478 | n3803 ;
  assign n5739 = ~n3804 ;
  assign n3806 = n5739 & n3805 ;
  assign n5740 = ~n3672 ;
  assign n3807 = n3670 & n5740 ;
  assign n481 = x10 & x52 ;
  assign n482 = x11 & x51 ;
  assign n483 = x12 & x50 ;
  assign n730 = n482 & n483 ;
  assign n3808 = n482 | n483 ;
  assign n5741 = ~n730 ;
  assign n3809 = n5741 & n3808 ;
  assign n3810 = n481 & n3809 ;
  assign n3811 = n481 | n3809 ;
  assign n5742 = ~n3810 ;
  assign n3812 = n5742 & n3811 ;
  assign n3813 = n3807 & n3812 ;
  assign n3814 = n3807 | n3812 ;
  assign n5743 = ~n3813 ;
  assign n3815 = n5743 & n3814 ;
  assign n3816 = n3806 & n3815 ;
  assign n3817 = n3806 | n3815 ;
  assign n5744 = ~n3816 ;
  assign n3818 = n5744 & n3817 ;
  assign n5745 = ~n3692 ;
  assign n3819 = n3689 & n5745 ;
  assign n5746 = ~n3641 ;
  assign n3820 = n3639 & n5746 ;
  assign n484 = x13 & x49 ;
  assign n485 = x15 & x47 ;
  assign n731 = x14 & x48 ;
  assign n5747 = ~n731 ;
  assign n3821 = n485 & n5747 ;
  assign n5748 = ~n485 ;
  assign n3822 = n5748 & n731 ;
  assign n3823 = n3821 | n3822 ;
  assign n5749 = ~n3823 ;
  assign n3824 = n484 & n5749 ;
  assign n5750 = ~n484 ;
  assign n3825 = n5750 & n3823 ;
  assign n3826 = n3824 | n3825 ;
  assign n5751 = ~n3820 ;
  assign n3827 = n5751 & n3826 ;
  assign n5752 = ~n3826 ;
  assign n3828 = n3820 & n5752 ;
  assign n3829 = n3827 | n3828 ;
  assign n3830 = n3819 | n3829 ;
  assign n3831 = n3819 & n3829 ;
  assign n5753 = ~n3831 ;
  assign n3832 = n3830 & n5753 ;
  assign n3833 = n3688 | n3693 ;
  assign n5754 = ~n3697 ;
  assign n3834 = n5754 & n3833 ;
  assign n3835 = n3832 & n3834 ;
  assign n3836 = n3832 | n3834 ;
  assign n5755 = ~n3835 ;
  assign n3837 = n5755 & n3836 ;
  assign n3838 = n3818 & n3837 ;
  assign n3839 = n3818 | n3837 ;
  assign n5756 = ~n3838 ;
  assign n3840 = n5756 & n3839 ;
  assign n5757 = ~n3649 ;
  assign n3841 = n5757 & n3656 ;
  assign n5758 = ~n3841 ;
  assign n3842 = n3654 & n5758 ;
  assign n5759 = ~n3685 ;
  assign n3843 = n5759 & n3704 ;
  assign n5760 = ~n3843 ;
  assign n3844 = n3702 & n5760 ;
  assign n5761 = ~n3842 ;
  assign n3845 = n5761 & n3844 ;
  assign n5762 = ~n3844 ;
  assign n3846 = n3842 & n5762 ;
  assign n3847 = n3845 | n3846 ;
  assign n5763 = ~n3840 ;
  assign n3848 = n5763 & n3847 ;
  assign n5764 = ~n3847 ;
  assign n3849 = n3840 & n5764 ;
  assign n3850 = n3848 | n3849 ;
  assign n5765 = ~n3664 ;
  assign n3851 = n3662 & n5765 ;
  assign n3852 = n3850 & n3851 ;
  assign n3853 = n3850 | n3851 ;
  assign n5766 = ~n3852 ;
  assign n3854 = n5766 & n3853 ;
  assign n3855 = n3801 & n3854 ;
  assign n3856 = n3801 | n3854 ;
  assign n5767 = ~n3855 ;
  assign n3857 = n5767 & n3856 ;
  assign n5768 = ~n3857 ;
  assign n3858 = n3799 & n5768 ;
  assign n5769 = ~n3799 ;
  assign n3859 = n5769 & n3857 ;
  assign n3860 = n3858 | n3859 ;
  assign n3861 = n3798 & n3860 ;
  assign n3862 = n3798 | n3860 ;
  assign n5770 = ~n3861 ;
  assign n3863 = n5770 & n3862 ;
  assign n3788 = n3779 & n3786 ;
  assign n3864 = n3781 & n3783 ;
  assign n3865 = n3788 | n3864 ;
  assign n3866 = n3740 | n3742 ;
  assign n489 = x0 & x62 ;
  assign n486 = x1 & x61 ;
  assign n487 = x3 & x59 ;
  assign n488 = x2 & x60 ;
  assign n732 = n487 & n488 ;
  assign n3867 = n487 | n488 ;
  assign n5771 = ~n732 ;
  assign n3868 = n5771 & n3867 ;
  assign n3869 = n486 & n3868 ;
  assign n3870 = n486 | n3868 ;
  assign n5772 = ~n3869 ;
  assign n3871 = n5772 & n3870 ;
  assign n733 = n428 & n477 ;
  assign n3872 = n733 | n3753 ;
  assign n5773 = ~n3872 ;
  assign n3873 = n3871 & n5773 ;
  assign n5774 = ~n3871 ;
  assign n3874 = n5774 & n3872 ;
  assign n3875 = n3873 | n3874 ;
  assign n3876 = n489 & n3875 ;
  assign n3877 = n489 | n3875 ;
  assign n5775 = ~n3876 ;
  assign n3878 = n5775 & n3877 ;
  assign n5776 = ~n3749 ;
  assign n3879 = n452 & n5776 ;
  assign n3880 = n3878 | n3879 ;
  assign n3881 = n3878 & n3879 ;
  assign n5777 = ~n3881 ;
  assign n3882 = n3880 & n5777 ;
  assign n5778 = ~n3866 ;
  assign n3883 = n5778 & n3882 ;
  assign n5779 = ~n3882 ;
  assign n3884 = n3866 & n5779 ;
  assign n3885 = n3883 | n3884 ;
  assign n5780 = ~n3712 ;
  assign n3886 = n3710 & n5780 ;
  assign n5781 = ~n3744 ;
  assign n3761 = n5781 & n3759 ;
  assign n3887 = n3747 | n3756 ;
  assign n5782 = ~n3761 ;
  assign n3888 = n5782 & n3887 ;
  assign n5783 = ~n3678 ;
  assign n3889 = n3675 & n5783 ;
  assign n5784 = ~n3729 ;
  assign n3890 = n3727 & n5784 ;
  assign n3891 = n3889 & n3890 ;
  assign n3892 = n3889 | n3890 ;
  assign n5785 = ~n3891 ;
  assign n3893 = n5785 & n3892 ;
  assign n492 = x4 & x58 ;
  assign n490 = x5 & x57 ;
  assign n491 = x6 & x56 ;
  assign n734 = n490 & n491 ;
  assign n3894 = n490 | n491 ;
  assign n5786 = ~n734 ;
  assign n3895 = n5786 & n3894 ;
  assign n3896 = n492 & n3895 ;
  assign n3897 = n492 | n3895 ;
  assign n5787 = ~n3896 ;
  assign n3898 = n5787 & n3897 ;
  assign n5788 = ~n3898 ;
  assign n3899 = n3893 & n5788 ;
  assign n5789 = ~n3893 ;
  assign n3900 = n5789 & n3898 ;
  assign n3901 = n3899 | n3900 ;
  assign n3902 = n3681 | n3683 ;
  assign n3903 = n3725 & n3734 ;
  assign n3904 = n3733 | n3903 ;
  assign n5790 = ~n3904 ;
  assign n3905 = n3902 & n5790 ;
  assign n5791 = ~n3902 ;
  assign n3906 = n5791 & n3904 ;
  assign n3907 = n3905 | n3906 ;
  assign n5792 = ~n3901 ;
  assign n3908 = n5792 & n3907 ;
  assign n5793 = ~n3907 ;
  assign n3909 = n3901 & n5793 ;
  assign n3910 = n3908 | n3909 ;
  assign n5794 = ~n3910 ;
  assign n3911 = n3888 & n5794 ;
  assign n5795 = ~n3888 ;
  assign n3912 = n5795 & n3910 ;
  assign n3913 = n3911 | n3912 ;
  assign n3914 = n3886 & n3913 ;
  assign n3915 = n3886 | n3913 ;
  assign n5796 = ~n3914 ;
  assign n3916 = n5796 & n3915 ;
  assign n3917 = n3885 & n3916 ;
  assign n3918 = n3885 | n3916 ;
  assign n5797 = ~n3917 ;
  assign n3919 = n5797 & n3918 ;
  assign n5798 = ~n3769 ;
  assign n3920 = n3767 & n5798 ;
  assign n493 = x27 & x35 ;
  assign n494 = x30 & x32 ;
  assign n735 = x29 & x33 ;
  assign n5799 = ~n735 ;
  assign n3921 = n494 & n5799 ;
  assign n5800 = ~n494 ;
  assign n3922 = n5800 & n735 ;
  assign n3923 = n3921 | n3922 ;
  assign n5801 = ~n3923 ;
  assign n3924 = n493 & n5801 ;
  assign n5802 = ~n493 ;
  assign n3925 = n5802 & n3923 ;
  assign n3926 = n3924 | n3925 ;
  assign n5803 = ~n453 ;
  assign n3927 = n5803 & n3595 ;
  assign n5804 = ~n3927 ;
  assign n3928 = n3594 & n5804 ;
  assign n5805 = ~n3928 ;
  assign n3929 = n3926 & n5805 ;
  assign n5806 = ~n3926 ;
  assign n3930 = n5806 & n3928 ;
  assign n3931 = n3929 | n3930 ;
  assign n736 = x26 & x36 ;
  assign n495 = x25 & x37 ;
  assign n496 = x28 & x34 ;
  assign n737 = n495 & n496 ;
  assign n3932 = n495 | n496 ;
  assign n5807 = ~n737 ;
  assign n3933 = n5807 & n3932 ;
  assign n5808 = ~n736 ;
  assign n3934 = n5808 & n3933 ;
  assign n5809 = ~n3933 ;
  assign n3935 = n736 & n5809 ;
  assign n3936 = n3934 | n3935 ;
  assign n5810 = ~n3936 ;
  assign n3937 = n3931 & n5810 ;
  assign n5811 = ~n3931 ;
  assign n3938 = n5811 & n3936 ;
  assign n3939 = n3937 | n3938 ;
  assign n5812 = ~n3606 ;
  assign n3940 = n3603 & n5812 ;
  assign n5813 = ~n3617 ;
  assign n3941 = n3614 & n5813 ;
  assign n5814 = ~n3941 ;
  assign n3942 = n3940 & n5814 ;
  assign n5815 = ~n3940 ;
  assign n3943 = n5815 & n3941 ;
  assign n3944 = n3942 | n3943 ;
  assign n499 = x22 & x40 ;
  assign n497 = x23 & x39 ;
  assign n498 = x24 & x38 ;
  assign n738 = n497 & n498 ;
  assign n3945 = n497 | n498 ;
  assign n5816 = ~n738 ;
  assign n3946 = n5816 & n3945 ;
  assign n5817 = ~n3946 ;
  assign n3947 = n499 & n5817 ;
  assign n5818 = ~n499 ;
  assign n3948 = n5818 & n3946 ;
  assign n3949 = n3947 | n3948 ;
  assign n3950 = n3944 & n3949 ;
  assign n3951 = n3944 | n3949 ;
  assign n5819 = ~n3950 ;
  assign n3952 = n5819 & n3951 ;
  assign n3953 = n3598 | n3599 ;
  assign n5820 = ~n3608 ;
  assign n3954 = n5820 & n3953 ;
  assign n3955 = n3952 & n3954 ;
  assign n3956 = n3952 | n3954 ;
  assign n5821 = ~n3955 ;
  assign n3957 = n5821 & n3956 ;
  assign n3958 = n3939 & n3957 ;
  assign n3959 = n3939 | n3957 ;
  assign n5822 = ~n3958 ;
  assign n3960 = n5822 & n3959 ;
  assign n3961 = n3645 | n3647 ;
  assign n500 = x21 & x41 ;
  assign n501 = x19 & x43 ;
  assign n739 = x20 & x42 ;
  assign n5823 = ~n739 ;
  assign n3962 = n501 & n5823 ;
  assign n5824 = ~n501 ;
  assign n3963 = n5824 & n739 ;
  assign n3964 = n3962 | n3963 ;
  assign n5825 = ~n3964 ;
  assign n3965 = n500 & n5825 ;
  assign n5826 = ~n500 ;
  assign n3966 = n5826 & n3964 ;
  assign n3967 = n3965 | n3966 ;
  assign n5827 = ~n462 ;
  assign n3968 = n5827 & n3635 ;
  assign n5828 = ~n3968 ;
  assign n3969 = n3634 & n5828 ;
  assign n504 = x16 & x46 ;
  assign n502 = x17 & x45 ;
  assign n503 = x18 & x44 ;
  assign n740 = n502 & n503 ;
  assign n3970 = n502 | n503 ;
  assign n5829 = ~n740 ;
  assign n3971 = n5829 & n3970 ;
  assign n3972 = n504 & n3971 ;
  assign n3973 = n504 | n3971 ;
  assign n5830 = ~n3972 ;
  assign n3974 = n5830 & n3973 ;
  assign n3975 = n3969 | n3974 ;
  assign n3976 = n3969 & n3974 ;
  assign n5831 = ~n3976 ;
  assign n3977 = n3975 & n5831 ;
  assign n5832 = ~n3967 ;
  assign n3978 = n5832 & n3977 ;
  assign n5833 = ~n3977 ;
  assign n3979 = n3967 & n5833 ;
  assign n3980 = n3978 | n3979 ;
  assign n3981 = n3611 & n3621 ;
  assign n3982 = n3620 | n3981 ;
  assign n3983 = n3980 | n3982 ;
  assign n3984 = n3980 & n3982 ;
  assign n5834 = ~n3984 ;
  assign n3985 = n3983 & n5834 ;
  assign n5835 = ~n3961 ;
  assign n3986 = n5835 & n3985 ;
  assign n5836 = ~n3985 ;
  assign n3987 = n3961 & n5836 ;
  assign n3988 = n3986 | n3987 ;
  assign n3989 = n3628 | n3630 ;
  assign n3990 = n3988 | n3989 ;
  assign n3991 = n3988 & n3989 ;
  assign n5837 = ~n3991 ;
  assign n3992 = n3990 & n5837 ;
  assign n5838 = ~n3960 ;
  assign n3993 = n5838 & n3992 ;
  assign n5839 = ~n3992 ;
  assign n3994 = n3960 & n5839 ;
  assign n3995 = n3993 | n3994 ;
  assign n3996 = n3920 & n3995 ;
  assign n3997 = n3920 | n3995 ;
  assign n5840 = ~n3996 ;
  assign n3998 = n5840 & n3997 ;
  assign n3999 = n3919 & n3998 ;
  assign n4000 = n3919 | n3998 ;
  assign n5841 = ~n3999 ;
  assign n4001 = n5841 & n4000 ;
  assign n5842 = ~n3865 ;
  assign n4002 = n5842 & n4001 ;
  assign n5843 = ~n4001 ;
  assign n4003 = n3865 & n5843 ;
  assign n4004 = n4002 | n4003 ;
  assign n4005 = n3863 | n4004 ;
  assign n4006 = n3863 & n4004 ;
  assign n5844 = ~n4006 ;
  assign n95 = n4005 & n5844 ;
  assign n4008 = n3865 & n4001 ;
  assign n4009 = n4006 | n4008 ;
  assign n741 = x15 & x48 ;
  assign n4010 = n484 & n3823 ;
  assign n5845 = ~n741 ;
  assign n4011 = n5845 & n4010 ;
  assign n4012 = n472 | n4010 ;
  assign n5846 = ~n4012 ;
  assign n4013 = n741 & n5846 ;
  assign n4014 = n4011 | n4013 ;
  assign n505 = x26 & x37 ;
  assign n4015 = n3842 & n3844 ;
  assign n4016 = n3840 & n3847 ;
  assign n4017 = n4015 | n4016 ;
  assign n4018 = n505 & n4017 ;
  assign n4019 = n505 | n4017 ;
  assign n5847 = ~n4018 ;
  assign n4020 = n5847 & n4019 ;
  assign n4021 = n4014 & n4020 ;
  assign n4022 = n4014 | n4020 ;
  assign n5848 = ~n4021 ;
  assign n4023 = n5848 & n4022 ;
  assign n506 = x9 & x54 ;
  assign n507 = x10 & x53 ;
  assign n742 = n506 & n507 ;
  assign n4024 = n506 | n507 ;
  assign n5849 = ~n742 ;
  assign n4025 = n5849 & n4024 ;
  assign n508 = x25 & x38 ;
  assign n509 = x8 & x55 ;
  assign n510 = x16 & x47 ;
  assign n743 = n509 & n510 ;
  assign n4026 = n509 | n510 ;
  assign n5850 = ~n743 ;
  assign n4027 = n5850 & n4026 ;
  assign n4028 = n452 & n3878 ;
  assign n5851 = ~n4028 ;
  assign n4029 = n477 & n5851 ;
  assign n5852 = ~n3748 ;
  assign n4030 = n5852 & n4028 ;
  assign n4031 = n4029 | n4030 ;
  assign n4032 = n4027 & n4031 ;
  assign n4033 = n4027 | n4031 ;
  assign n5853 = ~n4032 ;
  assign n4034 = n5853 & n4033 ;
  assign n4035 = n508 & n4034 ;
  assign n4036 = n508 | n4034 ;
  assign n5854 = ~n4035 ;
  assign n4037 = n5854 & n4036 ;
  assign n4038 = n4025 & n4037 ;
  assign n4039 = n4025 | n4037 ;
  assign n5855 = ~n4038 ;
  assign n4040 = n5855 & n4039 ;
  assign n4041 = n4023 & n4040 ;
  assign n4042 = n4023 | n4040 ;
  assign n5856 = ~n4041 ;
  assign n4043 = n5856 & n4042 ;
  assign n511 = x29 & x34 ;
  assign n4044 = n3940 | n3941 ;
  assign n5857 = ~n3949 ;
  assign n4045 = n3944 & n5857 ;
  assign n5858 = ~n4045 ;
  assign n4046 = n4044 & n5858 ;
  assign n4047 = n511 & n4046 ;
  assign n4048 = n511 | n4046 ;
  assign n5859 = ~n4047 ;
  assign n4049 = n5859 & n4048 ;
  assign n4050 = n730 | n3810 ;
  assign n4051 = n3960 & n3992 ;
  assign n4052 = n3991 | n4051 ;
  assign n744 = x12 & x51 ;
  assign n745 = x20 & x43 ;
  assign n4053 = n500 & n3964 ;
  assign n5860 = ~n745 ;
  assign n4054 = n5860 & n4053 ;
  assign n4055 = n463 | n4053 ;
  assign n5861 = ~n4055 ;
  assign n4056 = n745 & n5861 ;
  assign n4057 = n4054 | n4056 ;
  assign n5862 = ~n744 ;
  assign n4058 = n5862 & n4057 ;
  assign n5863 = ~n4057 ;
  assign n4059 = n744 & n5863 ;
  assign n4060 = n4058 | n4059 ;
  assign n5864 = ~n4060 ;
  assign n4061 = n4052 & n5864 ;
  assign n5865 = ~n4052 ;
  assign n4062 = n5865 & n4060 ;
  assign n4063 = n4061 | n4062 ;
  assign n512 = x7 & x56 ;
  assign n4064 = n3820 & n3826 ;
  assign n4065 = n3831 | n4064 ;
  assign n4066 = n3926 & n3928 ;
  assign n4067 = n3931 & n3936 ;
  assign n4068 = n4066 | n4067 ;
  assign n5866 = ~n4068 ;
  assign n4069 = n4065 & n5866 ;
  assign n5867 = ~n4065 ;
  assign n4070 = n5867 & n4068 ;
  assign n4071 = n4069 | n4070 ;
  assign n5868 = ~n4071 ;
  assign n4072 = n512 & n5868 ;
  assign n5869 = ~n512 ;
  assign n4073 = n5869 & n4071 ;
  assign n4074 = n4072 | n4073 ;
  assign n513 = x4 & x59 ;
  assign n746 = x21 & x42 ;
  assign n5870 = ~n746 ;
  assign n4075 = n513 & n5870 ;
  assign n5871 = ~n513 ;
  assign n4076 = n5871 & n746 ;
  assign n4077 = n4075 | n4076 ;
  assign n747 = x30 & x33 ;
  assign n4078 = n493 & n3923 ;
  assign n5872 = ~n747 ;
  assign n4079 = n5872 & n4078 ;
  assign n4080 = n455 | n4078 ;
  assign n5873 = ~n4080 ;
  assign n4081 = n747 & n5873 ;
  assign n4082 = n4079 | n4081 ;
  assign n5874 = ~n4077 ;
  assign n4083 = n5874 & n4082 ;
  assign n5875 = ~n4082 ;
  assign n4084 = n4077 & n5875 ;
  assign n4085 = n4083 | n4084 ;
  assign n514 = x19 & x44 ;
  assign n4086 = n499 & n3946 ;
  assign n5876 = ~n4086 ;
  assign n4087 = n514 & n5876 ;
  assign n5877 = ~n514 ;
  assign n4088 = n5877 & n4086 ;
  assign n4089 = n4087 | n4088 ;
  assign n4090 = n4085 | n4089 ;
  assign n4091 = n4085 & n4089 ;
  assign n5878 = ~n4091 ;
  assign n4092 = n4090 & n5878 ;
  assign n5879 = ~n4074 ;
  assign n4093 = n5879 & n4092 ;
  assign n5880 = ~n4092 ;
  assign n4094 = n4074 & n5880 ;
  assign n4095 = n4093 | n4094 ;
  assign n4096 = n3902 | n3904 ;
  assign n5881 = ~n3908 ;
  assign n4097 = n5881 & n4096 ;
  assign n515 = x28 & x35 ;
  assign n748 = x14 & x49 ;
  assign n5882 = ~n748 ;
  assign n4098 = n515 & n5882 ;
  assign n5883 = ~n515 ;
  assign n4099 = n5883 & n748 ;
  assign n4100 = n4098 | n4099 ;
  assign n4101 = n4097 | n4100 ;
  assign n4102 = n4097 & n4100 ;
  assign n5884 = ~n4102 ;
  assign n4103 = n4101 & n5884 ;
  assign n5885 = ~n4095 ;
  assign n4104 = n5885 & n4103 ;
  assign n5886 = ~n4103 ;
  assign n4105 = n4095 & n5886 ;
  assign n4106 = n4104 | n4105 ;
  assign n4107 = n4063 | n4106 ;
  assign n4108 = n4063 & n4106 ;
  assign n5887 = ~n4108 ;
  assign n4109 = n4107 & n5887 ;
  assign n4110 = n4050 & n4109 ;
  assign n4111 = n4050 | n4109 ;
  assign n5888 = ~n4110 ;
  assign n4112 = n5888 & n4111 ;
  assign n4113 = n4049 & n4112 ;
  assign n4114 = n4049 | n4112 ;
  assign n5889 = ~n4113 ;
  assign n4115 = n5889 & n4114 ;
  assign n4116 = n4043 & n4115 ;
  assign n4117 = n4043 | n4115 ;
  assign n5890 = ~n4116 ;
  assign n4118 = n5890 & n4117 ;
  assign n5891 = ~n478 ;
  assign n4119 = n5891 & n3803 ;
  assign n5892 = ~n4119 ;
  assign n4120 = n3802 & n5892 ;
  assign n5893 = ~n504 ;
  assign n4121 = n5893 & n3971 ;
  assign n5894 = ~n4121 ;
  assign n4122 = n3970 & n5894 ;
  assign n5895 = ~n4120 ;
  assign n4123 = n5895 & n4122 ;
  assign n5896 = ~n4122 ;
  assign n4124 = n4120 & n5896 ;
  assign n4125 = n4123 | n4124 ;
  assign n5897 = ~n4125 ;
  assign n4126 = n4118 & n5897 ;
  assign n5898 = ~n4118 ;
  assign n4127 = n5898 & n4125 ;
  assign n4128 = n4126 | n4127 ;
  assign n5899 = ~n4128 ;
  assign n4129 = n4009 & n5899 ;
  assign n5900 = ~n4009 ;
  assign n4130 = n5900 & n4128 ;
  assign n4131 = n4129 | n4130 ;
  assign n4132 = n3996 | n3999 ;
  assign n4133 = n3799 & n3857 ;
  assign n4134 = n3861 | n4133 ;
  assign n4135 = n4132 | n4134 ;
  assign n4136 = n4132 & n4134 ;
  assign n5901 = ~n4136 ;
  assign n4137 = n4135 & n5901 ;
  assign n5902 = ~n3801 ;
  assign n4138 = n5902 & n3854 ;
  assign n5903 = ~n4138 ;
  assign n4139 = n3853 & n5903 ;
  assign n4140 = n3888 & n3910 ;
  assign n4141 = n3914 | n4140 ;
  assign n4142 = n3866 | n3882 ;
  assign n5904 = ~n3916 ;
  assign n4143 = n3885 & n5904 ;
  assign n5905 = ~n4143 ;
  assign n4144 = n4142 & n5905 ;
  assign n5906 = ~n4141 ;
  assign n4145 = n5906 & n4144 ;
  assign n5907 = ~n4144 ;
  assign n4146 = n4141 & n5907 ;
  assign n4147 = n4145 | n4146 ;
  assign n5908 = ~n486 ;
  assign n4148 = n5908 & n3868 ;
  assign n5909 = ~n4148 ;
  assign n4149 = n3867 & n5909 ;
  assign n516 = x0 & x63 ;
  assign n749 = x11 & x52 ;
  assign n5910 = ~n749 ;
  assign n4150 = n516 & n5910 ;
  assign n5911 = ~n516 ;
  assign n4151 = n5911 & n749 ;
  assign n4152 = n4150 | n4151 ;
  assign n517 = x13 & x50 ;
  assign n750 = x5 & x58 ;
  assign n5912 = ~n750 ;
  assign n4153 = n517 & n5912 ;
  assign n5913 = ~n517 ;
  assign n4154 = n5913 & n750 ;
  assign n4155 = n4153 | n4154 ;
  assign n4156 = n4152 | n4155 ;
  assign n4157 = n4152 & n4155 ;
  assign n5914 = ~n4157 ;
  assign n4158 = n4156 & n5914 ;
  assign n518 = x17 & x46 ;
  assign n5915 = ~n3978 ;
  assign n4159 = n3975 & n5915 ;
  assign n4160 = n518 & n4159 ;
  assign n4161 = n518 | n4159 ;
  assign n5916 = ~n4160 ;
  assign n4162 = n5916 & n4161 ;
  assign n519 = x22 & x41 ;
  assign n5917 = ~n3986 ;
  assign n4163 = n3983 & n5917 ;
  assign n4164 = n519 & n4163 ;
  assign n4165 = n519 | n4163 ;
  assign n5918 = ~n4164 ;
  assign n4166 = n5918 & n4165 ;
  assign n5919 = ~n3934 ;
  assign n4167 = n3932 & n5919 ;
  assign n4168 = n4166 & n4167 ;
  assign n4169 = n4166 | n4167 ;
  assign n5920 = ~n4168 ;
  assign n4170 = n5920 & n4169 ;
  assign n4171 = n4162 & n4170 ;
  assign n4172 = n4162 | n4170 ;
  assign n5921 = ~n4171 ;
  assign n4173 = n5921 & n4172 ;
  assign n521 = x1 & x62 ;
  assign n520 = x23 & x40 ;
  assign n4174 = n3893 & n3898 ;
  assign n4175 = n3891 | n4174 ;
  assign n5922 = ~n4175 ;
  assign n4176 = n520 & n5922 ;
  assign n5923 = ~n520 ;
  assign n4177 = n5923 & n4175 ;
  assign n4178 = n4176 | n4177 ;
  assign n5924 = ~n4178 ;
  assign n4179 = n521 & n5924 ;
  assign n5925 = ~n521 ;
  assign n4180 = n5925 & n4178 ;
  assign n4181 = n4179 | n4180 ;
  assign n5926 = ~n4181 ;
  assign n4182 = n4173 & n5926 ;
  assign n5927 = ~n4173 ;
  assign n4183 = n5927 & n4181 ;
  assign n4184 = n4182 | n4183 ;
  assign n5928 = ~n4184 ;
  assign n4185 = n4158 & n5928 ;
  assign n5929 = ~n4158 ;
  assign n4186 = n5929 & n4184 ;
  assign n4187 = n4185 | n4186 ;
  assign n751 = x6 & x57 ;
  assign n4188 = n3813 | n3816 ;
  assign n4189 = n751 | n4188 ;
  assign n4190 = n751 & n4188 ;
  assign n5930 = ~n4190 ;
  assign n4191 = n4189 & n5930 ;
  assign n5931 = ~n4187 ;
  assign n4192 = n5931 & n4191 ;
  assign n5932 = ~n4191 ;
  assign n4193 = n4187 & n5932 ;
  assign n4194 = n4192 | n4193 ;
  assign n522 = x3 & x60 ;
  assign n752 = x18 & x45 ;
  assign n4195 = n3871 | n3872 ;
  assign n5933 = ~n489 ;
  assign n4196 = n5933 & n3875 ;
  assign n5934 = ~n4196 ;
  assign n4197 = n4195 & n5934 ;
  assign n5935 = ~n752 ;
  assign n4198 = n5935 & n4197 ;
  assign n5936 = ~n4197 ;
  assign n4199 = n752 & n5936 ;
  assign n4200 = n4198 | n4199 ;
  assign n5937 = ~n4200 ;
  assign n4201 = n522 & n5937 ;
  assign n5938 = ~n522 ;
  assign n4202 = n5938 & n4200 ;
  assign n4203 = n4201 | n4202 ;
  assign n5939 = ~n3818 ;
  assign n4204 = n5939 & n3837 ;
  assign n5940 = ~n4204 ;
  assign n4205 = n3836 & n5940 ;
  assign n523 = x31 & x32 ;
  assign n524 = x24 & x39 ;
  assign n5941 = ~n460 ;
  assign n4206 = n5941 & n524 ;
  assign n4207 = n523 & n4206 ;
  assign n4208 = n523 | n4206 ;
  assign n5942 = ~n4207 ;
  assign n4209 = n5942 & n4208 ;
  assign n5943 = ~n492 ;
  assign n4210 = n5943 & n3895 ;
  assign n5944 = ~n4210 ;
  assign n4211 = n3894 & n5944 ;
  assign n4212 = n4209 & n4211 ;
  assign n4213 = n4209 | n4211 ;
  assign n5945 = ~n4212 ;
  assign n4214 = n5945 & n4213 ;
  assign n5946 = ~n4205 ;
  assign n4215 = n5946 & n4214 ;
  assign n5947 = ~n4214 ;
  assign n4216 = n4205 & n5947 ;
  assign n4217 = n4215 | n4216 ;
  assign n4218 = n4203 | n4217 ;
  assign n4219 = n4203 & n4217 ;
  assign n5948 = ~n4219 ;
  assign n4220 = n4218 & n5948 ;
  assign n525 = x27 & x36 ;
  assign n5949 = ~n3939 ;
  assign n4221 = n5949 & n3957 ;
  assign n5950 = ~n4221 ;
  assign n4222 = n3956 & n5950 ;
  assign n5951 = ~n4222 ;
  assign n4223 = n525 & n5951 ;
  assign n5952 = ~n525 ;
  assign n4224 = n5952 & n4222 ;
  assign n4225 = n4223 | n4224 ;
  assign n5953 = ~n4225 ;
  assign n4226 = n4220 & n5953 ;
  assign n5954 = ~n4220 ;
  assign n4227 = n5954 & n4225 ;
  assign n4228 = n4226 | n4227 ;
  assign n4229 = n4194 | n4228 ;
  assign n4230 = n4194 & n4228 ;
  assign n5955 = ~n4230 ;
  assign n4231 = n4229 & n5955 ;
  assign n5956 = ~n4149 ;
  assign n4232 = n5956 & n4231 ;
  assign n5957 = ~n4231 ;
  assign n4233 = n4149 & n5957 ;
  assign n4234 = n4232 | n4233 ;
  assign n4235 = n4147 | n4234 ;
  assign n4236 = n4147 & n4234 ;
  assign n5958 = ~n4236 ;
  assign n4237 = n4235 & n5958 ;
  assign n5959 = ~n4139 ;
  assign n4238 = n5959 & n4237 ;
  assign n5960 = ~n4237 ;
  assign n4239 = n4139 & n5960 ;
  assign n4240 = n4238 | n4239 ;
  assign n5961 = ~n4240 ;
  assign n4241 = n4137 & n5961 ;
  assign n5962 = ~n4137 ;
  assign n4242 = n5962 & n4240 ;
  assign n4243 = n4241 | n4242 ;
  assign n4244 = n4131 | n4243 ;
  assign n4245 = n4131 & n4243 ;
  assign n5963 = ~n4245 ;
  assign n96 = n4244 & n5963 ;
  assign y0 = n65 ;
  assign y1 = n66 ;
  assign y2 = n67 ;
  assign y3 = n68 ;
  assign y4 = n69 ;
  assign y5 = n70 ;
  assign y6 = n71 ;
  assign y7 = n72 ;
  assign y8 = n73 ;
  assign y9 = n74 ;
  assign y10 = n75 ;
  assign y11 = n76 ;
  assign y12 = n77 ;
  assign y13 = n78 ;
  assign y14 = n79 ;
  assign y15 = n80 ;
  assign y16 = n81 ;
  assign y17 = n82 ;
  assign y18 = n83 ;
  assign y19 = n84 ;
  assign y20 = n85 ;
  assign y21 = n86 ;
  assign y22 = n87 ;
  assign y23 = n88 ;
  assign y24 = n89 ;
  assign y25 = n90 ;
  assign y26 = n91 ;
  assign y27 = n92 ;
  assign y28 = n93 ;
  assign y29 = n94 ;
  assign y30 = n95 ;
  assign y31 = n96 ;
endmodule
