module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 ;
  assign n4602 = x32 & x33 ;
  assign n4597 = ~x1 ;
  assign n109 = n4597 & n4602 ;
  assign n112 = x62 | x63 ;
  assign n113 = x61 | n112 ;
  assign n114 = x60 | n113 ;
  assign n115 = x59 | n114 ;
  assign n116 = x58 | n115 ;
  assign n117 = x57 | n116 ;
  assign n118 = x56 | n117 ;
  assign n119 = x55 | n118 ;
  assign n120 = x54 | n119 ;
  assign n121 = x53 | n120 ;
  assign n122 = x52 | n121 ;
  assign n123 = x51 | n122 ;
  assign n124 = x50 | n123 ;
  assign n125 = x49 | n124 ;
  assign n126 = x48 | n125 ;
  assign n127 = x47 | n126 ;
  assign n128 = x46 | n127 ;
  assign n129 = x45 | n128 ;
  assign n130 = x44 | n129 ;
  assign n131 = x43 | n130 ;
  assign n132 = x42 | n131 ;
  assign n133 = x41 | n132 ;
  assign n134 = x40 | n133 ;
  assign n135 = x39 | n134 ;
  assign n136 = x38 | n135 ;
  assign n137 = x35 | x36 ;
  assign n138 = x37 | n137 ;
  assign n139 = n136 | n138 ;
  assign n4598 = ~x30 ;
  assign n144 = n4598 & x32 ;
  assign n145 = x34 | n144 ;
  assign n146 = n139 | n145 ;
  assign n4599 = ~n146 ;
  assign n147 = x33 & n4599 ;
  assign n4600 = ~n147 ;
  assign n148 = x31 & n4600 ;
  assign n140 = x33 | x34 ;
  assign n4601 = ~x31 ;
  assign n141 = n4601 & x32 ;
  assign n142 = n140 | n141 ;
  assign n143 = n139 | n142 ;
  assign n96 = ~n143 ;
  assign n149 = x32 & n96 ;
  assign n4603 = ~n149 ;
  assign n150 = n148 & n4603 ;
  assign n4604 = ~x29 ;
  assign n4612 = n4604 & n4602 ;
  assign n151 = n4601 & x33 ;
  assign n152 = n146 | n151 ;
  assign n95 = ~n152 ;
  assign n153 = x32 & n95 ;
  assign n4606 = ~n153 ;
  assign n154 = x30 & n4606 ;
  assign n4605 = n4604 & x32 ;
  assign n155 = x33 | n4605 ;
  assign n4607 = ~n154 ;
  assign n156 = n4607 & n155 ;
  assign n157 = n4612 | n156 ;
  assign n158 = x34 | n157 ;
  assign n159 = x34 & n157 ;
  assign n160 = n139 | n159 ;
  assign n4608 = ~n160 ;
  assign n162 = n158 & n4608 ;
  assign n4609 = ~n162 ;
  assign n163 = n150 & n4609 ;
  assign n4610 = ~x28 ;
  assign n4622 = n4610 & n4602 ;
  assign n4611 = ~n150 ;
  assign n161 = n4611 & n158 ;
  assign n165 = n160 | n161 ;
  assign n94 = ~n165 ;
  assign n166 = x32 & n94 ;
  assign n167 = n4604 & n166 ;
  assign n4613 = ~n166 ;
  assign n168 = x29 & n4613 ;
  assign n169 = n167 | n168 ;
  assign n170 = n4610 & x32 ;
  assign n171 = x33 | n170 ;
  assign n4614 = ~n169 ;
  assign n172 = n4614 & n171 ;
  assign n173 = n4622 | n172 ;
  assign n175 = x34 & n173 ;
  assign n174 = x34 | n173 ;
  assign n4615 = ~n4612 ;
  assign n176 = n4615 & n155 ;
  assign n177 = n94 & n176 ;
  assign n178 = n4607 & n177 ;
  assign n4616 = ~n177 ;
  assign n179 = n154 & n4616 ;
  assign n180 = n178 | n179 ;
  assign n4617 = ~n180 ;
  assign n181 = n174 & n4617 ;
  assign n182 = n175 | n181 ;
  assign n183 = x35 | n182 ;
  assign n4618 = ~n163 ;
  assign n164 = x35 & n4618 ;
  assign n184 = x37 | n136 ;
  assign n185 = x36 | n184 ;
  assign n186 = n164 | n185 ;
  assign n187 = x35 & n182 ;
  assign n188 = n186 | n187 ;
  assign n4619 = ~n188 ;
  assign n189 = n183 & n4619 ;
  assign n4620 = ~n189 ;
  assign n190 = n163 & n4620 ;
  assign n4621 = ~x27 ;
  assign n4635 = n4621 & n4602 ;
  assign n191 = n4618 & n182 ;
  assign n192 = n188 | n191 ;
  assign n93 = ~n192 ;
  assign n193 = x32 & n93 ;
  assign n194 = n4610 & n193 ;
  assign n4623 = ~n193 ;
  assign n195 = x28 & n4623 ;
  assign n196 = n194 | n195 ;
  assign n197 = n4621 & x32 ;
  assign n198 = x33 | n197 ;
  assign n4624 = ~n196 ;
  assign n199 = n4624 & n198 ;
  assign n200 = n4635 | n199 ;
  assign n201 = x34 & n200 ;
  assign n4625 = ~n4622 ;
  assign n202 = n4625 & n171 ;
  assign n203 = n93 & n202 ;
  assign n204 = n4614 & n203 ;
  assign n4626 = ~n203 ;
  assign n205 = n169 & n4626 ;
  assign n206 = n204 | n205 ;
  assign n207 = x34 | n200 ;
  assign n4627 = ~n206 ;
  assign n208 = n4627 & n207 ;
  assign n209 = n201 | n208 ;
  assign n210 = x35 & n209 ;
  assign n211 = x35 | n209 ;
  assign n4628 = ~n175 ;
  assign n212 = n174 & n4628 ;
  assign n213 = n93 & n212 ;
  assign n214 = n4617 & n213 ;
  assign n4629 = ~n213 ;
  assign n215 = n180 & n4629 ;
  assign n216 = n214 | n215 ;
  assign n4630 = ~n216 ;
  assign n217 = n211 & n4630 ;
  assign n218 = n210 | n217 ;
  assign n219 = x36 | n218 ;
  assign n220 = x36 & n218 ;
  assign n221 = n184 | n220 ;
  assign n4631 = ~n221 ;
  assign n223 = n219 & n4631 ;
  assign n4632 = ~n223 ;
  assign n224 = n190 & n4632 ;
  assign n4633 = ~x26 ;
  assign n4650 = n4633 & n4602 ;
  assign n4634 = ~n190 ;
  assign n222 = n4634 & n219 ;
  assign n225 = n221 | n222 ;
  assign n92 = ~n225 ;
  assign n226 = x32 & n92 ;
  assign n227 = n4621 & n226 ;
  assign n4636 = ~n226 ;
  assign n228 = x27 & n4636 ;
  assign n229 = n227 | n228 ;
  assign n230 = n4633 & x32 ;
  assign n231 = x33 | n230 ;
  assign n4637 = ~n229 ;
  assign n232 = n4637 & n231 ;
  assign n233 = n4650 | n232 ;
  assign n234 = x34 & n233 ;
  assign n4638 = ~n4635 ;
  assign n235 = n4638 & n198 ;
  assign n236 = n92 & n235 ;
  assign n237 = n4624 & n236 ;
  assign n4639 = ~n236 ;
  assign n238 = n196 & n4639 ;
  assign n239 = n237 | n238 ;
  assign n240 = x34 | n233 ;
  assign n4640 = ~n239 ;
  assign n241 = n4640 & n240 ;
  assign n242 = n234 | n241 ;
  assign n243 = x35 & n242 ;
  assign n244 = x35 | n242 ;
  assign n4641 = ~n201 ;
  assign n245 = n4641 & n207 ;
  assign n246 = n92 & n245 ;
  assign n247 = n206 & n246 ;
  assign n248 = n206 | n246 ;
  assign n4642 = ~n247 ;
  assign n249 = n4642 & n248 ;
  assign n4643 = ~n249 ;
  assign n250 = n244 & n4643 ;
  assign n251 = n243 | n250 ;
  assign n252 = x36 & n251 ;
  assign n253 = x36 | n251 ;
  assign n4644 = ~n210 ;
  assign n254 = n4644 & n211 ;
  assign n255 = n92 & n254 ;
  assign n256 = n4630 & n255 ;
  assign n4645 = ~n255 ;
  assign n257 = n216 & n4645 ;
  assign n258 = n256 | n257 ;
  assign n4646 = ~n258 ;
  assign n259 = n253 & n4646 ;
  assign n260 = n252 | n259 ;
  assign n261 = x37 | n260 ;
  assign n262 = x37 & n260 ;
  assign n263 = n136 | n262 ;
  assign n4647 = ~n263 ;
  assign n265 = n261 & n4647 ;
  assign n4648 = ~n265 ;
  assign n266 = n224 & n4648 ;
  assign n4649 = ~n224 ;
  assign n264 = n4649 & n261 ;
  assign n267 = n263 | n264 ;
  assign n91 = ~n267 ;
  assign n268 = x32 & n91 ;
  assign n269 = n4633 & n268 ;
  assign n4651 = ~n268 ;
  assign n270 = x26 & n4651 ;
  assign n271 = n269 | n270 ;
  assign n4652 = ~x25 ;
  assign n4673 = n4652 & x32 ;
  assign n272 = x33 | n4673 ;
  assign n4653 = ~n271 ;
  assign n273 = n4653 & n272 ;
  assign n274 = n4652 & n4602 ;
  assign n275 = n273 | n274 ;
  assign n277 = x34 & n275 ;
  assign n276 = x34 | n275 ;
  assign n4654 = ~n4650 ;
  assign n278 = n4654 & n231 ;
  assign n279 = n91 & n278 ;
  assign n280 = n4637 & n279 ;
  assign n4655 = ~n279 ;
  assign n281 = n229 & n4655 ;
  assign n282 = n280 | n281 ;
  assign n4656 = ~n282 ;
  assign n283 = n276 & n4656 ;
  assign n284 = n277 | n283 ;
  assign n285 = x35 | n284 ;
  assign n286 = x35 & n284 ;
  assign n4657 = ~n234 ;
  assign n287 = n4657 & n240 ;
  assign n288 = n91 & n287 ;
  assign n4658 = ~n288 ;
  assign n289 = n239 & n4658 ;
  assign n290 = n4640 & n288 ;
  assign n291 = n289 | n290 ;
  assign n4659 = ~n286 ;
  assign n292 = n4659 & n291 ;
  assign n4660 = ~n292 ;
  assign n293 = n285 & n4660 ;
  assign n294 = x36 | n293 ;
  assign n295 = x36 & n293 ;
  assign n4661 = ~n243 ;
  assign n296 = n4661 & n244 ;
  assign n297 = n91 & n296 ;
  assign n298 = n249 & n297 ;
  assign n299 = n249 | n297 ;
  assign n4662 = ~n298 ;
  assign n300 = n4662 & n299 ;
  assign n4663 = ~n295 ;
  assign n301 = n4663 & n300 ;
  assign n4664 = ~n301 ;
  assign n302 = n294 & n4664 ;
  assign n303 = x37 | n302 ;
  assign n304 = x37 & n302 ;
  assign n4665 = ~n252 ;
  assign n305 = n4665 & n253 ;
  assign n306 = n91 & n305 ;
  assign n307 = n4646 & n306 ;
  assign n4666 = ~n306 ;
  assign n308 = n258 & n4666 ;
  assign n309 = n307 | n308 ;
  assign n4667 = ~n304 ;
  assign n310 = n4667 & n309 ;
  assign n4668 = ~n310 ;
  assign n311 = n303 & n4668 ;
  assign n312 = x38 | n311 ;
  assign n313 = x38 & n311 ;
  assign n314 = n135 | n313 ;
  assign n4669 = ~n314 ;
  assign n315 = n312 & n4669 ;
  assign n4670 = ~n315 ;
  assign n316 = n266 & n4670 ;
  assign n4671 = ~x24 ;
  assign n4695 = n4671 & n4602 ;
  assign n4672 = ~n266 ;
  assign n317 = n4672 & n312 ;
  assign n318 = n314 | n317 ;
  assign n90 = ~n318 ;
  assign n319 = x32 & n90 ;
  assign n320 = n4652 & n319 ;
  assign n4674 = ~n319 ;
  assign n321 = x25 & n4674 ;
  assign n322 = n320 | n321 ;
  assign n323 = n4671 & x32 ;
  assign n324 = x33 | n323 ;
  assign n4675 = ~n322 ;
  assign n325 = n4675 & n324 ;
  assign n326 = n4695 | n325 ;
  assign n327 = x34 & n326 ;
  assign n4676 = ~n274 ;
  assign n328 = n272 & n4676 ;
  assign n329 = n90 & n328 ;
  assign n330 = n4653 & n329 ;
  assign n4677 = ~n329 ;
  assign n331 = n271 & n4677 ;
  assign n332 = n330 | n331 ;
  assign n333 = x34 | n326 ;
  assign n4678 = ~n332 ;
  assign n334 = n4678 & n333 ;
  assign n335 = n327 | n334 ;
  assign n336 = x35 & n335 ;
  assign n337 = x35 | n335 ;
  assign n338 = n277 | n318 ;
  assign n4679 = ~n338 ;
  assign n339 = n276 & n4679 ;
  assign n4680 = ~n339 ;
  assign n340 = n282 & n4680 ;
  assign n341 = n283 & n4679 ;
  assign n342 = n340 | n341 ;
  assign n4681 = ~n342 ;
  assign n343 = n337 & n4681 ;
  assign n344 = n336 | n343 ;
  assign n345 = x36 & n344 ;
  assign n346 = x36 | n344 ;
  assign n347 = n285 & n4659 ;
  assign n348 = n90 & n347 ;
  assign n4682 = ~n291 ;
  assign n349 = n4682 & n348 ;
  assign n4683 = ~n348 ;
  assign n350 = n291 & n4683 ;
  assign n351 = n349 | n350 ;
  assign n4684 = ~n351 ;
  assign n352 = n346 & n4684 ;
  assign n353 = n345 | n352 ;
  assign n354 = x37 & n353 ;
  assign n355 = x37 | n353 ;
  assign n356 = n294 & n4663 ;
  assign n357 = n90 & n356 ;
  assign n4685 = ~n300 ;
  assign n358 = n4685 & n357 ;
  assign n4686 = ~n357 ;
  assign n359 = n300 & n4686 ;
  assign n360 = n358 | n359 ;
  assign n4687 = ~n360 ;
  assign n361 = n355 & n4687 ;
  assign n362 = n354 | n361 ;
  assign n363 = x38 & n362 ;
  assign n364 = x38 | n362 ;
  assign n365 = n303 & n4667 ;
  assign n366 = n90 & n365 ;
  assign n4688 = ~n309 ;
  assign n367 = n4688 & n366 ;
  assign n4689 = ~n366 ;
  assign n368 = n309 & n4689 ;
  assign n369 = n367 | n368 ;
  assign n4690 = ~n369 ;
  assign n370 = n364 & n4690 ;
  assign n371 = n363 | n370 ;
  assign n372 = x39 | n371 ;
  assign n373 = x39 & n371 ;
  assign n374 = n134 | n373 ;
  assign n4691 = ~n374 ;
  assign n376 = n372 & n4691 ;
  assign n4692 = ~n376 ;
  assign n377 = n316 & n4692 ;
  assign n4693 = ~x23 ;
  assign n4720 = n4693 & n4602 ;
  assign n4694 = ~n316 ;
  assign n375 = n4694 & n372 ;
  assign n378 = n374 | n375 ;
  assign n89 = ~n378 ;
  assign n379 = x32 & n89 ;
  assign n380 = n4671 & n379 ;
  assign n4696 = ~n379 ;
  assign n381 = x24 & n4696 ;
  assign n382 = n380 | n381 ;
  assign n383 = n4693 & x32 ;
  assign n384 = x33 | n383 ;
  assign n4697 = ~n382 ;
  assign n385 = n4697 & n384 ;
  assign n386 = n4720 | n385 ;
  assign n387 = x34 & n386 ;
  assign n4698 = ~n4695 ;
  assign n388 = n4698 & n324 ;
  assign n389 = n89 & n388 ;
  assign n390 = n4675 & n389 ;
  assign n4699 = ~n389 ;
  assign n391 = n322 & n4699 ;
  assign n392 = n390 | n391 ;
  assign n393 = x34 | n386 ;
  assign n4700 = ~n392 ;
  assign n394 = n4700 & n393 ;
  assign n395 = n387 | n394 ;
  assign n396 = x35 & n395 ;
  assign n397 = x35 | n395 ;
  assign n4701 = ~n327 ;
  assign n398 = n4701 & n333 ;
  assign n399 = n89 & n398 ;
  assign n400 = n332 & n399 ;
  assign n401 = n332 | n399 ;
  assign n4702 = ~n400 ;
  assign n402 = n4702 & n401 ;
  assign n4703 = ~n402 ;
  assign n403 = n397 & n4703 ;
  assign n404 = n396 | n403 ;
  assign n405 = x36 & n404 ;
  assign n406 = x36 | n404 ;
  assign n4704 = ~n336 ;
  assign n407 = n4704 & n337 ;
  assign n408 = n89 & n407 ;
  assign n409 = n342 & n408 ;
  assign n410 = n342 | n408 ;
  assign n4705 = ~n409 ;
  assign n411 = n4705 & n410 ;
  assign n4706 = ~n411 ;
  assign n412 = n406 & n4706 ;
  assign n413 = n405 | n412 ;
  assign n414 = x37 & n413 ;
  assign n415 = x37 | n413 ;
  assign n4707 = ~n345 ;
  assign n416 = n4707 & n346 ;
  assign n417 = n89 & n416 ;
  assign n418 = n4684 & n417 ;
  assign n4708 = ~n417 ;
  assign n419 = n351 & n4708 ;
  assign n420 = n418 | n419 ;
  assign n4709 = ~n420 ;
  assign n421 = n415 & n4709 ;
  assign n422 = n414 | n421 ;
  assign n423 = x38 & n422 ;
  assign n424 = x38 | n422 ;
  assign n4710 = ~n354 ;
  assign n425 = n4710 & n355 ;
  assign n426 = n89 & n425 ;
  assign n427 = n360 & n426 ;
  assign n428 = n360 | n426 ;
  assign n4711 = ~n427 ;
  assign n429 = n4711 & n428 ;
  assign n4712 = ~n429 ;
  assign n430 = n424 & n4712 ;
  assign n431 = n423 | n430 ;
  assign n432 = x39 & n431 ;
  assign n433 = x39 | n431 ;
  assign n4713 = ~n363 ;
  assign n434 = n4713 & n364 ;
  assign n435 = n89 & n434 ;
  assign n436 = n369 & n435 ;
  assign n437 = n369 | n435 ;
  assign n4714 = ~n436 ;
  assign n438 = n4714 & n437 ;
  assign n4715 = ~n438 ;
  assign n439 = n433 & n4715 ;
  assign n440 = n432 | n439 ;
  assign n441 = x40 | n440 ;
  assign n442 = x40 & n440 ;
  assign n443 = n133 | n442 ;
  assign n4716 = ~n443 ;
  assign n445 = n441 & n4716 ;
  assign n4717 = ~n445 ;
  assign n446 = n377 & n4717 ;
  assign n4718 = ~x22 ;
  assign n4783 = n4718 & n4602 ;
  assign n4719 = ~n377 ;
  assign n444 = n4719 & n441 ;
  assign n447 = n443 | n444 ;
  assign n88 = ~n447 ;
  assign n448 = x32 & n88 ;
  assign n449 = x23 & n448 ;
  assign n451 = x23 | n448 ;
  assign n4721 = ~n449 ;
  assign n452 = n4721 & n451 ;
  assign n4750 = n4718 & x32 ;
  assign n453 = x33 | n4750 ;
  assign n4722 = ~n452 ;
  assign n454 = n4722 & n453 ;
  assign n455 = n4783 | n454 ;
  assign n456 = x34 & n455 ;
  assign n450 = n4693 & n448 ;
  assign n4723 = ~n448 ;
  assign n457 = x23 & n4723 ;
  assign n458 = n450 | n457 ;
  assign n4724 = ~n458 ;
  assign n459 = n453 & n4724 ;
  assign n460 = n4783 | n459 ;
  assign n461 = x34 | n460 ;
  assign n4725 = ~n4720 ;
  assign n462 = n4725 & n384 ;
  assign n463 = n88 & n462 ;
  assign n464 = n4697 & n463 ;
  assign n4726 = ~n463 ;
  assign n465 = n382 & n4726 ;
  assign n466 = n464 | n465 ;
  assign n4727 = ~n466 ;
  assign n467 = n461 & n4727 ;
  assign n468 = n456 | n467 ;
  assign n469 = x35 & n468 ;
  assign n470 = x35 | n468 ;
  assign n4728 = ~n387 ;
  assign n471 = n4728 & n393 ;
  assign n472 = n88 & n471 ;
  assign n473 = n392 & n472 ;
  assign n474 = n392 | n472 ;
  assign n4729 = ~n473 ;
  assign n475 = n4729 & n474 ;
  assign n4730 = ~n475 ;
  assign n476 = n470 & n4730 ;
  assign n477 = n469 | n476 ;
  assign n478 = x36 & n477 ;
  assign n479 = x36 | n477 ;
  assign n4731 = ~n396 ;
  assign n480 = n4731 & n397 ;
  assign n481 = n88 & n480 ;
  assign n482 = n402 & n481 ;
  assign n483 = n402 | n481 ;
  assign n4732 = ~n482 ;
  assign n484 = n4732 & n483 ;
  assign n4733 = ~n484 ;
  assign n485 = n479 & n4733 ;
  assign n486 = n478 | n485 ;
  assign n487 = x37 & n486 ;
  assign n488 = x37 | n486 ;
  assign n4734 = ~n405 ;
  assign n489 = n4734 & n406 ;
  assign n490 = n88 & n489 ;
  assign n491 = n411 & n490 ;
  assign n492 = n411 | n490 ;
  assign n4735 = ~n491 ;
  assign n493 = n4735 & n492 ;
  assign n4736 = ~n493 ;
  assign n494 = n488 & n4736 ;
  assign n495 = n487 | n494 ;
  assign n496 = x38 & n495 ;
  assign n497 = x38 | n495 ;
  assign n4737 = ~n414 ;
  assign n498 = n4737 & n415 ;
  assign n499 = n88 & n498 ;
  assign n500 = n4709 & n499 ;
  assign n4738 = ~n499 ;
  assign n501 = n420 & n4738 ;
  assign n502 = n500 | n501 ;
  assign n4739 = ~n502 ;
  assign n503 = n497 & n4739 ;
  assign n504 = n496 | n503 ;
  assign n505 = x39 & n504 ;
  assign n506 = x39 | n504 ;
  assign n4740 = ~n423 ;
  assign n507 = n4740 & n424 ;
  assign n508 = n88 & n507 ;
  assign n509 = n429 & n508 ;
  assign n510 = n429 | n508 ;
  assign n4741 = ~n509 ;
  assign n511 = n4741 & n510 ;
  assign n4742 = ~n511 ;
  assign n512 = n506 & n4742 ;
  assign n513 = n505 | n512 ;
  assign n514 = x40 & n513 ;
  assign n515 = x40 | n513 ;
  assign n4743 = ~n432 ;
  assign n516 = n4743 & n433 ;
  assign n517 = n88 & n516 ;
  assign n518 = n438 & n517 ;
  assign n519 = n438 | n517 ;
  assign n4744 = ~n518 ;
  assign n520 = n4744 & n519 ;
  assign n4745 = ~n520 ;
  assign n521 = n515 & n4745 ;
  assign n522 = n514 | n521 ;
  assign n523 = x41 | n522 ;
  assign n524 = x41 & n522 ;
  assign n525 = n132 | n524 ;
  assign n4746 = ~n525 ;
  assign n527 = n523 & n4746 ;
  assign n4747 = ~n527 ;
  assign n528 = n446 & n4747 ;
  assign n4748 = ~x21 ;
  assign n4856 = n4748 & n4602 ;
  assign n4749 = ~n446 ;
  assign n526 = n4749 & n523 ;
  assign n529 = n525 | n526 ;
  assign n87 = ~n529 ;
  assign n530 = x32 & n87 ;
  assign n531 = x22 & n530 ;
  assign n533 = x22 | n530 ;
  assign n4751 = ~n531 ;
  assign n534 = n4751 & n533 ;
  assign n4817 = n4748 & x32 ;
  assign n535 = x33 | n4817 ;
  assign n4752 = ~n534 ;
  assign n536 = n4752 & n535 ;
  assign n537 = n4856 | n536 ;
  assign n538 = x34 & n537 ;
  assign n532 = n4718 & n530 ;
  assign n4753 = ~n530 ;
  assign n539 = x22 & n4753 ;
  assign n540 = n532 | n539 ;
  assign n4754 = ~n540 ;
  assign n541 = n535 & n4754 ;
  assign n542 = n4856 | n541 ;
  assign n543 = x34 | n542 ;
  assign n4755 = ~n4783 ;
  assign n544 = n4755 & n453 ;
  assign n545 = n87 & n544 ;
  assign n546 = n452 & n545 ;
  assign n547 = n452 | n545 ;
  assign n4756 = ~n546 ;
  assign n548 = n4756 & n547 ;
  assign n4757 = ~n548 ;
  assign n549 = n543 & n4757 ;
  assign n550 = n538 | n549 ;
  assign n551 = x35 & n550 ;
  assign n552 = x35 | n550 ;
  assign n553 = x34 | n455 ;
  assign n554 = n456 | n529 ;
  assign n4758 = ~n554 ;
  assign n555 = n553 & n4758 ;
  assign n4759 = ~n555 ;
  assign n556 = n466 & n4759 ;
  assign n557 = n467 & n4758 ;
  assign n558 = n556 | n557 ;
  assign n4760 = ~n558 ;
  assign n559 = n552 & n4760 ;
  assign n560 = n551 | n559 ;
  assign n561 = x36 & n560 ;
  assign n562 = x36 | n560 ;
  assign n4761 = ~n469 ;
  assign n563 = n4761 & n470 ;
  assign n564 = n87 & n563 ;
  assign n565 = n475 & n564 ;
  assign n566 = n475 | n564 ;
  assign n4762 = ~n565 ;
  assign n567 = n4762 & n566 ;
  assign n4763 = ~n567 ;
  assign n568 = n562 & n4763 ;
  assign n569 = n561 | n568 ;
  assign n570 = x37 & n569 ;
  assign n571 = x37 | n569 ;
  assign n4764 = ~n478 ;
  assign n572 = n4764 & n479 ;
  assign n573 = n87 & n572 ;
  assign n574 = n4733 & n573 ;
  assign n4765 = ~n573 ;
  assign n575 = n484 & n4765 ;
  assign n576 = n574 | n575 ;
  assign n4766 = ~n576 ;
  assign n577 = n571 & n4766 ;
  assign n578 = n570 | n577 ;
  assign n579 = x38 & n578 ;
  assign n580 = x38 | n578 ;
  assign n4767 = ~n487 ;
  assign n581 = n4767 & n488 ;
  assign n582 = n87 & n581 ;
  assign n583 = n493 & n582 ;
  assign n584 = n493 | n582 ;
  assign n4768 = ~n583 ;
  assign n585 = n4768 & n584 ;
  assign n4769 = ~n585 ;
  assign n586 = n580 & n4769 ;
  assign n587 = n579 | n586 ;
  assign n588 = x39 & n587 ;
  assign n589 = x39 | n587 ;
  assign n4770 = ~n496 ;
  assign n590 = n4770 & n497 ;
  assign n591 = n87 & n590 ;
  assign n592 = n502 & n591 ;
  assign n593 = n502 | n591 ;
  assign n4771 = ~n592 ;
  assign n594 = n4771 & n593 ;
  assign n4772 = ~n594 ;
  assign n595 = n589 & n4772 ;
  assign n596 = n588 | n595 ;
  assign n597 = x40 & n596 ;
  assign n598 = x40 | n596 ;
  assign n4773 = ~n505 ;
  assign n599 = n4773 & n506 ;
  assign n600 = n87 & n599 ;
  assign n601 = n511 & n600 ;
  assign n602 = n511 | n600 ;
  assign n4774 = ~n601 ;
  assign n603 = n4774 & n602 ;
  assign n4775 = ~n603 ;
  assign n604 = n598 & n4775 ;
  assign n605 = n597 | n604 ;
  assign n606 = x41 & n605 ;
  assign n607 = x41 | n605 ;
  assign n4776 = ~n514 ;
  assign n608 = n4776 & n515 ;
  assign n609 = n87 & n608 ;
  assign n610 = n4745 & n609 ;
  assign n4777 = ~n609 ;
  assign n611 = n520 & n4777 ;
  assign n612 = n610 | n611 ;
  assign n4778 = ~n612 ;
  assign n613 = n607 & n4778 ;
  assign n614 = n606 | n613 ;
  assign n615 = x42 | n614 ;
  assign n616 = x42 & n614 ;
  assign n617 = n131 | n616 ;
  assign n4779 = ~n617 ;
  assign n619 = n615 & n4779 ;
  assign n4780 = ~n619 ;
  assign n620 = n528 & n4780 ;
  assign n4781 = ~x20 ;
  assign n4899 = n4781 & n4602 ;
  assign n4782 = ~n528 ;
  assign n618 = n4782 & n615 ;
  assign n621 = n617 | n618 ;
  assign n86 = ~n621 ;
  assign n622 = x32 & n86 ;
  assign n623 = n4748 & n622 ;
  assign n4784 = ~n622 ;
  assign n624 = x21 & n4784 ;
  assign n625 = n623 | n624 ;
  assign n626 = n4781 & x32 ;
  assign n627 = x33 | n626 ;
  assign n4785 = ~n625 ;
  assign n628 = n4785 & n627 ;
  assign n629 = n4899 | n628 ;
  assign n630 = x34 & n629 ;
  assign n4786 = ~n4856 ;
  assign n631 = n4786 & n535 ;
  assign n632 = n86 & n631 ;
  assign n633 = n534 & n632 ;
  assign n634 = n534 | n632 ;
  assign n4787 = ~n633 ;
  assign n635 = n4787 & n634 ;
  assign n636 = x34 | n629 ;
  assign n4788 = ~n635 ;
  assign n637 = n4788 & n636 ;
  assign n638 = n630 | n637 ;
  assign n639 = x35 & n638 ;
  assign n640 = x35 | n638 ;
  assign n641 = x34 | n537 ;
  assign n642 = n538 | n621 ;
  assign n4789 = ~n642 ;
  assign n643 = n641 & n4789 ;
  assign n4790 = ~n643 ;
  assign n644 = n548 & n4790 ;
  assign n645 = n549 & n4789 ;
  assign n646 = n644 | n645 ;
  assign n4791 = ~n646 ;
  assign n647 = n640 & n4791 ;
  assign n648 = n639 | n647 ;
  assign n649 = x36 & n648 ;
  assign n650 = x36 | n648 ;
  assign n4792 = ~n551 ;
  assign n651 = n4792 & n552 ;
  assign n652 = n86 & n651 ;
  assign n653 = n4760 & n652 ;
  assign n4793 = ~n652 ;
  assign n654 = n558 & n4793 ;
  assign n655 = n653 | n654 ;
  assign n4794 = ~n655 ;
  assign n656 = n650 & n4794 ;
  assign n657 = n649 | n656 ;
  assign n658 = x37 & n657 ;
  assign n659 = x37 | n657 ;
  assign n4795 = ~n561 ;
  assign n660 = n4795 & n562 ;
  assign n661 = n86 & n660 ;
  assign n662 = n4763 & n661 ;
  assign n4796 = ~n661 ;
  assign n663 = n567 & n4796 ;
  assign n664 = n662 | n663 ;
  assign n4797 = ~n664 ;
  assign n665 = n659 & n4797 ;
  assign n666 = n658 | n665 ;
  assign n667 = x38 & n666 ;
  assign n668 = x38 | n666 ;
  assign n4798 = ~n570 ;
  assign n669 = n4798 & n571 ;
  assign n670 = n86 & n669 ;
  assign n671 = n576 & n670 ;
  assign n672 = n576 | n670 ;
  assign n4799 = ~n671 ;
  assign n673 = n4799 & n672 ;
  assign n4800 = ~n673 ;
  assign n674 = n668 & n4800 ;
  assign n675 = n667 | n674 ;
  assign n676 = x39 & n675 ;
  assign n677 = x39 | n675 ;
  assign n4801 = ~n579 ;
  assign n678 = n4801 & n580 ;
  assign n679 = n86 & n678 ;
  assign n680 = n585 & n679 ;
  assign n681 = n585 | n679 ;
  assign n4802 = ~n680 ;
  assign n682 = n4802 & n681 ;
  assign n4803 = ~n682 ;
  assign n683 = n677 & n4803 ;
  assign n684 = n676 | n683 ;
  assign n685 = x40 & n684 ;
  assign n686 = x40 | n684 ;
  assign n4804 = ~n588 ;
  assign n687 = n4804 & n589 ;
  assign n688 = n86 & n687 ;
  assign n689 = n594 & n688 ;
  assign n690 = n594 | n688 ;
  assign n4805 = ~n689 ;
  assign n691 = n4805 & n690 ;
  assign n4806 = ~n691 ;
  assign n692 = n686 & n4806 ;
  assign n693 = n685 | n692 ;
  assign n694 = x41 & n693 ;
  assign n695 = x41 | n693 ;
  assign n4807 = ~n597 ;
  assign n696 = n4807 & n598 ;
  assign n697 = n86 & n696 ;
  assign n698 = n603 & n697 ;
  assign n699 = n603 | n697 ;
  assign n4808 = ~n698 ;
  assign n700 = n4808 & n699 ;
  assign n4809 = ~n700 ;
  assign n701 = n695 & n4809 ;
  assign n702 = n694 | n701 ;
  assign n703 = x42 & n702 ;
  assign n704 = x42 | n702 ;
  assign n4810 = ~n606 ;
  assign n705 = n4810 & n607 ;
  assign n706 = n86 & n705 ;
  assign n707 = n4778 & n706 ;
  assign n4811 = ~n706 ;
  assign n708 = n612 & n4811 ;
  assign n709 = n707 | n708 ;
  assign n4812 = ~n709 ;
  assign n710 = n704 & n4812 ;
  assign n711 = n703 | n710 ;
  assign n712 = x43 | n711 ;
  assign n713 = x43 & n711 ;
  assign n714 = n130 | n713 ;
  assign n4813 = ~n714 ;
  assign n716 = n712 & n4813 ;
  assign n4814 = ~n716 ;
  assign n717 = n620 & n4814 ;
  assign n4815 = ~x19 ;
  assign n4990 = n4815 & n4602 ;
  assign n4816 = ~n620 ;
  assign n715 = n4816 & n712 ;
  assign n718 = n714 | n715 ;
  assign n85 = ~n718 ;
  assign n719 = x32 & n85 ;
  assign n720 = x20 & n719 ;
  assign n722 = x20 | n719 ;
  assign n4818 = ~n720 ;
  assign n723 = n4818 & n722 ;
  assign n4944 = n4815 & x32 ;
  assign n724 = x33 | n4944 ;
  assign n4819 = ~n723 ;
  assign n725 = n4819 & n724 ;
  assign n726 = n4990 | n725 ;
  assign n727 = x34 & n726 ;
  assign n721 = n4781 & n719 ;
  assign n4820 = ~n719 ;
  assign n728 = x20 & n4820 ;
  assign n729 = n721 | n728 ;
  assign n4821 = ~n729 ;
  assign n730 = n724 & n4821 ;
  assign n731 = n4990 | n730 ;
  assign n732 = x34 | n731 ;
  assign n4822 = ~n4899 ;
  assign n733 = n4822 & n627 ;
  assign n734 = n85 & n733 ;
  assign n735 = n4785 & n734 ;
  assign n4823 = ~n734 ;
  assign n736 = n625 & n4823 ;
  assign n737 = n735 | n736 ;
  assign n4824 = ~n737 ;
  assign n738 = n732 & n4824 ;
  assign n739 = n727 | n738 ;
  assign n740 = x35 & n739 ;
  assign n741 = x35 | n739 ;
  assign n4825 = ~n630 ;
  assign n742 = n4825 & n636 ;
  assign n743 = n85 & n742 ;
  assign n744 = n635 & n743 ;
  assign n745 = n635 | n743 ;
  assign n4826 = ~n744 ;
  assign n746 = n4826 & n745 ;
  assign n4827 = ~n746 ;
  assign n747 = n741 & n4827 ;
  assign n748 = n740 | n747 ;
  assign n749 = x36 & n748 ;
  assign n750 = x36 | n748 ;
  assign n4828 = ~n639 ;
  assign n751 = n4828 & n640 ;
  assign n752 = n85 & n751 ;
  assign n753 = n646 & n752 ;
  assign n754 = n646 | n752 ;
  assign n4829 = ~n753 ;
  assign n755 = n4829 & n754 ;
  assign n4830 = ~n755 ;
  assign n756 = n750 & n4830 ;
  assign n757 = n749 | n756 ;
  assign n758 = x37 & n757 ;
  assign n759 = x37 | n757 ;
  assign n4831 = ~n649 ;
  assign n760 = n4831 & n650 ;
  assign n761 = n85 & n760 ;
  assign n762 = n4794 & n761 ;
  assign n4832 = ~n761 ;
  assign n763 = n655 & n4832 ;
  assign n764 = n762 | n763 ;
  assign n4833 = ~n764 ;
  assign n765 = n759 & n4833 ;
  assign n766 = n758 | n765 ;
  assign n767 = x38 & n766 ;
  assign n768 = x38 | n766 ;
  assign n4834 = ~n658 ;
  assign n769 = n4834 & n659 ;
  assign n770 = n85 & n769 ;
  assign n771 = n664 & n770 ;
  assign n772 = n664 | n770 ;
  assign n4835 = ~n771 ;
  assign n773 = n4835 & n772 ;
  assign n4836 = ~n773 ;
  assign n774 = n768 & n4836 ;
  assign n775 = n767 | n774 ;
  assign n776 = x39 & n775 ;
  assign n777 = x39 | n775 ;
  assign n4837 = ~n667 ;
  assign n778 = n4837 & n668 ;
  assign n779 = n85 & n778 ;
  assign n780 = n673 & n779 ;
  assign n781 = n673 | n779 ;
  assign n4838 = ~n780 ;
  assign n782 = n4838 & n781 ;
  assign n4839 = ~n782 ;
  assign n783 = n777 & n4839 ;
  assign n784 = n776 | n783 ;
  assign n785 = x40 & n784 ;
  assign n786 = x40 | n784 ;
  assign n4840 = ~n676 ;
  assign n787 = n4840 & n677 ;
  assign n788 = n85 & n787 ;
  assign n789 = n4803 & n788 ;
  assign n4841 = ~n788 ;
  assign n790 = n682 & n4841 ;
  assign n791 = n789 | n790 ;
  assign n4842 = ~n791 ;
  assign n792 = n786 & n4842 ;
  assign n793 = n785 | n792 ;
  assign n794 = x41 & n793 ;
  assign n795 = x41 | n793 ;
  assign n4843 = ~n685 ;
  assign n796 = n4843 & n686 ;
  assign n797 = n85 & n796 ;
  assign n798 = n691 & n797 ;
  assign n799 = n691 | n797 ;
  assign n4844 = ~n798 ;
  assign n800 = n4844 & n799 ;
  assign n4845 = ~n800 ;
  assign n801 = n795 & n4845 ;
  assign n802 = n794 | n801 ;
  assign n803 = x42 & n802 ;
  assign n804 = x42 | n802 ;
  assign n4846 = ~n694 ;
  assign n805 = n4846 & n695 ;
  assign n806 = n85 & n805 ;
  assign n807 = n4809 & n806 ;
  assign n4847 = ~n806 ;
  assign n808 = n700 & n4847 ;
  assign n809 = n807 | n808 ;
  assign n4848 = ~n809 ;
  assign n810 = n804 & n4848 ;
  assign n811 = n803 | n810 ;
  assign n812 = x43 & n811 ;
  assign n813 = x43 | n811 ;
  assign n4849 = ~n703 ;
  assign n814 = n4849 & n704 ;
  assign n815 = n85 & n814 ;
  assign n816 = n4812 & n815 ;
  assign n4850 = ~n815 ;
  assign n817 = n709 & n4850 ;
  assign n818 = n816 | n817 ;
  assign n4851 = ~n818 ;
  assign n819 = n813 & n4851 ;
  assign n820 = n812 | n819 ;
  assign n821 = x44 | n820 ;
  assign n822 = x44 & n820 ;
  assign n823 = n129 | n822 ;
  assign n4852 = ~n823 ;
  assign n825 = n821 & n4852 ;
  assign n4853 = ~n825 ;
  assign n826 = n717 & n4853 ;
  assign n4854 = ~x18 ;
  assign n5091 = n4854 & n4602 ;
  assign n4855 = ~n717 ;
  assign n824 = n4855 & n821 ;
  assign n827 = n823 | n824 ;
  assign n84 = ~n827 ;
  assign n828 = x32 & n84 ;
  assign n829 = x19 & n828 ;
  assign n831 = x19 | n828 ;
  assign n4857 = ~n829 ;
  assign n832 = n4857 & n831 ;
  assign n5039 = n4854 & x32 ;
  assign n833 = x33 | n5039 ;
  assign n4858 = ~n832 ;
  assign n834 = n4858 & n833 ;
  assign n835 = n5091 | n834 ;
  assign n836 = x34 & n835 ;
  assign n830 = n4815 & n828 ;
  assign n4859 = ~n828 ;
  assign n837 = x19 & n4859 ;
  assign n838 = n830 | n837 ;
  assign n4860 = ~n838 ;
  assign n839 = n833 & n4860 ;
  assign n840 = n5091 | n839 ;
  assign n841 = x34 | n840 ;
  assign n4861 = ~n4990 ;
  assign n842 = n4861 & n724 ;
  assign n843 = n84 & n842 ;
  assign n844 = n723 & n843 ;
  assign n845 = n723 | n843 ;
  assign n4862 = ~n844 ;
  assign n846 = n4862 & n845 ;
  assign n4863 = ~n846 ;
  assign n847 = n841 & n4863 ;
  assign n848 = n836 | n847 ;
  assign n849 = x35 | n848 ;
  assign n850 = x35 & n848 ;
  assign n851 = n727 | n827 ;
  assign n4864 = ~n851 ;
  assign n852 = n738 & n4864 ;
  assign n853 = x34 | n726 ;
  assign n854 = n4864 & n853 ;
  assign n4865 = ~n854 ;
  assign n855 = n737 & n4865 ;
  assign n856 = n852 | n855 ;
  assign n4866 = ~n850 ;
  assign n857 = n4866 & n856 ;
  assign n4867 = ~n857 ;
  assign n858 = n849 & n4867 ;
  assign n859 = x36 & n858 ;
  assign n860 = x36 | n858 ;
  assign n4868 = ~n740 ;
  assign n861 = n4868 & n741 ;
  assign n862 = n84 & n861 ;
  assign n863 = n746 & n862 ;
  assign n864 = n746 | n862 ;
  assign n4869 = ~n863 ;
  assign n865 = n4869 & n864 ;
  assign n4870 = ~n865 ;
  assign n866 = n860 & n4870 ;
  assign n867 = n859 | n866 ;
  assign n868 = x37 & n867 ;
  assign n869 = x37 | n867 ;
  assign n4871 = ~n749 ;
  assign n870 = n4871 & n750 ;
  assign n871 = n84 & n870 ;
  assign n872 = n755 & n871 ;
  assign n873 = n755 | n871 ;
  assign n4872 = ~n872 ;
  assign n874 = n4872 & n873 ;
  assign n4873 = ~n874 ;
  assign n875 = n869 & n4873 ;
  assign n876 = n868 | n875 ;
  assign n877 = x38 & n876 ;
  assign n878 = x38 | n876 ;
  assign n4874 = ~n758 ;
  assign n879 = n4874 & n759 ;
  assign n880 = n84 & n879 ;
  assign n881 = n4833 & n880 ;
  assign n4875 = ~n880 ;
  assign n882 = n764 & n4875 ;
  assign n883 = n881 | n882 ;
  assign n4876 = ~n883 ;
  assign n884 = n878 & n4876 ;
  assign n885 = n877 | n884 ;
  assign n886 = x39 & n885 ;
  assign n887 = x39 | n885 ;
  assign n4877 = ~n767 ;
  assign n888 = n4877 & n768 ;
  assign n889 = n84 & n888 ;
  assign n890 = n773 & n889 ;
  assign n891 = n773 | n889 ;
  assign n4878 = ~n890 ;
  assign n892 = n4878 & n891 ;
  assign n4879 = ~n892 ;
  assign n893 = n887 & n4879 ;
  assign n894 = n886 | n893 ;
  assign n895 = x40 & n894 ;
  assign n896 = x40 | n894 ;
  assign n4880 = ~n776 ;
  assign n897 = n4880 & n777 ;
  assign n898 = n84 & n897 ;
  assign n899 = n782 & n898 ;
  assign n900 = n782 | n898 ;
  assign n4881 = ~n899 ;
  assign n901 = n4881 & n900 ;
  assign n4882 = ~n901 ;
  assign n902 = n896 & n4882 ;
  assign n903 = n895 | n902 ;
  assign n904 = x41 & n903 ;
  assign n905 = x41 | n903 ;
  assign n4883 = ~n785 ;
  assign n906 = n4883 & n786 ;
  assign n907 = n84 & n906 ;
  assign n908 = n4842 & n907 ;
  assign n4884 = ~n907 ;
  assign n909 = n791 & n4884 ;
  assign n910 = n908 | n909 ;
  assign n4885 = ~n910 ;
  assign n911 = n905 & n4885 ;
  assign n912 = n904 | n911 ;
  assign n913 = x42 & n912 ;
  assign n914 = x42 | n912 ;
  assign n4886 = ~n794 ;
  assign n915 = n4886 & n795 ;
  assign n916 = n84 & n915 ;
  assign n917 = n800 & n916 ;
  assign n918 = n800 | n916 ;
  assign n4887 = ~n917 ;
  assign n919 = n4887 & n918 ;
  assign n4888 = ~n919 ;
  assign n920 = n914 & n4888 ;
  assign n921 = n913 | n920 ;
  assign n922 = x43 & n921 ;
  assign n923 = x43 | n921 ;
  assign n4889 = ~n803 ;
  assign n924 = n4889 & n804 ;
  assign n925 = n84 & n924 ;
  assign n926 = n4848 & n925 ;
  assign n4890 = ~n925 ;
  assign n927 = n809 & n4890 ;
  assign n928 = n926 | n927 ;
  assign n4891 = ~n928 ;
  assign n929 = n923 & n4891 ;
  assign n930 = n922 | n929 ;
  assign n931 = x44 & n930 ;
  assign n932 = x44 | n930 ;
  assign n4892 = ~n812 ;
  assign n933 = n4892 & n813 ;
  assign n934 = n84 & n933 ;
  assign n935 = n4851 & n934 ;
  assign n4893 = ~n934 ;
  assign n936 = n818 & n4893 ;
  assign n937 = n935 | n936 ;
  assign n4894 = ~n937 ;
  assign n938 = n932 & n4894 ;
  assign n939 = n931 | n938 ;
  assign n940 = x45 | n939 ;
  assign n941 = x45 & n939 ;
  assign n942 = n128 | n941 ;
  assign n4895 = ~n942 ;
  assign n944 = n940 & n4895 ;
  assign n4896 = ~n944 ;
  assign n945 = n826 & n4896 ;
  assign n4897 = ~x17 ;
  assign n5206 = n4897 & n4602 ;
  assign n4898 = ~n826 ;
  assign n943 = n4898 & n940 ;
  assign n946 = n942 | n943 ;
  assign n83 = ~n946 ;
  assign n947 = x32 & n83 ;
  assign n948 = x18 & n947 ;
  assign n950 = x18 | n947 ;
  assign n4900 = ~n948 ;
  assign n951 = n4900 & n950 ;
  assign n5148 = n4897 & x32 ;
  assign n952 = x33 | n5148 ;
  assign n4901 = ~n951 ;
  assign n953 = n4901 & n952 ;
  assign n954 = n5206 | n953 ;
  assign n955 = x34 & n954 ;
  assign n949 = n4854 & n947 ;
  assign n4902 = ~n947 ;
  assign n956 = x18 & n4902 ;
  assign n957 = n949 | n956 ;
  assign n4903 = ~n957 ;
  assign n958 = n952 & n4903 ;
  assign n959 = n5206 | n958 ;
  assign n960 = x34 | n959 ;
  assign n4904 = ~n5091 ;
  assign n961 = n4904 & n833 ;
  assign n962 = n83 & n961 ;
  assign n963 = n832 & n962 ;
  assign n964 = n832 | n962 ;
  assign n4905 = ~n963 ;
  assign n965 = n4905 & n964 ;
  assign n4906 = ~n965 ;
  assign n966 = n960 & n4906 ;
  assign n967 = n955 | n966 ;
  assign n968 = x35 & n967 ;
  assign n969 = x35 | n967 ;
  assign n970 = x34 | n835 ;
  assign n971 = n836 | n946 ;
  assign n4907 = ~n971 ;
  assign n972 = n970 & n4907 ;
  assign n4908 = ~n972 ;
  assign n973 = n846 & n4908 ;
  assign n974 = n847 & n4907 ;
  assign n975 = n973 | n974 ;
  assign n4909 = ~n975 ;
  assign n976 = n969 & n4909 ;
  assign n977 = n968 | n976 ;
  assign n978 = x36 & n977 ;
  assign n979 = x36 | n977 ;
  assign n980 = n849 & n4866 ;
  assign n981 = n83 & n980 ;
  assign n4910 = ~n856 ;
  assign n982 = n4910 & n981 ;
  assign n4911 = ~n981 ;
  assign n983 = n856 & n4911 ;
  assign n984 = n982 | n983 ;
  assign n4912 = ~n984 ;
  assign n985 = n979 & n4912 ;
  assign n986 = n978 | n985 ;
  assign n987 = x37 & n986 ;
  assign n988 = x37 | n986 ;
  assign n4913 = ~n859 ;
  assign n989 = n4913 & n860 ;
  assign n990 = n83 & n989 ;
  assign n991 = n865 & n990 ;
  assign n992 = n865 | n990 ;
  assign n4914 = ~n991 ;
  assign n993 = n4914 & n992 ;
  assign n4915 = ~n993 ;
  assign n994 = n988 & n4915 ;
  assign n995 = n987 | n994 ;
  assign n996 = x38 & n995 ;
  assign n997 = x38 | n995 ;
  assign n4916 = ~n868 ;
  assign n998 = n4916 & n869 ;
  assign n999 = n83 & n998 ;
  assign n1000 = n874 & n999 ;
  assign n1001 = n874 | n999 ;
  assign n4917 = ~n1000 ;
  assign n1002 = n4917 & n1001 ;
  assign n4918 = ~n1002 ;
  assign n1003 = n997 & n4918 ;
  assign n1004 = n996 | n1003 ;
  assign n1005 = x39 & n1004 ;
  assign n1006 = x39 | n1004 ;
  assign n4919 = ~n877 ;
  assign n1007 = n4919 & n878 ;
  assign n1008 = n83 & n1007 ;
  assign n1009 = n883 & n1008 ;
  assign n1010 = n883 | n1008 ;
  assign n4920 = ~n1009 ;
  assign n1011 = n4920 & n1010 ;
  assign n4921 = ~n1011 ;
  assign n1012 = n1006 & n4921 ;
  assign n1013 = n1005 | n1012 ;
  assign n1014 = x40 & n1013 ;
  assign n1015 = x40 | n1013 ;
  assign n4922 = ~n886 ;
  assign n1016 = n4922 & n887 ;
  assign n1017 = n83 & n1016 ;
  assign n1018 = n892 & n1017 ;
  assign n1019 = n892 | n1017 ;
  assign n4923 = ~n1018 ;
  assign n1020 = n4923 & n1019 ;
  assign n4924 = ~n1020 ;
  assign n1021 = n1015 & n4924 ;
  assign n1022 = n1014 | n1021 ;
  assign n1023 = x41 & n1022 ;
  assign n1024 = x41 | n1022 ;
  assign n4925 = ~n895 ;
  assign n1025 = n4925 & n896 ;
  assign n1026 = n83 & n1025 ;
  assign n1027 = n901 & n1026 ;
  assign n1028 = n901 | n1026 ;
  assign n4926 = ~n1027 ;
  assign n1029 = n4926 & n1028 ;
  assign n4927 = ~n1029 ;
  assign n1030 = n1024 & n4927 ;
  assign n1031 = n1023 | n1030 ;
  assign n1032 = x42 & n1031 ;
  assign n1033 = x42 | n1031 ;
  assign n4928 = ~n904 ;
  assign n1034 = n4928 & n905 ;
  assign n1035 = n83 & n1034 ;
  assign n1036 = n910 & n1035 ;
  assign n1037 = n910 | n1035 ;
  assign n4929 = ~n1036 ;
  assign n1038 = n4929 & n1037 ;
  assign n4930 = ~n1038 ;
  assign n1039 = n1033 & n4930 ;
  assign n1040 = n1032 | n1039 ;
  assign n1041 = x43 & n1040 ;
  assign n1042 = x43 | n1040 ;
  assign n4931 = ~n913 ;
  assign n1043 = n4931 & n914 ;
  assign n1044 = n83 & n1043 ;
  assign n1045 = n919 & n1044 ;
  assign n1046 = n919 | n1044 ;
  assign n4932 = ~n1045 ;
  assign n1047 = n4932 & n1046 ;
  assign n4933 = ~n1047 ;
  assign n1048 = n1042 & n4933 ;
  assign n1049 = n1041 | n1048 ;
  assign n1050 = x44 & n1049 ;
  assign n1051 = x44 | n1049 ;
  assign n4934 = ~n922 ;
  assign n1052 = n4934 & n923 ;
  assign n1053 = n83 & n1052 ;
  assign n1054 = n4891 & n1053 ;
  assign n4935 = ~n1053 ;
  assign n1055 = n928 & n4935 ;
  assign n1056 = n1054 | n1055 ;
  assign n4936 = ~n1056 ;
  assign n1057 = n1051 & n4936 ;
  assign n1058 = n1050 | n1057 ;
  assign n1059 = x45 & n1058 ;
  assign n1060 = x45 | n1058 ;
  assign n4937 = ~n931 ;
  assign n1061 = n4937 & n932 ;
  assign n1062 = n83 & n1061 ;
  assign n1063 = n4894 & n1062 ;
  assign n4938 = ~n1062 ;
  assign n1064 = n937 & n4938 ;
  assign n1065 = n1063 | n1064 ;
  assign n4939 = ~n1065 ;
  assign n1066 = n1060 & n4939 ;
  assign n1067 = n1059 | n1066 ;
  assign n1068 = x46 | n1067 ;
  assign n1069 = x46 & n1067 ;
  assign n1070 = n127 | n1069 ;
  assign n4940 = ~n1070 ;
  assign n1072 = n1068 & n4940 ;
  assign n4941 = ~n1072 ;
  assign n1073 = n945 & n4941 ;
  assign n4942 = ~x16 ;
  assign n5269 = n4942 & n4602 ;
  assign n4943 = ~n945 ;
  assign n1071 = n4943 & n1068 ;
  assign n1074 = n1070 | n1071 ;
  assign n82 = ~n1074 ;
  assign n1075 = x32 & n82 ;
  assign n1076 = n4897 & n1075 ;
  assign n4945 = ~n1075 ;
  assign n1077 = x17 & n4945 ;
  assign n1078 = n1076 | n1077 ;
  assign n1079 = n4942 & x32 ;
  assign n1080 = x33 | n1079 ;
  assign n4946 = ~n1078 ;
  assign n1081 = n4946 & n1080 ;
  assign n1082 = n5269 | n1081 ;
  assign n1083 = x34 & n1082 ;
  assign n4947 = ~n5206 ;
  assign n1084 = n4947 & n952 ;
  assign n1085 = n82 & n1084 ;
  assign n1086 = n951 & n1085 ;
  assign n1087 = n951 | n1085 ;
  assign n4948 = ~n1086 ;
  assign n1088 = n4948 & n1087 ;
  assign n1089 = x34 | n1082 ;
  assign n4949 = ~n1088 ;
  assign n1090 = n4949 & n1089 ;
  assign n1091 = n1083 | n1090 ;
  assign n1092 = x35 & n1091 ;
  assign n1093 = x35 | n1091 ;
  assign n1094 = x34 | n954 ;
  assign n1095 = n955 | n1074 ;
  assign n4950 = ~n1095 ;
  assign n1096 = n1094 & n4950 ;
  assign n4951 = ~n1096 ;
  assign n1097 = n965 & n4951 ;
  assign n1098 = n966 & n4950 ;
  assign n1099 = n1097 | n1098 ;
  assign n4952 = ~n1099 ;
  assign n1100 = n1093 & n4952 ;
  assign n1101 = n1092 | n1100 ;
  assign n1102 = x36 & n1101 ;
  assign n1103 = x36 | n1101 ;
  assign n4953 = ~n968 ;
  assign n1104 = n4953 & n969 ;
  assign n1105 = n82 & n1104 ;
  assign n1106 = n975 & n1105 ;
  assign n1107 = n975 | n1105 ;
  assign n4954 = ~n1106 ;
  assign n1108 = n4954 & n1107 ;
  assign n4955 = ~n1108 ;
  assign n1109 = n1103 & n4955 ;
  assign n1110 = n1102 | n1109 ;
  assign n1111 = x37 & n1110 ;
  assign n1112 = x37 | n1110 ;
  assign n4956 = ~n978 ;
  assign n1113 = n4956 & n979 ;
  assign n1114 = n82 & n1113 ;
  assign n1115 = n984 & n1114 ;
  assign n1116 = n984 | n1114 ;
  assign n4957 = ~n1115 ;
  assign n1117 = n4957 & n1116 ;
  assign n4958 = ~n1117 ;
  assign n1118 = n1112 & n4958 ;
  assign n1119 = n1111 | n1118 ;
  assign n1120 = x38 & n1119 ;
  assign n1121 = x38 | n1119 ;
  assign n4959 = ~n987 ;
  assign n1122 = n4959 & n988 ;
  assign n1123 = n82 & n1122 ;
  assign n1124 = n993 & n1123 ;
  assign n1125 = n993 | n1123 ;
  assign n4960 = ~n1124 ;
  assign n1126 = n4960 & n1125 ;
  assign n4961 = ~n1126 ;
  assign n1127 = n1121 & n4961 ;
  assign n1128 = n1120 | n1127 ;
  assign n1129 = x39 & n1128 ;
  assign n1130 = x39 | n1128 ;
  assign n4962 = ~n996 ;
  assign n1131 = n4962 & n997 ;
  assign n1132 = n82 & n1131 ;
  assign n1133 = n1002 & n1132 ;
  assign n1134 = n1002 | n1132 ;
  assign n4963 = ~n1133 ;
  assign n1135 = n4963 & n1134 ;
  assign n4964 = ~n1135 ;
  assign n1136 = n1130 & n4964 ;
  assign n1137 = n1129 | n1136 ;
  assign n1138 = x40 & n1137 ;
  assign n1139 = x40 | n1137 ;
  assign n4965 = ~n1005 ;
  assign n1140 = n4965 & n1006 ;
  assign n1141 = n82 & n1140 ;
  assign n1142 = n1011 & n1141 ;
  assign n1143 = n1011 | n1141 ;
  assign n4966 = ~n1142 ;
  assign n1144 = n4966 & n1143 ;
  assign n4967 = ~n1144 ;
  assign n1145 = n1139 & n4967 ;
  assign n1146 = n1138 | n1145 ;
  assign n1147 = x41 & n1146 ;
  assign n1148 = x41 | n1146 ;
  assign n4968 = ~n1014 ;
  assign n1149 = n4968 & n1015 ;
  assign n1150 = n82 & n1149 ;
  assign n1151 = n1020 & n1150 ;
  assign n1152 = n1020 | n1150 ;
  assign n4969 = ~n1151 ;
  assign n1153 = n4969 & n1152 ;
  assign n4970 = ~n1153 ;
  assign n1154 = n1148 & n4970 ;
  assign n1155 = n1147 | n1154 ;
  assign n1156 = x42 & n1155 ;
  assign n1157 = x42 | n1155 ;
  assign n4971 = ~n1023 ;
  assign n1158 = n4971 & n1024 ;
  assign n1159 = n82 & n1158 ;
  assign n1160 = n4927 & n1159 ;
  assign n4972 = ~n1159 ;
  assign n1161 = n1029 & n4972 ;
  assign n1162 = n1160 | n1161 ;
  assign n4973 = ~n1162 ;
  assign n1163 = n1157 & n4973 ;
  assign n1164 = n1156 | n1163 ;
  assign n1165 = x43 & n1164 ;
  assign n1166 = x43 | n1164 ;
  assign n4974 = ~n1032 ;
  assign n1167 = n4974 & n1033 ;
  assign n1168 = n82 & n1167 ;
  assign n1169 = n1038 & n1168 ;
  assign n1170 = n1038 | n1168 ;
  assign n4975 = ~n1169 ;
  assign n1171 = n4975 & n1170 ;
  assign n4976 = ~n1171 ;
  assign n1172 = n1166 & n4976 ;
  assign n1173 = n1165 | n1172 ;
  assign n1174 = x44 & n1173 ;
  assign n1175 = x44 | n1173 ;
  assign n4977 = ~n1041 ;
  assign n1176 = n4977 & n1042 ;
  assign n1177 = n82 & n1176 ;
  assign n1178 = n4933 & n1177 ;
  assign n4978 = ~n1177 ;
  assign n1179 = n1047 & n4978 ;
  assign n1180 = n1178 | n1179 ;
  assign n4979 = ~n1180 ;
  assign n1181 = n1175 & n4979 ;
  assign n1182 = n1174 | n1181 ;
  assign n1183 = x45 & n1182 ;
  assign n1184 = x45 | n1182 ;
  assign n4980 = ~n1050 ;
  assign n1185 = n4980 & n1051 ;
  assign n1186 = n82 & n1185 ;
  assign n1187 = n1056 & n1186 ;
  assign n1188 = n1056 | n1186 ;
  assign n4981 = ~n1187 ;
  assign n1189 = n4981 & n1188 ;
  assign n4982 = ~n1189 ;
  assign n1190 = n1184 & n4982 ;
  assign n1191 = n1183 | n1190 ;
  assign n1192 = x46 & n1191 ;
  assign n1193 = x46 | n1191 ;
  assign n4983 = ~n1059 ;
  assign n1194 = n4983 & n1060 ;
  assign n1195 = n82 & n1194 ;
  assign n1196 = n1065 & n1195 ;
  assign n1197 = n1065 | n1195 ;
  assign n4984 = ~n1196 ;
  assign n1198 = n4984 & n1197 ;
  assign n4985 = ~n1198 ;
  assign n1199 = n1193 & n4985 ;
  assign n1200 = n1192 | n1199 ;
  assign n1201 = x47 | n1200 ;
  assign n1202 = x47 & n1200 ;
  assign n1203 = n126 | n1202 ;
  assign n4986 = ~n1203 ;
  assign n1205 = n1201 & n4986 ;
  assign n4987 = ~n1205 ;
  assign n1206 = n1073 & n4987 ;
  assign n4988 = ~x15 ;
  assign n5336 = n4988 & n4602 ;
  assign n4989 = ~n1073 ;
  assign n1204 = n4989 & n1201 ;
  assign n1207 = n1203 | n1204 ;
  assign n81 = ~n1207 ;
  assign n1208 = x32 & n81 ;
  assign n1209 = n4942 & n1208 ;
  assign n4991 = ~n1208 ;
  assign n1210 = x16 & n4991 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = n4988 & x32 ;
  assign n1213 = x33 | n1212 ;
  assign n4992 = ~n1211 ;
  assign n1214 = n4992 & n1213 ;
  assign n1215 = n5336 | n1214 ;
  assign n1216 = x34 & n1215 ;
  assign n4993 = ~n5269 ;
  assign n1217 = n4993 & n1080 ;
  assign n1218 = n81 & n1217 ;
  assign n1219 = n4946 & n1218 ;
  assign n4994 = ~n1218 ;
  assign n1220 = n1078 & n4994 ;
  assign n1221 = n1219 | n1220 ;
  assign n1222 = x34 | n1215 ;
  assign n4995 = ~n1221 ;
  assign n1223 = n4995 & n1222 ;
  assign n1224 = n1216 | n1223 ;
  assign n1225 = x35 & n1224 ;
  assign n1226 = x35 | n1224 ;
  assign n4996 = ~n1083 ;
  assign n1227 = n4996 & n1089 ;
  assign n1228 = n81 & n1227 ;
  assign n1229 = n1088 & n1228 ;
  assign n1230 = n1088 | n1228 ;
  assign n4997 = ~n1229 ;
  assign n1231 = n4997 & n1230 ;
  assign n4998 = ~n1231 ;
  assign n1232 = n1226 & n4998 ;
  assign n1233 = n1225 | n1232 ;
  assign n1234 = x36 & n1233 ;
  assign n1235 = x36 | n1233 ;
  assign n4999 = ~n1092 ;
  assign n1236 = n4999 & n1093 ;
  assign n1237 = n81 & n1236 ;
  assign n1238 = n1099 & n1237 ;
  assign n1239 = n1099 | n1237 ;
  assign n5000 = ~n1238 ;
  assign n1240 = n5000 & n1239 ;
  assign n5001 = ~n1240 ;
  assign n1241 = n1235 & n5001 ;
  assign n1242 = n1234 | n1241 ;
  assign n1243 = x37 & n1242 ;
  assign n1244 = x37 | n1242 ;
  assign n5002 = ~n1102 ;
  assign n1245 = n5002 & n1103 ;
  assign n1246 = n81 & n1245 ;
  assign n1247 = n1108 & n1246 ;
  assign n1248 = n1108 | n1246 ;
  assign n5003 = ~n1247 ;
  assign n1249 = n5003 & n1248 ;
  assign n5004 = ~n1249 ;
  assign n1250 = n1244 & n5004 ;
  assign n1251 = n1243 | n1250 ;
  assign n1252 = x38 & n1251 ;
  assign n1253 = x38 | n1251 ;
  assign n5005 = ~n1111 ;
  assign n1254 = n5005 & n1112 ;
  assign n1255 = n81 & n1254 ;
  assign n1256 = n1117 & n1255 ;
  assign n1257 = n1117 | n1255 ;
  assign n5006 = ~n1256 ;
  assign n1258 = n5006 & n1257 ;
  assign n5007 = ~n1258 ;
  assign n1259 = n1253 & n5007 ;
  assign n1260 = n1252 | n1259 ;
  assign n1261 = x39 & n1260 ;
  assign n1262 = x39 | n1260 ;
  assign n5008 = ~n1120 ;
  assign n1263 = n5008 & n1121 ;
  assign n1264 = n81 & n1263 ;
  assign n1265 = n1126 & n1264 ;
  assign n1266 = n1126 | n1264 ;
  assign n5009 = ~n1265 ;
  assign n1267 = n5009 & n1266 ;
  assign n5010 = ~n1267 ;
  assign n1268 = n1262 & n5010 ;
  assign n1269 = n1261 | n1268 ;
  assign n1270 = x40 & n1269 ;
  assign n1271 = x40 | n1269 ;
  assign n5011 = ~n1129 ;
  assign n1272 = n5011 & n1130 ;
  assign n1273 = n81 & n1272 ;
  assign n1274 = n4964 & n1273 ;
  assign n5012 = ~n1273 ;
  assign n1275 = n1135 & n5012 ;
  assign n1276 = n1274 | n1275 ;
  assign n5013 = ~n1276 ;
  assign n1277 = n1271 & n5013 ;
  assign n1278 = n1270 | n1277 ;
  assign n1279 = x41 & n1278 ;
  assign n1280 = x41 | n1278 ;
  assign n5014 = ~n1138 ;
  assign n1281 = n5014 & n1139 ;
  assign n1282 = n81 & n1281 ;
  assign n1283 = n1144 & n1282 ;
  assign n1284 = n1144 | n1282 ;
  assign n5015 = ~n1283 ;
  assign n1285 = n5015 & n1284 ;
  assign n5016 = ~n1285 ;
  assign n1286 = n1280 & n5016 ;
  assign n1287 = n1279 | n1286 ;
  assign n1288 = x42 & n1287 ;
  assign n1289 = x42 | n1287 ;
  assign n5017 = ~n1147 ;
  assign n1290 = n5017 & n1148 ;
  assign n1291 = n81 & n1290 ;
  assign n1292 = n4970 & n1291 ;
  assign n5018 = ~n1291 ;
  assign n1293 = n1153 & n5018 ;
  assign n1294 = n1292 | n1293 ;
  assign n5019 = ~n1294 ;
  assign n1295 = n1289 & n5019 ;
  assign n1296 = n1288 | n1295 ;
  assign n1297 = x43 & n1296 ;
  assign n1298 = x43 | n1296 ;
  assign n5020 = ~n1156 ;
  assign n1299 = n5020 & n1157 ;
  assign n1300 = n81 & n1299 ;
  assign n1301 = n4973 & n1300 ;
  assign n5021 = ~n1300 ;
  assign n1302 = n1162 & n5021 ;
  assign n1303 = n1301 | n1302 ;
  assign n5022 = ~n1303 ;
  assign n1304 = n1298 & n5022 ;
  assign n1305 = n1297 | n1304 ;
  assign n1306 = x44 & n1305 ;
  assign n1307 = x44 | n1305 ;
  assign n5023 = ~n1165 ;
  assign n1308 = n5023 & n1166 ;
  assign n1309 = n81 & n1308 ;
  assign n1310 = n1171 & n1309 ;
  assign n1311 = n1171 | n1309 ;
  assign n5024 = ~n1310 ;
  assign n1312 = n5024 & n1311 ;
  assign n5025 = ~n1312 ;
  assign n1313 = n1307 & n5025 ;
  assign n1314 = n1306 | n1313 ;
  assign n1315 = x45 & n1314 ;
  assign n1316 = x45 | n1314 ;
  assign n5026 = ~n1174 ;
  assign n1317 = n5026 & n1175 ;
  assign n1318 = n81 & n1317 ;
  assign n1319 = n4979 & n1318 ;
  assign n5027 = ~n1318 ;
  assign n1320 = n1180 & n5027 ;
  assign n1321 = n1319 | n1320 ;
  assign n5028 = ~n1321 ;
  assign n1322 = n1316 & n5028 ;
  assign n1323 = n1315 | n1322 ;
  assign n1324 = x46 & n1323 ;
  assign n1325 = x46 | n1323 ;
  assign n5029 = ~n1183 ;
  assign n1326 = n5029 & n1184 ;
  assign n1327 = n81 & n1326 ;
  assign n1328 = n1189 & n1327 ;
  assign n1329 = n1189 | n1327 ;
  assign n5030 = ~n1328 ;
  assign n1330 = n5030 & n1329 ;
  assign n5031 = ~n1330 ;
  assign n1331 = n1325 & n5031 ;
  assign n1332 = n1324 | n1331 ;
  assign n1333 = x47 & n1332 ;
  assign n1334 = x47 | n1332 ;
  assign n5032 = ~n1192 ;
  assign n1335 = n5032 & n1193 ;
  assign n1336 = n81 & n1335 ;
  assign n1337 = n1198 & n1336 ;
  assign n1338 = n1198 | n1336 ;
  assign n5033 = ~n1337 ;
  assign n1339 = n5033 & n1338 ;
  assign n5034 = ~n1339 ;
  assign n1340 = n1334 & n5034 ;
  assign n1341 = n1333 | n1340 ;
  assign n1342 = x48 | n1341 ;
  assign n1343 = x48 & n1341 ;
  assign n1344 = n125 | n1343 ;
  assign n5035 = ~n1344 ;
  assign n1346 = n1342 & n5035 ;
  assign n5036 = ~n1346 ;
  assign n1347 = n1206 & n5036 ;
  assign n5037 = ~x14 ;
  assign n5404 = n5037 & n4602 ;
  assign n5038 = ~n1206 ;
  assign n1345 = n5038 & n1342 ;
  assign n1348 = n1344 | n1345 ;
  assign n80 = ~n1348 ;
  assign n1349 = x32 & n80 ;
  assign n1350 = n4988 & n1349 ;
  assign n5040 = ~n1349 ;
  assign n1351 = x15 & n5040 ;
  assign n1352 = n1350 | n1351 ;
  assign n1353 = n5037 & x32 ;
  assign n1354 = x33 | n1353 ;
  assign n5041 = ~n1352 ;
  assign n1355 = n5041 & n1354 ;
  assign n1356 = n5404 | n1355 ;
  assign n1357 = x34 & n1356 ;
  assign n5042 = ~n5336 ;
  assign n1358 = n5042 & n1213 ;
  assign n1359 = n80 & n1358 ;
  assign n1360 = n4992 & n1359 ;
  assign n5043 = ~n1359 ;
  assign n1361 = n1211 & n5043 ;
  assign n1362 = n1360 | n1361 ;
  assign n1363 = x34 | n1356 ;
  assign n5044 = ~n1362 ;
  assign n1364 = n5044 & n1363 ;
  assign n1365 = n1357 | n1364 ;
  assign n1366 = x35 & n1365 ;
  assign n1367 = x35 | n1365 ;
  assign n5045 = ~n1216 ;
  assign n1368 = n5045 & n1222 ;
  assign n1369 = n80 & n1368 ;
  assign n1370 = n1221 & n1369 ;
  assign n1371 = n1221 | n1369 ;
  assign n5046 = ~n1370 ;
  assign n1372 = n5046 & n1371 ;
  assign n5047 = ~n1372 ;
  assign n1373 = n1367 & n5047 ;
  assign n1374 = n1366 | n1373 ;
  assign n1375 = x36 & n1374 ;
  assign n1376 = x36 | n1374 ;
  assign n5048 = ~n1225 ;
  assign n1377 = n5048 & n1226 ;
  assign n1378 = n80 & n1377 ;
  assign n1379 = n1231 & n1378 ;
  assign n1380 = n1231 | n1378 ;
  assign n5049 = ~n1379 ;
  assign n1381 = n5049 & n1380 ;
  assign n5050 = ~n1381 ;
  assign n1382 = n1376 & n5050 ;
  assign n1383 = n1375 | n1382 ;
  assign n1384 = x37 & n1383 ;
  assign n1385 = x37 | n1383 ;
  assign n5051 = ~n1234 ;
  assign n1386 = n5051 & n1235 ;
  assign n1387 = n80 & n1386 ;
  assign n1388 = n1240 & n1387 ;
  assign n1389 = n1240 | n1387 ;
  assign n5052 = ~n1388 ;
  assign n1390 = n5052 & n1389 ;
  assign n5053 = ~n1390 ;
  assign n1391 = n1385 & n5053 ;
  assign n1392 = n1384 | n1391 ;
  assign n1393 = x38 & n1392 ;
  assign n1394 = x38 | n1392 ;
  assign n5054 = ~n1243 ;
  assign n1395 = n5054 & n1244 ;
  assign n1396 = n80 & n1395 ;
  assign n1397 = n1249 & n1396 ;
  assign n1398 = n1249 | n1396 ;
  assign n5055 = ~n1397 ;
  assign n1399 = n5055 & n1398 ;
  assign n5056 = ~n1399 ;
  assign n1400 = n1394 & n5056 ;
  assign n1401 = n1393 | n1400 ;
  assign n1402 = x39 & n1401 ;
  assign n1403 = x39 | n1401 ;
  assign n5057 = ~n1252 ;
  assign n1404 = n5057 & n1253 ;
  assign n1405 = n80 & n1404 ;
  assign n1406 = n1258 & n1405 ;
  assign n1407 = n1258 | n1405 ;
  assign n5058 = ~n1406 ;
  assign n1408 = n5058 & n1407 ;
  assign n5059 = ~n1408 ;
  assign n1409 = n1403 & n5059 ;
  assign n1410 = n1402 | n1409 ;
  assign n1411 = x40 & n1410 ;
  assign n1412 = x40 | n1410 ;
  assign n5060 = ~n1261 ;
  assign n1413 = n5060 & n1262 ;
  assign n1414 = n80 & n1413 ;
  assign n1415 = n1267 & n1414 ;
  assign n1416 = n1267 | n1414 ;
  assign n5061 = ~n1415 ;
  assign n1417 = n5061 & n1416 ;
  assign n5062 = ~n1417 ;
  assign n1418 = n1412 & n5062 ;
  assign n1419 = n1411 | n1418 ;
  assign n1420 = x41 & n1419 ;
  assign n1421 = x41 | n1419 ;
  assign n5063 = ~n1270 ;
  assign n1422 = n5063 & n1271 ;
  assign n1423 = n80 & n1422 ;
  assign n1424 = n5013 & n1423 ;
  assign n5064 = ~n1423 ;
  assign n1425 = n1276 & n5064 ;
  assign n1426 = n1424 | n1425 ;
  assign n5065 = ~n1426 ;
  assign n1427 = n1421 & n5065 ;
  assign n1428 = n1420 | n1427 ;
  assign n1429 = x42 & n1428 ;
  assign n1430 = x42 | n1428 ;
  assign n5066 = ~n1279 ;
  assign n1431 = n5066 & n1280 ;
  assign n1432 = n80 & n1431 ;
  assign n1433 = n1285 & n1432 ;
  assign n1434 = n1285 | n1432 ;
  assign n5067 = ~n1433 ;
  assign n1435 = n5067 & n1434 ;
  assign n5068 = ~n1435 ;
  assign n1436 = n1430 & n5068 ;
  assign n1437 = n1429 | n1436 ;
  assign n1438 = x43 & n1437 ;
  assign n1439 = x43 | n1437 ;
  assign n5069 = ~n1288 ;
  assign n1440 = n5069 & n1289 ;
  assign n1441 = n80 & n1440 ;
  assign n1442 = n5019 & n1441 ;
  assign n5070 = ~n1441 ;
  assign n1443 = n1294 & n5070 ;
  assign n1444 = n1442 | n1443 ;
  assign n5071 = ~n1444 ;
  assign n1445 = n1439 & n5071 ;
  assign n1446 = n1438 | n1445 ;
  assign n1447 = x44 & n1446 ;
  assign n1448 = x44 | n1446 ;
  assign n5072 = ~n1297 ;
  assign n1449 = n5072 & n1298 ;
  assign n1450 = n80 & n1449 ;
  assign n1451 = n1303 & n1450 ;
  assign n1452 = n1303 | n1450 ;
  assign n5073 = ~n1451 ;
  assign n1453 = n5073 & n1452 ;
  assign n5074 = ~n1453 ;
  assign n1454 = n1448 & n5074 ;
  assign n1455 = n1447 | n1454 ;
  assign n1456 = x45 & n1455 ;
  assign n1457 = x45 | n1455 ;
  assign n5075 = ~n1306 ;
  assign n1458 = n5075 & n1307 ;
  assign n1459 = n80 & n1458 ;
  assign n1460 = n1312 & n1459 ;
  assign n1461 = n1312 | n1459 ;
  assign n5076 = ~n1460 ;
  assign n1462 = n5076 & n1461 ;
  assign n5077 = ~n1462 ;
  assign n1463 = n1457 & n5077 ;
  assign n1464 = n1456 | n1463 ;
  assign n1465 = x46 & n1464 ;
  assign n1466 = x46 | n1464 ;
  assign n5078 = ~n1315 ;
  assign n1467 = n5078 & n1316 ;
  assign n1468 = n80 & n1467 ;
  assign n1469 = n5028 & n1468 ;
  assign n5079 = ~n1468 ;
  assign n1470 = n1321 & n5079 ;
  assign n1471 = n1469 | n1470 ;
  assign n5080 = ~n1471 ;
  assign n1472 = n1466 & n5080 ;
  assign n1473 = n1465 | n1472 ;
  assign n1474 = x47 & n1473 ;
  assign n1475 = x47 | n1473 ;
  assign n5081 = ~n1324 ;
  assign n1476 = n5081 & n1325 ;
  assign n1477 = n80 & n1476 ;
  assign n1478 = n1330 & n1477 ;
  assign n1479 = n1330 | n1477 ;
  assign n5082 = ~n1478 ;
  assign n1480 = n5082 & n1479 ;
  assign n5083 = ~n1480 ;
  assign n1481 = n1475 & n5083 ;
  assign n1482 = n1474 | n1481 ;
  assign n1483 = x48 & n1482 ;
  assign n1484 = x48 | n1482 ;
  assign n5084 = ~n1333 ;
  assign n1485 = n5084 & n1334 ;
  assign n1486 = n80 & n1485 ;
  assign n1487 = n1339 & n1486 ;
  assign n1488 = n1339 | n1486 ;
  assign n5085 = ~n1487 ;
  assign n1489 = n5085 & n1488 ;
  assign n5086 = ~n1489 ;
  assign n1490 = n1484 & n5086 ;
  assign n1491 = n1483 | n1490 ;
  assign n1492 = x49 | n1491 ;
  assign n1493 = x49 & n1491 ;
  assign n1494 = n124 | n1493 ;
  assign n5087 = ~n1494 ;
  assign n1496 = n1492 & n5087 ;
  assign n5088 = ~n1496 ;
  assign n1497 = n1347 & n5088 ;
  assign n5089 = ~x13 ;
  assign n5564 = n5089 & n4602 ;
  assign n5090 = ~n1347 ;
  assign n1495 = n5090 & n1492 ;
  assign n1498 = n1494 | n1495 ;
  assign n79 = ~n1498 ;
  assign n1499 = x32 & n79 ;
  assign n1500 = x14 & n1499 ;
  assign n1502 = x14 | n1499 ;
  assign n5092 = ~n1500 ;
  assign n1503 = n5092 & n1502 ;
  assign n5498 = n5089 & x32 ;
  assign n1504 = x33 | n5498 ;
  assign n5093 = ~n1503 ;
  assign n1505 = n5093 & n1504 ;
  assign n1506 = n5564 | n1505 ;
  assign n1507 = x34 & n1506 ;
  assign n1501 = n5037 & n1499 ;
  assign n5094 = ~n1499 ;
  assign n1508 = x14 & n5094 ;
  assign n1509 = n1501 | n1508 ;
  assign n5095 = ~n1509 ;
  assign n1510 = n1504 & n5095 ;
  assign n1511 = n5564 | n1510 ;
  assign n1512 = x34 | n1511 ;
  assign n5096 = ~n5404 ;
  assign n1513 = n5096 & n1354 ;
  assign n1514 = n79 & n1513 ;
  assign n1515 = n5041 & n1514 ;
  assign n5097 = ~n1514 ;
  assign n1516 = n1352 & n5097 ;
  assign n1517 = n1515 | n1516 ;
  assign n5098 = ~n1517 ;
  assign n1518 = n1512 & n5098 ;
  assign n1519 = n1507 | n1518 ;
  assign n1520 = x35 & n1519 ;
  assign n5099 = ~n1357 ;
  assign n1521 = n5099 & n1363 ;
  assign n1522 = n79 & n1521 ;
  assign n1523 = n1362 & n1522 ;
  assign n1524 = n1362 | n1522 ;
  assign n5100 = ~n1523 ;
  assign n1525 = n5100 & n1524 ;
  assign n1526 = x35 | n1519 ;
  assign n5101 = ~n1525 ;
  assign n1527 = n5101 & n1526 ;
  assign n1528 = n1520 | n1527 ;
  assign n1529 = x36 & n1528 ;
  assign n1530 = x36 | n1528 ;
  assign n5102 = ~n1366 ;
  assign n1531 = n5102 & n1367 ;
  assign n1532 = n79 & n1531 ;
  assign n1533 = n1372 & n1532 ;
  assign n1534 = n1372 | n1532 ;
  assign n5103 = ~n1533 ;
  assign n1535 = n5103 & n1534 ;
  assign n5104 = ~n1535 ;
  assign n1536 = n1530 & n5104 ;
  assign n1537 = n1529 | n1536 ;
  assign n1538 = x37 & n1537 ;
  assign n1539 = x37 | n1537 ;
  assign n5105 = ~n1375 ;
  assign n1540 = n5105 & n1376 ;
  assign n1541 = n79 & n1540 ;
  assign n1542 = n5050 & n1541 ;
  assign n5106 = ~n1541 ;
  assign n1543 = n1381 & n5106 ;
  assign n1544 = n1542 | n1543 ;
  assign n5107 = ~n1544 ;
  assign n1545 = n1539 & n5107 ;
  assign n1546 = n1538 | n1545 ;
  assign n1547 = x38 & n1546 ;
  assign n1548 = x38 | n1546 ;
  assign n5108 = ~n1384 ;
  assign n1549 = n5108 & n1385 ;
  assign n1550 = n79 & n1549 ;
  assign n1551 = n1390 & n1550 ;
  assign n1552 = n1390 | n1550 ;
  assign n5109 = ~n1551 ;
  assign n1553 = n5109 & n1552 ;
  assign n5110 = ~n1553 ;
  assign n1554 = n1548 & n5110 ;
  assign n1555 = n1547 | n1554 ;
  assign n1556 = x39 & n1555 ;
  assign n1557 = x39 | n1555 ;
  assign n5111 = ~n1393 ;
  assign n1558 = n5111 & n1394 ;
  assign n1559 = n79 & n1558 ;
  assign n1560 = n1399 & n1559 ;
  assign n1561 = n1399 | n1559 ;
  assign n5112 = ~n1560 ;
  assign n1562 = n5112 & n1561 ;
  assign n5113 = ~n1562 ;
  assign n1563 = n1557 & n5113 ;
  assign n1564 = n1556 | n1563 ;
  assign n1565 = x40 & n1564 ;
  assign n1566 = x40 | n1564 ;
  assign n5114 = ~n1402 ;
  assign n1567 = n5114 & n1403 ;
  assign n1568 = n79 & n1567 ;
  assign n1569 = n1408 & n1568 ;
  assign n1570 = n1408 | n1568 ;
  assign n5115 = ~n1569 ;
  assign n1571 = n5115 & n1570 ;
  assign n5116 = ~n1571 ;
  assign n1572 = n1566 & n5116 ;
  assign n1573 = n1565 | n1572 ;
  assign n1574 = x41 & n1573 ;
  assign n1575 = x41 | n1573 ;
  assign n5117 = ~n1411 ;
  assign n1576 = n5117 & n1412 ;
  assign n1577 = n79 & n1576 ;
  assign n1578 = n1417 & n1577 ;
  assign n1579 = n1417 | n1577 ;
  assign n5118 = ~n1578 ;
  assign n1580 = n5118 & n1579 ;
  assign n5119 = ~n1580 ;
  assign n1581 = n1575 & n5119 ;
  assign n1582 = n1574 | n1581 ;
  assign n1583 = x42 & n1582 ;
  assign n1584 = x42 | n1582 ;
  assign n5120 = ~n1420 ;
  assign n1585 = n5120 & n1421 ;
  assign n1586 = n79 & n1585 ;
  assign n1587 = n5065 & n1586 ;
  assign n5121 = ~n1586 ;
  assign n1588 = n1426 & n5121 ;
  assign n1589 = n1587 | n1588 ;
  assign n5122 = ~n1589 ;
  assign n1590 = n1584 & n5122 ;
  assign n1591 = n1583 | n1590 ;
  assign n1592 = x43 & n1591 ;
  assign n1593 = x43 | n1591 ;
  assign n5123 = ~n1429 ;
  assign n1594 = n5123 & n1430 ;
  assign n1595 = n79 & n1594 ;
  assign n1596 = n5068 & n1595 ;
  assign n5124 = ~n1595 ;
  assign n1597 = n1435 & n5124 ;
  assign n1598 = n1596 | n1597 ;
  assign n5125 = ~n1598 ;
  assign n1599 = n1593 & n5125 ;
  assign n1600 = n1592 | n1599 ;
  assign n1601 = x44 & n1600 ;
  assign n1602 = x44 | n1600 ;
  assign n5126 = ~n1438 ;
  assign n1603 = n5126 & n1439 ;
  assign n1604 = n79 & n1603 ;
  assign n1605 = n1444 & n1604 ;
  assign n1606 = n1444 | n1604 ;
  assign n5127 = ~n1605 ;
  assign n1607 = n5127 & n1606 ;
  assign n5128 = ~n1607 ;
  assign n1608 = n1602 & n5128 ;
  assign n1609 = n1601 | n1608 ;
  assign n1610 = x45 & n1609 ;
  assign n1611 = x45 | n1609 ;
  assign n5129 = ~n1447 ;
  assign n1612 = n5129 & n1448 ;
  assign n1613 = n79 & n1612 ;
  assign n1614 = n1453 & n1613 ;
  assign n1615 = n1453 | n1613 ;
  assign n5130 = ~n1614 ;
  assign n1616 = n5130 & n1615 ;
  assign n5131 = ~n1616 ;
  assign n1617 = n1611 & n5131 ;
  assign n1618 = n1610 | n1617 ;
  assign n1619 = x46 & n1618 ;
  assign n1620 = x46 | n1618 ;
  assign n5132 = ~n1456 ;
  assign n1621 = n5132 & n1457 ;
  assign n1622 = n79 & n1621 ;
  assign n1623 = n5077 & n1622 ;
  assign n5133 = ~n1622 ;
  assign n1624 = n1462 & n5133 ;
  assign n1625 = n1623 | n1624 ;
  assign n5134 = ~n1625 ;
  assign n1626 = n1620 & n5134 ;
  assign n1627 = n1619 | n1626 ;
  assign n1628 = x47 & n1627 ;
  assign n1629 = x47 | n1627 ;
  assign n5135 = ~n1465 ;
  assign n1630 = n5135 & n1466 ;
  assign n1631 = n79 & n1630 ;
  assign n1632 = n5080 & n1631 ;
  assign n5136 = ~n1631 ;
  assign n1633 = n1471 & n5136 ;
  assign n1634 = n1632 | n1633 ;
  assign n5137 = ~n1634 ;
  assign n1635 = n1629 & n5137 ;
  assign n1636 = n1628 | n1635 ;
  assign n1637 = x48 & n1636 ;
  assign n1638 = x48 | n1636 ;
  assign n5138 = ~n1474 ;
  assign n1639 = n5138 & n1475 ;
  assign n1640 = n79 & n1639 ;
  assign n1641 = n1480 & n1640 ;
  assign n1642 = n1480 | n1640 ;
  assign n5139 = ~n1641 ;
  assign n1643 = n5139 & n1642 ;
  assign n5140 = ~n1643 ;
  assign n1644 = n1638 & n5140 ;
  assign n1645 = n1637 | n1644 ;
  assign n1646 = x49 & n1645 ;
  assign n1647 = x49 | n1645 ;
  assign n5141 = ~n1483 ;
  assign n1648 = n5141 & n1484 ;
  assign n1649 = n79 & n1648 ;
  assign n1650 = n5086 & n1649 ;
  assign n5142 = ~n1649 ;
  assign n1651 = n1489 & n5142 ;
  assign n1652 = n1650 | n1651 ;
  assign n5143 = ~n1652 ;
  assign n1653 = n1647 & n5143 ;
  assign n1654 = n1646 | n1653 ;
  assign n1655 = x50 | n1654 ;
  assign n1656 = x50 & n1654 ;
  assign n1657 = n123 | n1656 ;
  assign n5144 = ~n1657 ;
  assign n1659 = n1655 & n5144 ;
  assign n5145 = ~n1659 ;
  assign n1660 = n1497 & n5145 ;
  assign n5146 = ~x12 ;
  assign n5641 = n5146 & n4602 ;
  assign n5147 = ~n1497 ;
  assign n1658 = n5147 & n1655 ;
  assign n1661 = n1657 | n1658 ;
  assign n78 = ~n1661 ;
  assign n1662 = x32 & n78 ;
  assign n1663 = n5089 & n1662 ;
  assign n5149 = ~n1662 ;
  assign n1664 = x13 & n5149 ;
  assign n1665 = n1663 | n1664 ;
  assign n1666 = n5146 & x32 ;
  assign n1667 = x33 | n1666 ;
  assign n5150 = ~n1665 ;
  assign n1668 = n5150 & n1667 ;
  assign n1669 = n5641 | n1668 ;
  assign n1670 = x34 & n1669 ;
  assign n5151 = ~n5564 ;
  assign n1671 = n5151 & n1504 ;
  assign n1672 = n78 & n1671 ;
  assign n1673 = n1503 & n1672 ;
  assign n1674 = n1503 | n1672 ;
  assign n5152 = ~n1673 ;
  assign n1675 = n5152 & n1674 ;
  assign n1676 = x34 | n1669 ;
  assign n5153 = ~n1675 ;
  assign n1677 = n5153 & n1676 ;
  assign n1678 = n1670 | n1677 ;
  assign n1679 = x35 & n1678 ;
  assign n1680 = x34 | n1506 ;
  assign n1681 = n1507 | n1661 ;
  assign n5154 = ~n1681 ;
  assign n1682 = n1680 & n5154 ;
  assign n5155 = ~n1682 ;
  assign n1683 = n1517 & n5155 ;
  assign n1684 = n1518 & n5154 ;
  assign n1685 = n1683 | n1684 ;
  assign n1686 = x35 | n1678 ;
  assign n5156 = ~n1685 ;
  assign n1687 = n5156 & n1686 ;
  assign n1688 = n1679 | n1687 ;
  assign n1689 = x36 & n1688 ;
  assign n5157 = ~n1520 ;
  assign n1690 = n5157 & n1526 ;
  assign n1691 = n78 & n1690 ;
  assign n1692 = n1525 & n1691 ;
  assign n1693 = n1525 | n1691 ;
  assign n5158 = ~n1692 ;
  assign n1694 = n5158 & n1693 ;
  assign n1695 = x36 | n1688 ;
  assign n5159 = ~n1694 ;
  assign n1696 = n5159 & n1695 ;
  assign n1697 = n1689 | n1696 ;
  assign n1698 = x37 & n1697 ;
  assign n1699 = x37 | n1697 ;
  assign n5160 = ~n1529 ;
  assign n1700 = n5160 & n1530 ;
  assign n1701 = n78 & n1700 ;
  assign n1702 = n5104 & n1701 ;
  assign n5161 = ~n1701 ;
  assign n1703 = n1535 & n5161 ;
  assign n1704 = n1702 | n1703 ;
  assign n5162 = ~n1704 ;
  assign n1705 = n1699 & n5162 ;
  assign n1706 = n1698 | n1705 ;
  assign n1707 = x38 & n1706 ;
  assign n1708 = x38 | n1706 ;
  assign n5163 = ~n1538 ;
  assign n1709 = n5163 & n1539 ;
  assign n1710 = n78 & n1709 ;
  assign n1711 = n1544 & n1710 ;
  assign n1712 = n1544 | n1710 ;
  assign n5164 = ~n1711 ;
  assign n1713 = n5164 & n1712 ;
  assign n5165 = ~n1713 ;
  assign n1714 = n1708 & n5165 ;
  assign n1715 = n1707 | n1714 ;
  assign n1716 = x39 & n1715 ;
  assign n1717 = x39 | n1715 ;
  assign n5166 = ~n1547 ;
  assign n1718 = n5166 & n1548 ;
  assign n1719 = n78 & n1718 ;
  assign n1720 = n1553 & n1719 ;
  assign n1721 = n1553 | n1719 ;
  assign n5167 = ~n1720 ;
  assign n1722 = n5167 & n1721 ;
  assign n5168 = ~n1722 ;
  assign n1723 = n1717 & n5168 ;
  assign n1724 = n1716 | n1723 ;
  assign n1725 = x40 & n1724 ;
  assign n1726 = x40 | n1724 ;
  assign n5169 = ~n1556 ;
  assign n1727 = n5169 & n1557 ;
  assign n1728 = n78 & n1727 ;
  assign n1729 = n5113 & n1728 ;
  assign n5170 = ~n1728 ;
  assign n1730 = n1562 & n5170 ;
  assign n1731 = n1729 | n1730 ;
  assign n5171 = ~n1731 ;
  assign n1732 = n1726 & n5171 ;
  assign n1733 = n1725 | n1732 ;
  assign n1734 = x41 & n1733 ;
  assign n1735 = x41 | n1733 ;
  assign n5172 = ~n1565 ;
  assign n1736 = n5172 & n1566 ;
  assign n1737 = n78 & n1736 ;
  assign n1738 = n5116 & n1737 ;
  assign n5173 = ~n1737 ;
  assign n1739 = n1571 & n5173 ;
  assign n1740 = n1738 | n1739 ;
  assign n5174 = ~n1740 ;
  assign n1741 = n1735 & n5174 ;
  assign n1742 = n1734 | n1741 ;
  assign n1743 = x42 & n1742 ;
  assign n1744 = x42 | n1742 ;
  assign n5175 = ~n1574 ;
  assign n1745 = n5175 & n1575 ;
  assign n1746 = n78 & n1745 ;
  assign n1747 = n1580 & n1746 ;
  assign n1748 = n1580 | n1746 ;
  assign n5176 = ~n1747 ;
  assign n1749 = n5176 & n1748 ;
  assign n5177 = ~n1749 ;
  assign n1750 = n1744 & n5177 ;
  assign n1751 = n1743 | n1750 ;
  assign n1752 = x43 & n1751 ;
  assign n1753 = x43 | n1751 ;
  assign n5178 = ~n1583 ;
  assign n1754 = n5178 & n1584 ;
  assign n1755 = n78 & n1754 ;
  assign n1756 = n1589 & n1755 ;
  assign n1757 = n1589 | n1755 ;
  assign n5179 = ~n1756 ;
  assign n1758 = n5179 & n1757 ;
  assign n5180 = ~n1758 ;
  assign n1759 = n1753 & n5180 ;
  assign n1760 = n1752 | n1759 ;
  assign n1761 = x44 & n1760 ;
  assign n1762 = x44 | n1760 ;
  assign n5181 = ~n1592 ;
  assign n1763 = n5181 & n1593 ;
  assign n1764 = n78 & n1763 ;
  assign n1765 = n5125 & n1764 ;
  assign n5182 = ~n1764 ;
  assign n1766 = n1598 & n5182 ;
  assign n1767 = n1765 | n1766 ;
  assign n5183 = ~n1767 ;
  assign n1768 = n1762 & n5183 ;
  assign n1769 = n1761 | n1768 ;
  assign n1770 = x45 & n1769 ;
  assign n1771 = x45 | n1769 ;
  assign n5184 = ~n1601 ;
  assign n1772 = n5184 & n1602 ;
  assign n1773 = n78 & n1772 ;
  assign n1774 = n1607 & n1773 ;
  assign n1775 = n1607 | n1773 ;
  assign n5185 = ~n1774 ;
  assign n1776 = n5185 & n1775 ;
  assign n5186 = ~n1776 ;
  assign n1777 = n1771 & n5186 ;
  assign n1778 = n1770 | n1777 ;
  assign n1779 = x46 & n1778 ;
  assign n1780 = x46 | n1778 ;
  assign n5187 = ~n1610 ;
  assign n1781 = n5187 & n1611 ;
  assign n1782 = n78 & n1781 ;
  assign n1783 = n1616 & n1782 ;
  assign n1784 = n1616 | n1782 ;
  assign n5188 = ~n1783 ;
  assign n1785 = n5188 & n1784 ;
  assign n5189 = ~n1785 ;
  assign n1786 = n1780 & n5189 ;
  assign n1787 = n1779 | n1786 ;
  assign n1788 = x47 & n1787 ;
  assign n1789 = x47 | n1787 ;
  assign n5190 = ~n1619 ;
  assign n1790 = n5190 & n1620 ;
  assign n1791 = n78 & n1790 ;
  assign n1792 = n5134 & n1791 ;
  assign n5191 = ~n1791 ;
  assign n1793 = n1625 & n5191 ;
  assign n1794 = n1792 | n1793 ;
  assign n5192 = ~n1794 ;
  assign n1795 = n1789 & n5192 ;
  assign n1796 = n1788 | n1795 ;
  assign n1797 = x48 & n1796 ;
  assign n1798 = x48 | n1796 ;
  assign n5193 = ~n1628 ;
  assign n1799 = n5193 & n1629 ;
  assign n1800 = n78 & n1799 ;
  assign n1801 = n1634 & n1800 ;
  assign n1802 = n1634 | n1800 ;
  assign n5194 = ~n1801 ;
  assign n1803 = n5194 & n1802 ;
  assign n5195 = ~n1803 ;
  assign n1804 = n1798 & n5195 ;
  assign n1805 = n1797 | n1804 ;
  assign n1806 = x49 & n1805 ;
  assign n1807 = x49 | n1805 ;
  assign n5196 = ~n1637 ;
  assign n1808 = n5196 & n1638 ;
  assign n1809 = n78 & n1808 ;
  assign n1810 = n5140 & n1809 ;
  assign n5197 = ~n1809 ;
  assign n1811 = n1643 & n5197 ;
  assign n1812 = n1810 | n1811 ;
  assign n5198 = ~n1812 ;
  assign n1813 = n1807 & n5198 ;
  assign n1814 = n1806 | n1813 ;
  assign n1815 = x50 & n1814 ;
  assign n1816 = x50 | n1814 ;
  assign n5199 = ~n1646 ;
  assign n1817 = n5199 & n1647 ;
  assign n1818 = n78 & n1817 ;
  assign n1819 = n5143 & n1818 ;
  assign n5200 = ~n1818 ;
  assign n1820 = n1652 & n5200 ;
  assign n1821 = n1819 | n1820 ;
  assign n5201 = ~n1821 ;
  assign n1822 = n1816 & n5201 ;
  assign n1823 = n1815 | n1822 ;
  assign n1824 = x51 | n1823 ;
  assign n1825 = x51 & n1823 ;
  assign n1826 = n122 | n1825 ;
  assign n5202 = ~n1826 ;
  assign n1828 = n1824 & n5202 ;
  assign n5203 = ~n1828 ;
  assign n1829 = n1660 & n5203 ;
  assign n5204 = ~x11 ;
  assign n5807 = n5204 & n4602 ;
  assign n5205 = ~n1660 ;
  assign n1827 = n5205 & n1824 ;
  assign n1830 = n1826 | n1827 ;
  assign n77 = ~n1830 ;
  assign n1831 = x32 & n77 ;
  assign n1832 = x12 & n1831 ;
  assign n1834 = x12 | n1831 ;
  assign n5207 = ~n1832 ;
  assign n1835 = n5207 & n1834 ;
  assign n5723 = n5204 & x32 ;
  assign n1836 = x33 | n5723 ;
  assign n5208 = ~n1835 ;
  assign n1837 = n5208 & n1836 ;
  assign n1838 = n5807 | n1837 ;
  assign n1839 = x34 & n1838 ;
  assign n1833 = n5146 & n1831 ;
  assign n5209 = ~n1831 ;
  assign n1840 = x12 & n5209 ;
  assign n1841 = n1833 | n1840 ;
  assign n5210 = ~n1841 ;
  assign n1842 = n1836 & n5210 ;
  assign n1843 = n5807 | n1842 ;
  assign n1844 = x34 | n1843 ;
  assign n5211 = ~n5641 ;
  assign n1845 = n5211 & n1667 ;
  assign n1846 = n77 & n1845 ;
  assign n1847 = n5150 & n1846 ;
  assign n5212 = ~n1846 ;
  assign n1848 = n1665 & n5212 ;
  assign n1849 = n1847 | n1848 ;
  assign n5213 = ~n1849 ;
  assign n1850 = n1844 & n5213 ;
  assign n1851 = n1839 | n1850 ;
  assign n1852 = x35 & n1851 ;
  assign n1853 = x35 | n1851 ;
  assign n5214 = ~n1670 ;
  assign n1854 = n5214 & n1676 ;
  assign n1855 = n77 & n1854 ;
  assign n1856 = n1675 & n1855 ;
  assign n1857 = n1675 | n1855 ;
  assign n5215 = ~n1856 ;
  assign n1858 = n5215 & n1857 ;
  assign n5216 = ~n1858 ;
  assign n1859 = n1853 & n5216 ;
  assign n1860 = n1852 | n1859 ;
  assign n1861 = x36 & n1860 ;
  assign n5217 = ~n1679 ;
  assign n1862 = n5217 & n1686 ;
  assign n1863 = n77 & n1862 ;
  assign n1864 = n1685 & n1863 ;
  assign n1865 = n1685 | n1863 ;
  assign n5218 = ~n1864 ;
  assign n1866 = n5218 & n1865 ;
  assign n1867 = x36 | n1860 ;
  assign n5219 = ~n1866 ;
  assign n1868 = n5219 & n1867 ;
  assign n1869 = n1861 | n1868 ;
  assign n1870 = x37 & n1869 ;
  assign n1871 = x37 | n1869 ;
  assign n5220 = ~n1689 ;
  assign n1872 = n5220 & n1695 ;
  assign n1873 = n77 & n1872 ;
  assign n1874 = n5159 & n1873 ;
  assign n5221 = ~n1873 ;
  assign n1875 = n1694 & n5221 ;
  assign n1876 = n1874 | n1875 ;
  assign n5222 = ~n1876 ;
  assign n1877 = n1871 & n5222 ;
  assign n1878 = n1870 | n1877 ;
  assign n1879 = x38 & n1878 ;
  assign n1880 = x38 | n1878 ;
  assign n5223 = ~n1698 ;
  assign n1881 = n5223 & n1699 ;
  assign n1882 = n77 & n1881 ;
  assign n1883 = n1704 & n1882 ;
  assign n1884 = n1704 | n1882 ;
  assign n5224 = ~n1883 ;
  assign n1885 = n5224 & n1884 ;
  assign n5225 = ~n1885 ;
  assign n1886 = n1880 & n5225 ;
  assign n1887 = n1879 | n1886 ;
  assign n1888 = x39 & n1887 ;
  assign n1889 = x39 | n1887 ;
  assign n5226 = ~n1707 ;
  assign n1890 = n5226 & n1708 ;
  assign n1891 = n77 & n1890 ;
  assign n1892 = n1713 & n1891 ;
  assign n1893 = n1713 | n1891 ;
  assign n5227 = ~n1892 ;
  assign n1894 = n5227 & n1893 ;
  assign n5228 = ~n1894 ;
  assign n1895 = n1889 & n5228 ;
  assign n1896 = n1888 | n1895 ;
  assign n1897 = x40 & n1896 ;
  assign n1898 = x40 | n1896 ;
  assign n5229 = ~n1716 ;
  assign n1899 = n5229 & n1717 ;
  assign n1900 = n77 & n1899 ;
  assign n1901 = n5168 & n1900 ;
  assign n5230 = ~n1900 ;
  assign n1902 = n1722 & n5230 ;
  assign n1903 = n1901 | n1902 ;
  assign n5231 = ~n1903 ;
  assign n1904 = n1898 & n5231 ;
  assign n1905 = n1897 | n1904 ;
  assign n1906 = x41 & n1905 ;
  assign n1907 = x41 | n1905 ;
  assign n5232 = ~n1725 ;
  assign n1908 = n5232 & n1726 ;
  assign n1909 = n77 & n1908 ;
  assign n1910 = n5171 & n1909 ;
  assign n5233 = ~n1909 ;
  assign n1911 = n1731 & n5233 ;
  assign n1912 = n1910 | n1911 ;
  assign n5234 = ~n1912 ;
  assign n1913 = n1907 & n5234 ;
  assign n1914 = n1906 | n1913 ;
  assign n1915 = x42 & n1914 ;
  assign n1916 = x42 | n1914 ;
  assign n5235 = ~n1734 ;
  assign n1917 = n5235 & n1735 ;
  assign n1918 = n77 & n1917 ;
  assign n1919 = n5174 & n1918 ;
  assign n5236 = ~n1918 ;
  assign n1920 = n1740 & n5236 ;
  assign n1921 = n1919 | n1920 ;
  assign n5237 = ~n1921 ;
  assign n1922 = n1916 & n5237 ;
  assign n1923 = n1915 | n1922 ;
  assign n1924 = x43 & n1923 ;
  assign n1925 = x43 | n1923 ;
  assign n5238 = ~n1743 ;
  assign n1926 = n5238 & n1744 ;
  assign n1927 = n77 & n1926 ;
  assign n1928 = n1749 & n1927 ;
  assign n1929 = n1749 | n1927 ;
  assign n5239 = ~n1928 ;
  assign n1930 = n5239 & n1929 ;
  assign n5240 = ~n1930 ;
  assign n1931 = n1925 & n5240 ;
  assign n1932 = n1924 | n1931 ;
  assign n1933 = x44 & n1932 ;
  assign n1934 = x44 | n1932 ;
  assign n5241 = ~n1752 ;
  assign n1935 = n5241 & n1753 ;
  assign n1936 = n77 & n1935 ;
  assign n1937 = n1758 & n1936 ;
  assign n1938 = n1758 | n1936 ;
  assign n5242 = ~n1937 ;
  assign n1939 = n5242 & n1938 ;
  assign n5243 = ~n1939 ;
  assign n1940 = n1934 & n5243 ;
  assign n1941 = n1933 | n1940 ;
  assign n1942 = x45 & n1941 ;
  assign n1943 = x45 | n1941 ;
  assign n5244 = ~n1761 ;
  assign n1944 = n5244 & n1762 ;
  assign n1945 = n77 & n1944 ;
  assign n1946 = n1767 & n1945 ;
  assign n1947 = n1767 | n1945 ;
  assign n5245 = ~n1946 ;
  assign n1948 = n5245 & n1947 ;
  assign n5246 = ~n1948 ;
  assign n1949 = n1943 & n5246 ;
  assign n1950 = n1942 | n1949 ;
  assign n1951 = x46 & n1950 ;
  assign n1952 = x46 | n1950 ;
  assign n5247 = ~n1770 ;
  assign n1953 = n5247 & n1771 ;
  assign n1954 = n77 & n1953 ;
  assign n1955 = n1776 & n1954 ;
  assign n1956 = n1776 | n1954 ;
  assign n5248 = ~n1955 ;
  assign n1957 = n5248 & n1956 ;
  assign n5249 = ~n1957 ;
  assign n1958 = n1952 & n5249 ;
  assign n1959 = n1951 | n1958 ;
  assign n1960 = x47 & n1959 ;
  assign n1961 = x47 | n1959 ;
  assign n5250 = ~n1779 ;
  assign n1962 = n5250 & n1780 ;
  assign n1963 = n77 & n1962 ;
  assign n1964 = n1785 & n1963 ;
  assign n1965 = n1785 | n1963 ;
  assign n5251 = ~n1964 ;
  assign n1966 = n5251 & n1965 ;
  assign n5252 = ~n1966 ;
  assign n1967 = n1961 & n5252 ;
  assign n1968 = n1960 | n1967 ;
  assign n1969 = x48 & n1968 ;
  assign n1970 = x48 | n1968 ;
  assign n5253 = ~n1788 ;
  assign n1971 = n5253 & n1789 ;
  assign n1972 = n77 & n1971 ;
  assign n1973 = n1794 & n1972 ;
  assign n1974 = n1794 | n1972 ;
  assign n5254 = ~n1973 ;
  assign n1975 = n5254 & n1974 ;
  assign n5255 = ~n1975 ;
  assign n1976 = n1970 & n5255 ;
  assign n1977 = n1969 | n1976 ;
  assign n1978 = x49 & n1977 ;
  assign n1979 = x49 | n1977 ;
  assign n5256 = ~n1797 ;
  assign n1980 = n5256 & n1798 ;
  assign n1981 = n77 & n1980 ;
  assign n1982 = n1803 & n1981 ;
  assign n1983 = n1803 | n1981 ;
  assign n5257 = ~n1982 ;
  assign n1984 = n5257 & n1983 ;
  assign n5258 = ~n1984 ;
  assign n1985 = n1979 & n5258 ;
  assign n1986 = n1978 | n1985 ;
  assign n1987 = x50 & n1986 ;
  assign n1988 = x50 | n1986 ;
  assign n5259 = ~n1806 ;
  assign n1989 = n5259 & n1807 ;
  assign n1990 = n77 & n1989 ;
  assign n1991 = n5198 & n1990 ;
  assign n5260 = ~n1990 ;
  assign n1992 = n1812 & n5260 ;
  assign n1993 = n1991 | n1992 ;
  assign n5261 = ~n1993 ;
  assign n1994 = n1988 & n5261 ;
  assign n1995 = n1987 | n1994 ;
  assign n1996 = x51 & n1995 ;
  assign n1997 = x51 | n1995 ;
  assign n5262 = ~n1815 ;
  assign n1998 = n5262 & n1816 ;
  assign n1999 = n77 & n1998 ;
  assign n2000 = n5201 & n1999 ;
  assign n5263 = ~n1999 ;
  assign n2001 = n1821 & n5263 ;
  assign n2002 = n2000 | n2001 ;
  assign n5264 = ~n2002 ;
  assign n2003 = n1997 & n5264 ;
  assign n2004 = n1996 | n2003 ;
  assign n2005 = x52 | n2004 ;
  assign n2006 = x52 & n2004 ;
  assign n2007 = n121 | n2006 ;
  assign n5265 = ~n2007 ;
  assign n2009 = n2005 & n5265 ;
  assign n5266 = ~n2009 ;
  assign n2010 = n1829 & n5266 ;
  assign n5267 = ~x10 ;
  assign n5986 = n5267 & n4602 ;
  assign n5268 = ~n1829 ;
  assign n2008 = n5268 & n2005 ;
  assign n2011 = n2007 | n2008 ;
  assign n76 = ~n2011 ;
  assign n2012 = x32 & n76 ;
  assign n2013 = x11 & n2012 ;
  assign n2015 = x11 | n2012 ;
  assign n5270 = ~n2013 ;
  assign n2016 = n5270 & n2015 ;
  assign n5896 = n5267 & x32 ;
  assign n2017 = x33 | n5896 ;
  assign n5271 = ~n2016 ;
  assign n2018 = n5271 & n2017 ;
  assign n2019 = n5986 | n2018 ;
  assign n2020 = x34 & n2019 ;
  assign n2014 = n5204 & n2012 ;
  assign n5272 = ~n2012 ;
  assign n2021 = x11 & n5272 ;
  assign n2022 = n2014 | n2021 ;
  assign n5273 = ~n2022 ;
  assign n2023 = n2017 & n5273 ;
  assign n2024 = n5986 | n2023 ;
  assign n2025 = x34 | n2024 ;
  assign n5274 = ~n5807 ;
  assign n2026 = n5274 & n1836 ;
  assign n2027 = n76 & n2026 ;
  assign n2028 = n1835 & n2027 ;
  assign n2029 = n1835 | n2027 ;
  assign n5275 = ~n2028 ;
  assign n2030 = n5275 & n2029 ;
  assign n5276 = ~n2030 ;
  assign n2031 = n2025 & n5276 ;
  assign n2032 = n2020 | n2031 ;
  assign n2033 = x35 | n2032 ;
  assign n2034 = x35 & n2032 ;
  assign n2035 = n1839 | n2011 ;
  assign n5277 = ~n2035 ;
  assign n2036 = n1850 & n5277 ;
  assign n2037 = x34 | n1838 ;
  assign n2038 = n5277 & n2037 ;
  assign n5278 = ~n2038 ;
  assign n2039 = n1849 & n5278 ;
  assign n2040 = n2036 | n2039 ;
  assign n5279 = ~n2034 ;
  assign n2041 = n5279 & n2040 ;
  assign n5280 = ~n2041 ;
  assign n2042 = n2033 & n5280 ;
  assign n2043 = x36 & n2042 ;
  assign n2044 = x36 | n2042 ;
  assign n5281 = ~n1852 ;
  assign n2045 = n5281 & n1853 ;
  assign n2046 = n76 & n2045 ;
  assign n2047 = n1858 & n2046 ;
  assign n2048 = n1858 | n2046 ;
  assign n5282 = ~n2047 ;
  assign n2049 = n5282 & n2048 ;
  assign n5283 = ~n2049 ;
  assign n2050 = n2044 & n5283 ;
  assign n2051 = n2043 | n2050 ;
  assign n2052 = x37 & n2051 ;
  assign n5284 = ~n1861 ;
  assign n2053 = n5284 & n1867 ;
  assign n2054 = n76 & n2053 ;
  assign n2055 = n1866 & n2054 ;
  assign n2056 = n1866 | n2054 ;
  assign n5285 = ~n2055 ;
  assign n2057 = n5285 & n2056 ;
  assign n2058 = x37 | n2051 ;
  assign n5286 = ~n2057 ;
  assign n2059 = n5286 & n2058 ;
  assign n2060 = n2052 | n2059 ;
  assign n2061 = x38 & n2060 ;
  assign n5287 = ~n1870 ;
  assign n2062 = n5287 & n1871 ;
  assign n2063 = n76 & n2062 ;
  assign n2064 = n1876 & n2063 ;
  assign n2065 = n1876 | n2063 ;
  assign n5288 = ~n2064 ;
  assign n2066 = n5288 & n2065 ;
  assign n2067 = x38 | n2060 ;
  assign n5289 = ~n2066 ;
  assign n2068 = n5289 & n2067 ;
  assign n2069 = n2061 | n2068 ;
  assign n2070 = x39 & n2069 ;
  assign n2071 = x39 | n2069 ;
  assign n5290 = ~n1879 ;
  assign n2072 = n5290 & n1880 ;
  assign n2073 = n76 & n2072 ;
  assign n2074 = n1885 & n2073 ;
  assign n2075 = n1885 | n2073 ;
  assign n5291 = ~n2074 ;
  assign n2076 = n5291 & n2075 ;
  assign n5292 = ~n2076 ;
  assign n2077 = n2071 & n5292 ;
  assign n2078 = n2070 | n2077 ;
  assign n2079 = x40 & n2078 ;
  assign n2080 = x40 | n2078 ;
  assign n5293 = ~n1888 ;
  assign n2081 = n5293 & n1889 ;
  assign n2082 = n76 & n2081 ;
  assign n2083 = n1894 & n2082 ;
  assign n2084 = n1894 | n2082 ;
  assign n5294 = ~n2083 ;
  assign n2085 = n5294 & n2084 ;
  assign n5295 = ~n2085 ;
  assign n2086 = n2080 & n5295 ;
  assign n2087 = n2079 | n2086 ;
  assign n2088 = x41 & n2087 ;
  assign n2089 = x41 | n2087 ;
  assign n5296 = ~n1897 ;
  assign n2090 = n5296 & n1898 ;
  assign n2091 = n76 & n2090 ;
  assign n2092 = n5231 & n2091 ;
  assign n5297 = ~n2091 ;
  assign n2093 = n1903 & n5297 ;
  assign n2094 = n2092 | n2093 ;
  assign n5298 = ~n2094 ;
  assign n2095 = n2089 & n5298 ;
  assign n2096 = n2088 | n2095 ;
  assign n2097 = x42 & n2096 ;
  assign n2098 = x42 | n2096 ;
  assign n5299 = ~n1906 ;
  assign n2099 = n5299 & n1907 ;
  assign n2100 = n76 & n2099 ;
  assign n2101 = n5234 & n2100 ;
  assign n5300 = ~n2100 ;
  assign n2102 = n1912 & n5300 ;
  assign n2103 = n2101 | n2102 ;
  assign n5301 = ~n2103 ;
  assign n2104 = n2098 & n5301 ;
  assign n2105 = n2097 | n2104 ;
  assign n2106 = x43 & n2105 ;
  assign n2107 = x43 | n2105 ;
  assign n5302 = ~n1915 ;
  assign n2108 = n5302 & n1916 ;
  assign n2109 = n76 & n2108 ;
  assign n2110 = n1921 & n2109 ;
  assign n2111 = n1921 | n2109 ;
  assign n5303 = ~n2110 ;
  assign n2112 = n5303 & n2111 ;
  assign n5304 = ~n2112 ;
  assign n2113 = n2107 & n5304 ;
  assign n2114 = n2106 | n2113 ;
  assign n2115 = x44 & n2114 ;
  assign n2116 = x44 | n2114 ;
  assign n5305 = ~n1924 ;
  assign n2117 = n5305 & n1925 ;
  assign n2118 = n76 & n2117 ;
  assign n2119 = n1930 & n2118 ;
  assign n2120 = n1930 | n2118 ;
  assign n5306 = ~n2119 ;
  assign n2121 = n5306 & n2120 ;
  assign n5307 = ~n2121 ;
  assign n2122 = n2116 & n5307 ;
  assign n2123 = n2115 | n2122 ;
  assign n2124 = x45 & n2123 ;
  assign n2125 = x45 | n2123 ;
  assign n5308 = ~n1933 ;
  assign n2126 = n5308 & n1934 ;
  assign n2127 = n76 & n2126 ;
  assign n2128 = n1939 & n2127 ;
  assign n2129 = n1939 | n2127 ;
  assign n5309 = ~n2128 ;
  assign n2130 = n5309 & n2129 ;
  assign n5310 = ~n2130 ;
  assign n2131 = n2125 & n5310 ;
  assign n2132 = n2124 | n2131 ;
  assign n2133 = x46 & n2132 ;
  assign n2134 = x46 | n2132 ;
  assign n5311 = ~n1942 ;
  assign n2135 = n5311 & n1943 ;
  assign n2136 = n76 & n2135 ;
  assign n2137 = n1948 & n2136 ;
  assign n2138 = n1948 | n2136 ;
  assign n5312 = ~n2137 ;
  assign n2139 = n5312 & n2138 ;
  assign n5313 = ~n2139 ;
  assign n2140 = n2134 & n5313 ;
  assign n2141 = n2133 | n2140 ;
  assign n2142 = x47 & n2141 ;
  assign n2143 = x47 | n2141 ;
  assign n5314 = ~n1951 ;
  assign n2144 = n5314 & n1952 ;
  assign n2145 = n76 & n2144 ;
  assign n2146 = n1957 & n2145 ;
  assign n2147 = n1957 | n2145 ;
  assign n5315 = ~n2146 ;
  assign n2148 = n5315 & n2147 ;
  assign n5316 = ~n2148 ;
  assign n2149 = n2143 & n5316 ;
  assign n2150 = n2142 | n2149 ;
  assign n2151 = x48 & n2150 ;
  assign n2152 = x48 | n2150 ;
  assign n5317 = ~n1960 ;
  assign n2153 = n5317 & n1961 ;
  assign n2154 = n76 & n2153 ;
  assign n2155 = n1966 & n2154 ;
  assign n2156 = n1966 | n2154 ;
  assign n5318 = ~n2155 ;
  assign n2157 = n5318 & n2156 ;
  assign n5319 = ~n2157 ;
  assign n2158 = n2152 & n5319 ;
  assign n2159 = n2151 | n2158 ;
  assign n2160 = x49 & n2159 ;
  assign n2161 = x49 | n2159 ;
  assign n5320 = ~n1969 ;
  assign n2162 = n5320 & n1970 ;
  assign n2163 = n76 & n2162 ;
  assign n2164 = n1975 & n2163 ;
  assign n2165 = n1975 | n2163 ;
  assign n5321 = ~n2164 ;
  assign n2166 = n5321 & n2165 ;
  assign n5322 = ~n2166 ;
  assign n2167 = n2161 & n5322 ;
  assign n2168 = n2160 | n2167 ;
  assign n2169 = x50 & n2168 ;
  assign n2170 = x50 | n2168 ;
  assign n5323 = ~n1978 ;
  assign n2171 = n5323 & n1979 ;
  assign n2172 = n76 & n2171 ;
  assign n2173 = n1984 & n2172 ;
  assign n2174 = n1984 | n2172 ;
  assign n5324 = ~n2173 ;
  assign n2175 = n5324 & n2174 ;
  assign n5325 = ~n2175 ;
  assign n2176 = n2170 & n5325 ;
  assign n2177 = n2169 | n2176 ;
  assign n2178 = x51 & n2177 ;
  assign n2179 = x51 | n2177 ;
  assign n5326 = ~n1987 ;
  assign n2180 = n5326 & n1988 ;
  assign n2181 = n76 & n2180 ;
  assign n2182 = n5261 & n2181 ;
  assign n5327 = ~n2181 ;
  assign n2183 = n1993 & n5327 ;
  assign n2184 = n2182 | n2183 ;
  assign n5328 = ~n2184 ;
  assign n2185 = n2179 & n5328 ;
  assign n2186 = n2178 | n2185 ;
  assign n2187 = x52 & n2186 ;
  assign n2188 = x52 | n2186 ;
  assign n5329 = ~n1996 ;
  assign n2189 = n5329 & n1997 ;
  assign n2190 = n76 & n2189 ;
  assign n2191 = n5264 & n2190 ;
  assign n5330 = ~n2190 ;
  assign n2192 = n2002 & n5330 ;
  assign n2193 = n2191 | n2192 ;
  assign n5331 = ~n2193 ;
  assign n2194 = n2188 & n5331 ;
  assign n2195 = n2187 | n2194 ;
  assign n2196 = x53 | n2195 ;
  assign n2197 = x53 & n2195 ;
  assign n2198 = n120 | n2197 ;
  assign n5332 = ~n2198 ;
  assign n2200 = n2196 & n5332 ;
  assign n5333 = ~n2200 ;
  assign n2201 = n2010 & n5333 ;
  assign n5334 = ~x9 ;
  assign n6084 = n5334 & n4602 ;
  assign n5335 = ~n2010 ;
  assign n2199 = n5335 & n2196 ;
  assign n2202 = n2198 | n2199 ;
  assign n75 = ~n2202 ;
  assign n2203 = x32 & n75 ;
  assign n2204 = n5267 & n2203 ;
  assign n5337 = ~n2203 ;
  assign n2205 = x10 & n5337 ;
  assign n2206 = n2204 | n2205 ;
  assign n2207 = n5334 & x32 ;
  assign n2208 = x33 | n2207 ;
  assign n5338 = ~n2206 ;
  assign n2209 = n5338 & n2208 ;
  assign n2210 = n6084 | n2209 ;
  assign n2211 = x34 & n2210 ;
  assign n5339 = ~n5986 ;
  assign n2212 = n5339 & n2017 ;
  assign n2213 = n75 & n2212 ;
  assign n2214 = n2016 & n2213 ;
  assign n2215 = n2016 | n2213 ;
  assign n5340 = ~n2214 ;
  assign n2216 = n5340 & n2215 ;
  assign n2217 = x34 | n2210 ;
  assign n5341 = ~n2216 ;
  assign n2218 = n5341 & n2217 ;
  assign n2219 = n2211 | n2218 ;
  assign n2222 = x35 | n2219 ;
  assign n2220 = x35 & n2219 ;
  assign n2223 = n2020 | n2202 ;
  assign n5342 = ~n2223 ;
  assign n2224 = n2031 & n5342 ;
  assign n2225 = x34 | n2019 ;
  assign n2226 = n5342 & n2225 ;
  assign n5343 = ~n2226 ;
  assign n2227 = n2030 & n5343 ;
  assign n2228 = n2224 | n2227 ;
  assign n5344 = ~n2220 ;
  assign n2229 = n5344 & n2228 ;
  assign n5345 = ~n2229 ;
  assign n2230 = n2222 & n5345 ;
  assign n2231 = x36 & n2230 ;
  assign n2232 = x36 | n2230 ;
  assign n2233 = n2033 & n5279 ;
  assign n2234 = n75 & n2233 ;
  assign n5346 = ~n2040 ;
  assign n2235 = n5346 & n2234 ;
  assign n5347 = ~n2234 ;
  assign n2236 = n2040 & n5347 ;
  assign n2237 = n2235 | n2236 ;
  assign n5348 = ~n2237 ;
  assign n2238 = n2232 & n5348 ;
  assign n2239 = n2231 | n2238 ;
  assign n2240 = x37 & n2239 ;
  assign n2241 = x37 | n2239 ;
  assign n5349 = ~n2043 ;
  assign n2242 = n5349 & n2044 ;
  assign n2243 = n75 & n2242 ;
  assign n2244 = n2049 & n2243 ;
  assign n2245 = n2049 | n2243 ;
  assign n5350 = ~n2244 ;
  assign n2246 = n5350 & n2245 ;
  assign n5351 = ~n2246 ;
  assign n2247 = n2241 & n5351 ;
  assign n2248 = n2240 | n2247 ;
  assign n2249 = x38 & n2248 ;
  assign n5352 = ~n2052 ;
  assign n2250 = n5352 & n2058 ;
  assign n2251 = n75 & n2250 ;
  assign n2252 = n2057 & n2251 ;
  assign n2253 = n2057 | n2251 ;
  assign n5353 = ~n2252 ;
  assign n2254 = n5353 & n2253 ;
  assign n2255 = x38 | n2248 ;
  assign n5354 = ~n2254 ;
  assign n2256 = n5354 & n2255 ;
  assign n2257 = n2249 | n2256 ;
  assign n2258 = x39 & n2257 ;
  assign n5355 = ~n2061 ;
  assign n2259 = n5355 & n2067 ;
  assign n2260 = n75 & n2259 ;
  assign n2261 = n2066 & n2260 ;
  assign n2262 = n2066 | n2260 ;
  assign n5356 = ~n2261 ;
  assign n2263 = n5356 & n2262 ;
  assign n2264 = x39 | n2257 ;
  assign n5357 = ~n2263 ;
  assign n2265 = n5357 & n2264 ;
  assign n2266 = n2258 | n2265 ;
  assign n2267 = x40 & n2266 ;
  assign n2268 = x40 | n2266 ;
  assign n5358 = ~n2070 ;
  assign n2269 = n5358 & n2071 ;
  assign n2270 = n75 & n2269 ;
  assign n2271 = n2076 & n2270 ;
  assign n2272 = n2076 | n2270 ;
  assign n5359 = ~n2271 ;
  assign n2273 = n5359 & n2272 ;
  assign n5360 = ~n2273 ;
  assign n2274 = n2268 & n5360 ;
  assign n2275 = n2267 | n2274 ;
  assign n2276 = x41 & n2275 ;
  assign n2277 = x41 | n2275 ;
  assign n5361 = ~n2079 ;
  assign n2278 = n5361 & n2080 ;
  assign n2279 = n75 & n2278 ;
  assign n2280 = n2085 & n2279 ;
  assign n2281 = n2085 | n2279 ;
  assign n5362 = ~n2280 ;
  assign n2282 = n5362 & n2281 ;
  assign n5363 = ~n2282 ;
  assign n2283 = n2277 & n5363 ;
  assign n2284 = n2276 | n2283 ;
  assign n2285 = x42 & n2284 ;
  assign n2286 = x42 | n2284 ;
  assign n5364 = ~n2088 ;
  assign n2287 = n5364 & n2089 ;
  assign n2288 = n75 & n2287 ;
  assign n2289 = n5298 & n2288 ;
  assign n5365 = ~n2288 ;
  assign n2290 = n2094 & n5365 ;
  assign n2291 = n2289 | n2290 ;
  assign n5366 = ~n2291 ;
  assign n2292 = n2286 & n5366 ;
  assign n2293 = n2285 | n2292 ;
  assign n2294 = x43 & n2293 ;
  assign n2295 = x43 | n2293 ;
  assign n5367 = ~n2097 ;
  assign n2296 = n5367 & n2098 ;
  assign n2297 = n75 & n2296 ;
  assign n2298 = n2103 & n2297 ;
  assign n2299 = n2103 | n2297 ;
  assign n5368 = ~n2298 ;
  assign n2300 = n5368 & n2299 ;
  assign n5369 = ~n2300 ;
  assign n2301 = n2295 & n5369 ;
  assign n2302 = n2294 | n2301 ;
  assign n2303 = x44 & n2302 ;
  assign n2304 = x44 | n2302 ;
  assign n5370 = ~n2106 ;
  assign n2305 = n5370 & n2107 ;
  assign n2306 = n75 & n2305 ;
  assign n2307 = n2112 & n2306 ;
  assign n2308 = n2112 | n2306 ;
  assign n5371 = ~n2307 ;
  assign n2309 = n5371 & n2308 ;
  assign n5372 = ~n2309 ;
  assign n2310 = n2304 & n5372 ;
  assign n2311 = n2303 | n2310 ;
  assign n2312 = x45 & n2311 ;
  assign n2313 = x45 | n2311 ;
  assign n5373 = ~n2115 ;
  assign n2314 = n5373 & n2116 ;
  assign n2315 = n75 & n2314 ;
  assign n2316 = n5307 & n2315 ;
  assign n5374 = ~n2315 ;
  assign n2317 = n2121 & n5374 ;
  assign n2318 = n2316 | n2317 ;
  assign n5375 = ~n2318 ;
  assign n2319 = n2313 & n5375 ;
  assign n2320 = n2312 | n2319 ;
  assign n2321 = x46 & n2320 ;
  assign n2322 = x46 | n2320 ;
  assign n5376 = ~n2124 ;
  assign n2323 = n5376 & n2125 ;
  assign n2324 = n75 & n2323 ;
  assign n2325 = n2130 & n2324 ;
  assign n2326 = n2130 | n2324 ;
  assign n5377 = ~n2325 ;
  assign n2327 = n5377 & n2326 ;
  assign n5378 = ~n2327 ;
  assign n2328 = n2322 & n5378 ;
  assign n2329 = n2321 | n2328 ;
  assign n2330 = x47 & n2329 ;
  assign n2331 = x47 | n2329 ;
  assign n5379 = ~n2133 ;
  assign n2332 = n5379 & n2134 ;
  assign n2333 = n75 & n2332 ;
  assign n2334 = n2139 & n2333 ;
  assign n2335 = n2139 | n2333 ;
  assign n5380 = ~n2334 ;
  assign n2336 = n5380 & n2335 ;
  assign n5381 = ~n2336 ;
  assign n2337 = n2331 & n5381 ;
  assign n2338 = n2330 | n2337 ;
  assign n2339 = x48 & n2338 ;
  assign n2340 = x48 | n2338 ;
  assign n5382 = ~n2142 ;
  assign n2341 = n5382 & n2143 ;
  assign n2342 = n75 & n2341 ;
  assign n2343 = n2148 & n2342 ;
  assign n2344 = n2148 | n2342 ;
  assign n5383 = ~n2343 ;
  assign n2345 = n5383 & n2344 ;
  assign n5384 = ~n2345 ;
  assign n2346 = n2340 & n5384 ;
  assign n2347 = n2339 | n2346 ;
  assign n2348 = x49 & n2347 ;
  assign n2349 = x49 | n2347 ;
  assign n5385 = ~n2151 ;
  assign n2350 = n5385 & n2152 ;
  assign n2351 = n75 & n2350 ;
  assign n2352 = n5319 & n2351 ;
  assign n5386 = ~n2351 ;
  assign n2353 = n2157 & n5386 ;
  assign n2354 = n2352 | n2353 ;
  assign n5387 = ~n2354 ;
  assign n2355 = n2349 & n5387 ;
  assign n2356 = n2348 | n2355 ;
  assign n2357 = x50 & n2356 ;
  assign n2358 = x50 | n2356 ;
  assign n5388 = ~n2160 ;
  assign n2359 = n5388 & n2161 ;
  assign n2360 = n75 & n2359 ;
  assign n2361 = n2166 & n2360 ;
  assign n2362 = n2166 | n2360 ;
  assign n5389 = ~n2361 ;
  assign n2363 = n5389 & n2362 ;
  assign n5390 = ~n2363 ;
  assign n2364 = n2358 & n5390 ;
  assign n2365 = n2357 | n2364 ;
  assign n2366 = x51 & n2365 ;
  assign n2367 = x51 | n2365 ;
  assign n5391 = ~n2169 ;
  assign n2368 = n5391 & n2170 ;
  assign n2369 = n75 & n2368 ;
  assign n2370 = n2175 & n2369 ;
  assign n2371 = n2175 | n2369 ;
  assign n5392 = ~n2370 ;
  assign n2372 = n5392 & n2371 ;
  assign n5393 = ~n2372 ;
  assign n2373 = n2367 & n5393 ;
  assign n2374 = n2366 | n2373 ;
  assign n2375 = x52 & n2374 ;
  assign n2376 = x52 | n2374 ;
  assign n5394 = ~n2178 ;
  assign n2377 = n5394 & n2179 ;
  assign n2378 = n75 & n2377 ;
  assign n2379 = n2184 & n2378 ;
  assign n2380 = n2184 | n2378 ;
  assign n5395 = ~n2379 ;
  assign n2381 = n5395 & n2380 ;
  assign n5396 = ~n2381 ;
  assign n2382 = n2376 & n5396 ;
  assign n2383 = n2375 | n2382 ;
  assign n2384 = x53 & n2383 ;
  assign n2385 = x53 | n2383 ;
  assign n5397 = ~n2187 ;
  assign n2386 = n5397 & n2188 ;
  assign n2387 = n75 & n2386 ;
  assign n2388 = n2193 & n2387 ;
  assign n2389 = n2193 | n2387 ;
  assign n5398 = ~n2388 ;
  assign n2390 = n5398 & n2389 ;
  assign n5399 = ~n2390 ;
  assign n2391 = n2385 & n5399 ;
  assign n2392 = n2384 | n2391 ;
  assign n2393 = x54 | n2392 ;
  assign n2394 = x54 & n2392 ;
  assign n2395 = n119 | n2394 ;
  assign n5400 = ~n2395 ;
  assign n2397 = n2393 & n5400 ;
  assign n5401 = ~n2397 ;
  assign n2398 = n2201 & n5401 ;
  assign n5402 = ~x8 ;
  assign n97 = n5402 & n4602 ;
  assign n5403 = ~n2201 ;
  assign n2396 = n5403 & n2393 ;
  assign n2399 = n2395 | n2396 ;
  assign n74 = ~n2399 ;
  assign n2400 = x32 & n74 ;
  assign n2401 = x9 & n2400 ;
  assign n2403 = x9 | n2400 ;
  assign n5405 = ~n2401 ;
  assign n2404 = n5405 & n2403 ;
  assign n6218 = n5402 & x32 ;
  assign n2405 = x33 | n6218 ;
  assign n5406 = ~n2404 ;
  assign n2406 = n5406 & n2405 ;
  assign n2407 = n97 | n2406 ;
  assign n2408 = x34 & n2407 ;
  assign n2402 = n5334 & n2400 ;
  assign n5407 = ~n2400 ;
  assign n2409 = x9 & n5407 ;
  assign n2410 = n2402 | n2409 ;
  assign n5408 = ~n2410 ;
  assign n2411 = n2405 & n5408 ;
  assign n2412 = n97 | n2411 ;
  assign n2413 = x34 | n2412 ;
  assign n5409 = ~n6084 ;
  assign n2414 = n5409 & n2208 ;
  assign n2415 = n74 & n2414 ;
  assign n2416 = n5338 & n2415 ;
  assign n5410 = ~n2415 ;
  assign n2417 = n2206 & n5410 ;
  assign n2418 = n2416 | n2417 ;
  assign n5411 = ~n2418 ;
  assign n2419 = n2413 & n5411 ;
  assign n2420 = n2408 | n2419 ;
  assign n2421 = x35 | n2420 ;
  assign n2422 = x35 & n2420 ;
  assign n5412 = ~n2211 ;
  assign n2423 = n5412 & n2217 ;
  assign n2424 = n74 & n2423 ;
  assign n5413 = ~n2424 ;
  assign n2425 = n2216 & n5413 ;
  assign n2426 = n5341 & n2424 ;
  assign n2427 = n2425 | n2426 ;
  assign n5414 = ~n2422 ;
  assign n2428 = n5414 & n2427 ;
  assign n5415 = ~n2428 ;
  assign n2429 = n2421 & n5415 ;
  assign n2430 = x36 | n2429 ;
  assign n2431 = x36 & n2429 ;
  assign n5416 = ~x35 ;
  assign n2221 = n5416 & n2219 ;
  assign n5417 = ~n2219 ;
  assign n2432 = x35 & n5417 ;
  assign n2433 = n2221 | n2432 ;
  assign n2434 = n74 & n2433 ;
  assign n5418 = ~n2228 ;
  assign n2435 = n5418 & n2434 ;
  assign n5419 = ~n2434 ;
  assign n2436 = n2228 & n5419 ;
  assign n2437 = n2435 | n2436 ;
  assign n5420 = ~n2431 ;
  assign n2438 = n5420 & n2437 ;
  assign n5421 = ~n2438 ;
  assign n2439 = n2430 & n5421 ;
  assign n2440 = x37 | n2439 ;
  assign n2441 = x37 & n2439 ;
  assign n5422 = ~n2231 ;
  assign n2442 = n5422 & n2232 ;
  assign n2443 = n74 & n2442 ;
  assign n2444 = n2237 & n2443 ;
  assign n2445 = n2237 | n2443 ;
  assign n5423 = ~n2444 ;
  assign n2446 = n5423 & n2445 ;
  assign n5424 = ~n2441 ;
  assign n2447 = n5424 & n2446 ;
  assign n5425 = ~n2447 ;
  assign n2448 = n2440 & n5425 ;
  assign n2449 = x38 | n2448 ;
  assign n2450 = x38 & n2448 ;
  assign n5426 = ~n2240 ;
  assign n2451 = n5426 & n2241 ;
  assign n2452 = n74 & n2451 ;
  assign n2453 = n5351 & n2452 ;
  assign n5427 = ~n2452 ;
  assign n2454 = n2246 & n5427 ;
  assign n2455 = n2453 | n2454 ;
  assign n5428 = ~n2450 ;
  assign n2456 = n5428 & n2455 ;
  assign n5429 = ~n2456 ;
  assign n2457 = n2449 & n5429 ;
  assign n2458 = x39 | n2457 ;
  assign n5430 = ~n2249 ;
  assign n2459 = n5430 & n2255 ;
  assign n2460 = n74 & n2459 ;
  assign n2461 = n2254 & n2460 ;
  assign n2462 = n2254 | n2460 ;
  assign n5431 = ~n2461 ;
  assign n2463 = n5431 & n2462 ;
  assign n2464 = x39 & n2457 ;
  assign n5432 = ~n2464 ;
  assign n2465 = n2463 & n5432 ;
  assign n5433 = ~n2465 ;
  assign n2466 = n2458 & n5433 ;
  assign n2467 = x40 | n2466 ;
  assign n2468 = x40 & n2466 ;
  assign n5434 = ~n2258 ;
  assign n2469 = n5434 & n2264 ;
  assign n2470 = n74 & n2469 ;
  assign n2471 = n2263 & n2470 ;
  assign n2472 = n2263 | n2470 ;
  assign n5435 = ~n2471 ;
  assign n2473 = n5435 & n2472 ;
  assign n5436 = ~n2468 ;
  assign n2474 = n5436 & n2473 ;
  assign n5437 = ~n2474 ;
  assign n2475 = n2467 & n5437 ;
  assign n2476 = x41 | n2475 ;
  assign n2477 = x41 & n2475 ;
  assign n5438 = ~n2267 ;
  assign n2478 = n5438 & n2268 ;
  assign n2479 = n74 & n2478 ;
  assign n2480 = n2273 & n2479 ;
  assign n2481 = n2273 | n2479 ;
  assign n5439 = ~n2480 ;
  assign n2482 = n5439 & n2481 ;
  assign n5440 = ~n2477 ;
  assign n2483 = n5440 & n2482 ;
  assign n5441 = ~n2483 ;
  assign n2484 = n2476 & n5441 ;
  assign n2485 = x42 | n2484 ;
  assign n2486 = x42 & n2484 ;
  assign n5442 = ~n2276 ;
  assign n2487 = n5442 & n2277 ;
  assign n2488 = n74 & n2487 ;
  assign n2489 = n2282 & n2488 ;
  assign n2490 = n2282 | n2488 ;
  assign n5443 = ~n2489 ;
  assign n2491 = n5443 & n2490 ;
  assign n5444 = ~n2486 ;
  assign n2492 = n5444 & n2491 ;
  assign n5445 = ~n2492 ;
  assign n2493 = n2485 & n5445 ;
  assign n2494 = x43 | n2493 ;
  assign n2495 = x43 & n2493 ;
  assign n5446 = ~n2285 ;
  assign n2496 = n5446 & n2286 ;
  assign n2497 = n74 & n2496 ;
  assign n2498 = n2291 & n2497 ;
  assign n2499 = n2291 | n2497 ;
  assign n5447 = ~n2498 ;
  assign n2500 = n5447 & n2499 ;
  assign n5448 = ~n2495 ;
  assign n2501 = n5448 & n2500 ;
  assign n5449 = ~n2501 ;
  assign n2502 = n2494 & n5449 ;
  assign n2503 = x44 | n2502 ;
  assign n2504 = x44 & n2502 ;
  assign n5450 = ~n2294 ;
  assign n2505 = n5450 & n2295 ;
  assign n2506 = n74 & n2505 ;
  assign n2507 = n2300 & n2506 ;
  assign n2508 = n2300 | n2506 ;
  assign n5451 = ~n2507 ;
  assign n2509 = n5451 & n2508 ;
  assign n5452 = ~n2504 ;
  assign n2510 = n5452 & n2509 ;
  assign n5453 = ~n2510 ;
  assign n2511 = n2503 & n5453 ;
  assign n2512 = x45 | n2511 ;
  assign n2513 = x45 & n2511 ;
  assign n5454 = ~n2303 ;
  assign n2514 = n5454 & n2304 ;
  assign n2515 = n74 & n2514 ;
  assign n2516 = n2309 & n2515 ;
  assign n2517 = n2309 | n2515 ;
  assign n5455 = ~n2516 ;
  assign n2518 = n5455 & n2517 ;
  assign n5456 = ~n2513 ;
  assign n2519 = n5456 & n2518 ;
  assign n5457 = ~n2519 ;
  assign n2520 = n2512 & n5457 ;
  assign n2521 = x46 | n2520 ;
  assign n2522 = x46 & n2520 ;
  assign n5458 = ~n2312 ;
  assign n2523 = n5458 & n2313 ;
  assign n2524 = n74 & n2523 ;
  assign n2525 = n5375 & n2524 ;
  assign n5459 = ~n2524 ;
  assign n2526 = n2318 & n5459 ;
  assign n2527 = n2525 | n2526 ;
  assign n5460 = ~n2522 ;
  assign n2528 = n5460 & n2527 ;
  assign n5461 = ~n2528 ;
  assign n2529 = n2521 & n5461 ;
  assign n2530 = x47 | n2529 ;
  assign n2531 = x47 & n2529 ;
  assign n5462 = ~n2321 ;
  assign n2532 = n5462 & n2322 ;
  assign n2533 = n74 & n2532 ;
  assign n2534 = n2327 & n2533 ;
  assign n2535 = n2327 | n2533 ;
  assign n5463 = ~n2534 ;
  assign n2536 = n5463 & n2535 ;
  assign n5464 = ~n2531 ;
  assign n2537 = n5464 & n2536 ;
  assign n5465 = ~n2537 ;
  assign n2538 = n2530 & n5465 ;
  assign n2539 = x48 | n2538 ;
  assign n2540 = x48 & n2538 ;
  assign n5466 = ~n2330 ;
  assign n2541 = n5466 & n2331 ;
  assign n2542 = n74 & n2541 ;
  assign n2543 = n2336 & n2542 ;
  assign n2544 = n2336 | n2542 ;
  assign n5467 = ~n2543 ;
  assign n2545 = n5467 & n2544 ;
  assign n5468 = ~n2540 ;
  assign n2546 = n5468 & n2545 ;
  assign n5469 = ~n2546 ;
  assign n2547 = n2539 & n5469 ;
  assign n2548 = x49 | n2547 ;
  assign n2549 = x49 & n2547 ;
  assign n5470 = ~n2339 ;
  assign n2550 = n5470 & n2340 ;
  assign n2551 = n74 & n2550 ;
  assign n2552 = n2345 & n2551 ;
  assign n2553 = n2345 | n2551 ;
  assign n5471 = ~n2552 ;
  assign n2554 = n5471 & n2553 ;
  assign n5472 = ~n2549 ;
  assign n2555 = n5472 & n2554 ;
  assign n5473 = ~n2555 ;
  assign n2556 = n2548 & n5473 ;
  assign n2557 = x50 | n2556 ;
  assign n2558 = x50 & n2556 ;
  assign n5474 = ~n2348 ;
  assign n2559 = n5474 & n2349 ;
  assign n2560 = n74 & n2559 ;
  assign n2561 = n5387 & n2560 ;
  assign n5475 = ~n2560 ;
  assign n2562 = n2354 & n5475 ;
  assign n2563 = n2561 | n2562 ;
  assign n5476 = ~n2558 ;
  assign n2564 = n5476 & n2563 ;
  assign n5477 = ~n2564 ;
  assign n2565 = n2557 & n5477 ;
  assign n2566 = x51 | n2565 ;
  assign n2567 = x51 & n2565 ;
  assign n5478 = ~n2357 ;
  assign n2568 = n5478 & n2358 ;
  assign n2569 = n74 & n2568 ;
  assign n2570 = n2363 & n2569 ;
  assign n2571 = n2363 | n2569 ;
  assign n5479 = ~n2570 ;
  assign n2572 = n5479 & n2571 ;
  assign n5480 = ~n2567 ;
  assign n2573 = n5480 & n2572 ;
  assign n5481 = ~n2573 ;
  assign n2574 = n2566 & n5481 ;
  assign n2575 = x52 | n2574 ;
  assign n2576 = x52 & n2574 ;
  assign n5482 = ~n2366 ;
  assign n2577 = n5482 & n2367 ;
  assign n2578 = n74 & n2577 ;
  assign n2579 = n5393 & n2578 ;
  assign n5483 = ~n2578 ;
  assign n2580 = n2372 & n5483 ;
  assign n2581 = n2579 | n2580 ;
  assign n5484 = ~n2576 ;
  assign n2582 = n5484 & n2581 ;
  assign n5485 = ~n2582 ;
  assign n2583 = n2575 & n5485 ;
  assign n2584 = x53 | n2583 ;
  assign n2585 = x53 & n2583 ;
  assign n5486 = ~n2375 ;
  assign n2586 = n5486 & n2376 ;
  assign n2587 = n74 & n2586 ;
  assign n2588 = n2381 & n2587 ;
  assign n2589 = n2381 | n2587 ;
  assign n5487 = ~n2588 ;
  assign n2590 = n5487 & n2589 ;
  assign n5488 = ~n2585 ;
  assign n2591 = n5488 & n2590 ;
  assign n5489 = ~n2591 ;
  assign n2592 = n2584 & n5489 ;
  assign n2593 = x54 | n2592 ;
  assign n2594 = x54 & n2592 ;
  assign n5490 = ~n2384 ;
  assign n2595 = n5490 & n2385 ;
  assign n2596 = n74 & n2595 ;
  assign n2597 = n2390 & n2596 ;
  assign n2598 = n2390 | n2596 ;
  assign n5491 = ~n2597 ;
  assign n2599 = n5491 & n2598 ;
  assign n5492 = ~n2594 ;
  assign n2600 = n5492 & n2599 ;
  assign n5493 = ~n2600 ;
  assign n2601 = n2593 & n5493 ;
  assign n2602 = x55 | n2601 ;
  assign n2603 = x55 & n2601 ;
  assign n2604 = n118 | n2603 ;
  assign n5494 = ~n2604 ;
  assign n2605 = n2602 & n5494 ;
  assign n5495 = ~n2605 ;
  assign n2606 = n2398 & n5495 ;
  assign n5496 = ~x7 ;
  assign n99 = n5496 & n4602 ;
  assign n5497 = ~n2398 ;
  assign n2607 = n5497 & n2602 ;
  assign n2608 = n2604 | n2607 ;
  assign n73 = ~n2608 ;
  assign n2609 = x32 & n73 ;
  assign n2610 = x8 & n2609 ;
  assign n2612 = x8 | n2609 ;
  assign n5499 = ~n2610 ;
  assign n2613 = n5499 & n2612 ;
  assign n98 = n5496 & x32 ;
  assign n2614 = x33 | n98 ;
  assign n5500 = ~n2613 ;
  assign n2615 = n5500 & n2614 ;
  assign n2616 = n99 | n2615 ;
  assign n2617 = x34 & n2616 ;
  assign n2611 = n5402 & n2609 ;
  assign n5501 = ~n2609 ;
  assign n2618 = x8 & n5501 ;
  assign n2619 = n2611 | n2618 ;
  assign n5502 = ~n2619 ;
  assign n2620 = n2614 & n5502 ;
  assign n2621 = n99 | n2620 ;
  assign n2622 = x34 | n2621 ;
  assign n5503 = ~n97 ;
  assign n2623 = n5503 & n2405 ;
  assign n2624 = n73 & n2623 ;
  assign n2625 = n2404 & n2624 ;
  assign n2626 = n2404 | n2624 ;
  assign n5504 = ~n2625 ;
  assign n2627 = n5504 & n2626 ;
  assign n5505 = ~n2627 ;
  assign n2628 = n2622 & n5505 ;
  assign n2629 = n2617 | n2628 ;
  assign n2630 = x35 & n2629 ;
  assign n2631 = x35 | n2629 ;
  assign n2632 = x34 | n2407 ;
  assign n2633 = n2408 | n2608 ;
  assign n5506 = ~n2633 ;
  assign n2634 = n2632 & n5506 ;
  assign n5507 = ~n2634 ;
  assign n2635 = n2418 & n5507 ;
  assign n2636 = n2419 & n5506 ;
  assign n2637 = n2635 | n2636 ;
  assign n5508 = ~n2637 ;
  assign n2638 = n2631 & n5508 ;
  assign n2639 = n2630 | n2638 ;
  assign n2640 = x36 & n2639 ;
  assign n2641 = x36 | n2639 ;
  assign n2642 = n2421 & n5414 ;
  assign n2643 = n73 & n2642 ;
  assign n5509 = ~n2427 ;
  assign n2644 = n5509 & n2643 ;
  assign n5510 = ~n2643 ;
  assign n2645 = n2427 & n5510 ;
  assign n2646 = n2644 | n2645 ;
  assign n5511 = ~n2646 ;
  assign n2647 = n2641 & n5511 ;
  assign n2648 = n2640 | n2647 ;
  assign n2649 = x37 & n2648 ;
  assign n2650 = x37 | n2648 ;
  assign n2651 = n2430 & n5420 ;
  assign n2652 = n73 & n2651 ;
  assign n2653 = n2437 & n2652 ;
  assign n2654 = n2437 | n2652 ;
  assign n5512 = ~n2653 ;
  assign n2655 = n5512 & n2654 ;
  assign n5513 = ~n2655 ;
  assign n2656 = n2650 & n5513 ;
  assign n2657 = n2649 | n2656 ;
  assign n2658 = x38 & n2657 ;
  assign n2659 = x38 | n2657 ;
  assign n2660 = n2440 & n5424 ;
  assign n2661 = n73 & n2660 ;
  assign n2662 = n2446 & n2661 ;
  assign n2663 = n2446 | n2661 ;
  assign n5514 = ~n2662 ;
  assign n2664 = n5514 & n2663 ;
  assign n5515 = ~n2664 ;
  assign n2665 = n2659 & n5515 ;
  assign n2666 = n2658 | n2665 ;
  assign n2667 = x39 & n2666 ;
  assign n2668 = x39 | n2666 ;
  assign n2669 = n2449 & n5428 ;
  assign n2670 = n73 & n2669 ;
  assign n5516 = ~n2455 ;
  assign n2671 = n5516 & n2670 ;
  assign n5517 = ~n2670 ;
  assign n2672 = n2455 & n5517 ;
  assign n2673 = n2671 | n2672 ;
  assign n5518 = ~n2673 ;
  assign n2674 = n2668 & n5518 ;
  assign n2675 = n2667 | n2674 ;
  assign n2676 = x40 & n2675 ;
  assign n2677 = n2458 & n5432 ;
  assign n2678 = n73 & n2677 ;
  assign n2679 = n2463 & n2678 ;
  assign n2680 = n2463 | n2678 ;
  assign n5519 = ~n2679 ;
  assign n2681 = n5519 & n2680 ;
  assign n2682 = x40 | n2675 ;
  assign n5520 = ~n2681 ;
  assign n2683 = n5520 & n2682 ;
  assign n2684 = n2676 | n2683 ;
  assign n2685 = x41 & n2684 ;
  assign n2686 = n2467 & n5436 ;
  assign n2687 = n73 & n2686 ;
  assign n5521 = ~n2473 ;
  assign n2688 = n5521 & n2687 ;
  assign n5522 = ~n2687 ;
  assign n2689 = n2473 & n5522 ;
  assign n2690 = n2688 | n2689 ;
  assign n2691 = x41 | n2684 ;
  assign n5523 = ~n2690 ;
  assign n2692 = n5523 & n2691 ;
  assign n2693 = n2685 | n2692 ;
  assign n2694 = x42 & n2693 ;
  assign n2695 = x42 | n2693 ;
  assign n2696 = n2476 & n5440 ;
  assign n2697 = n73 & n2696 ;
  assign n5524 = ~n2482 ;
  assign n2698 = n5524 & n2697 ;
  assign n5525 = ~n2697 ;
  assign n2699 = n2482 & n5525 ;
  assign n2700 = n2698 | n2699 ;
  assign n5526 = ~n2700 ;
  assign n2701 = n2695 & n5526 ;
  assign n2702 = n2694 | n2701 ;
  assign n2703 = x43 & n2702 ;
  assign n2704 = x43 | n2702 ;
  assign n2705 = n2485 & n5444 ;
  assign n2706 = n73 & n2705 ;
  assign n5527 = ~n2491 ;
  assign n2707 = n5527 & n2706 ;
  assign n5528 = ~n2706 ;
  assign n2708 = n2491 & n5528 ;
  assign n2709 = n2707 | n2708 ;
  assign n5529 = ~n2709 ;
  assign n2710 = n2704 & n5529 ;
  assign n2711 = n2703 | n2710 ;
  assign n2712 = x44 & n2711 ;
  assign n2713 = x44 | n2711 ;
  assign n2714 = n2494 & n5448 ;
  assign n2715 = n73 & n2714 ;
  assign n2716 = n2500 & n2715 ;
  assign n2717 = n2500 | n2715 ;
  assign n5530 = ~n2716 ;
  assign n2718 = n5530 & n2717 ;
  assign n5531 = ~n2718 ;
  assign n2719 = n2713 & n5531 ;
  assign n2720 = n2712 | n2719 ;
  assign n2721 = x45 & n2720 ;
  assign n2722 = x45 | n2720 ;
  assign n2723 = n2503 & n5452 ;
  assign n2724 = n73 & n2723 ;
  assign n2725 = n2509 & n2724 ;
  assign n2726 = n2509 | n2724 ;
  assign n5532 = ~n2725 ;
  assign n2727 = n5532 & n2726 ;
  assign n5533 = ~n2727 ;
  assign n2728 = n2722 & n5533 ;
  assign n2729 = n2721 | n2728 ;
  assign n2730 = x46 & n2729 ;
  assign n2731 = x46 | n2729 ;
  assign n2732 = n2512 & n5456 ;
  assign n2733 = n73 & n2732 ;
  assign n5534 = ~n2518 ;
  assign n2734 = n5534 & n2733 ;
  assign n5535 = ~n2733 ;
  assign n2735 = n2518 & n5535 ;
  assign n2736 = n2734 | n2735 ;
  assign n5536 = ~n2736 ;
  assign n2737 = n2731 & n5536 ;
  assign n2738 = n2730 | n2737 ;
  assign n2739 = x47 & n2738 ;
  assign n2740 = x47 | n2738 ;
  assign n2741 = n2521 & n5460 ;
  assign n2742 = n73 & n2741 ;
  assign n5537 = ~n2527 ;
  assign n2743 = n5537 & n2742 ;
  assign n5538 = ~n2742 ;
  assign n2744 = n2527 & n5538 ;
  assign n2745 = n2743 | n2744 ;
  assign n5539 = ~n2745 ;
  assign n2746 = n2740 & n5539 ;
  assign n2747 = n2739 | n2746 ;
  assign n2748 = x48 & n2747 ;
  assign n2749 = x48 | n2747 ;
  assign n2750 = n2530 & n5464 ;
  assign n2751 = n73 & n2750 ;
  assign n2752 = n2536 & n2751 ;
  assign n2753 = n2536 | n2751 ;
  assign n5540 = ~n2752 ;
  assign n2754 = n5540 & n2753 ;
  assign n5541 = ~n2754 ;
  assign n2755 = n2749 & n5541 ;
  assign n2756 = n2748 | n2755 ;
  assign n2757 = x49 & n2756 ;
  assign n2758 = x49 | n2756 ;
  assign n2759 = n2539 & n5468 ;
  assign n2760 = n73 & n2759 ;
  assign n5542 = ~n2545 ;
  assign n2761 = n5542 & n2760 ;
  assign n5543 = ~n2760 ;
  assign n2762 = n2545 & n5543 ;
  assign n2763 = n2761 | n2762 ;
  assign n5544 = ~n2763 ;
  assign n2764 = n2758 & n5544 ;
  assign n2765 = n2757 | n2764 ;
  assign n2766 = x50 & n2765 ;
  assign n2767 = x50 | n2765 ;
  assign n2768 = n2548 & n5472 ;
  assign n2769 = n73 & n2768 ;
  assign n5545 = ~n2554 ;
  assign n2770 = n5545 & n2769 ;
  assign n5546 = ~n2769 ;
  assign n2771 = n2554 & n5546 ;
  assign n2772 = n2770 | n2771 ;
  assign n5547 = ~n2772 ;
  assign n2773 = n2767 & n5547 ;
  assign n2774 = n2766 | n2773 ;
  assign n2775 = x51 & n2774 ;
  assign n2776 = x51 | n2774 ;
  assign n2777 = n2557 & n5476 ;
  assign n2778 = n73 & n2777 ;
  assign n5548 = ~n2563 ;
  assign n2779 = n5548 & n2778 ;
  assign n5549 = ~n2778 ;
  assign n2780 = n2563 & n5549 ;
  assign n2781 = n2779 | n2780 ;
  assign n5550 = ~n2781 ;
  assign n2782 = n2776 & n5550 ;
  assign n2783 = n2775 | n2782 ;
  assign n2784 = x52 & n2783 ;
  assign n2785 = x52 | n2783 ;
  assign n2786 = n2566 & n5480 ;
  assign n2787 = n73 & n2786 ;
  assign n2788 = n2572 & n2787 ;
  assign n2789 = n2572 | n2787 ;
  assign n5551 = ~n2788 ;
  assign n2790 = n5551 & n2789 ;
  assign n5552 = ~n2790 ;
  assign n2791 = n2785 & n5552 ;
  assign n2792 = n2784 | n2791 ;
  assign n2793 = x53 & n2792 ;
  assign n2794 = x53 | n2792 ;
  assign n2795 = n2575 & n5484 ;
  assign n2796 = n73 & n2795 ;
  assign n5553 = ~n2581 ;
  assign n2797 = n5553 & n2796 ;
  assign n5554 = ~n2796 ;
  assign n2798 = n2581 & n5554 ;
  assign n2799 = n2797 | n2798 ;
  assign n5555 = ~n2799 ;
  assign n2800 = n2794 & n5555 ;
  assign n2801 = n2793 | n2800 ;
  assign n2802 = x54 & n2801 ;
  assign n2803 = x54 | n2801 ;
  assign n2804 = n2584 & n5488 ;
  assign n2805 = n73 & n2804 ;
  assign n2806 = n2590 & n2805 ;
  assign n2807 = n2590 | n2805 ;
  assign n5556 = ~n2806 ;
  assign n2808 = n5556 & n2807 ;
  assign n5557 = ~n2808 ;
  assign n2809 = n2803 & n5557 ;
  assign n2810 = n2802 | n2809 ;
  assign n2811 = x55 & n2810 ;
  assign n2812 = x55 | n2810 ;
  assign n2813 = n2593 & n5492 ;
  assign n2814 = n73 & n2813 ;
  assign n2815 = n2599 & n2814 ;
  assign n2816 = n2599 | n2814 ;
  assign n5558 = ~n2815 ;
  assign n2817 = n5558 & n2816 ;
  assign n5559 = ~n2817 ;
  assign n2818 = n2812 & n5559 ;
  assign n2819 = n2811 | n2818 ;
  assign n2820 = x56 | n2819 ;
  assign n2821 = x56 & n2819 ;
  assign n2822 = n117 | n2821 ;
  assign n5560 = ~n2822 ;
  assign n2824 = n2820 & n5560 ;
  assign n5561 = ~n2824 ;
  assign n2825 = n2606 & n5561 ;
  assign n5562 = ~x6 ;
  assign n100 = n5562 & n4602 ;
  assign n5563 = ~n2606 ;
  assign n2823 = n5563 & n2820 ;
  assign n2826 = n2822 | n2823 ;
  assign n72 = ~n2826 ;
  assign n2827 = x32 & n72 ;
  assign n2828 = n5496 & n2827 ;
  assign n5565 = ~n2827 ;
  assign n2829 = x7 & n5565 ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = n5562 & x32 ;
  assign n2832 = x33 | n2831 ;
  assign n5566 = ~n2830 ;
  assign n2833 = n5566 & n2832 ;
  assign n2834 = n100 | n2833 ;
  assign n2835 = x34 & n2834 ;
  assign n5567 = ~n99 ;
  assign n2836 = n5567 & n2614 ;
  assign n2837 = n72 & n2836 ;
  assign n2838 = n2613 & n2837 ;
  assign n2839 = n2613 | n2837 ;
  assign n5568 = ~n2838 ;
  assign n2840 = n5568 & n2839 ;
  assign n2841 = x34 | n2834 ;
  assign n5569 = ~n2840 ;
  assign n2842 = n5569 & n2841 ;
  assign n2843 = n2835 | n2842 ;
  assign n2846 = x35 | n2843 ;
  assign n2844 = x35 & n2843 ;
  assign n2847 = n2617 | n2826 ;
  assign n5570 = ~n2847 ;
  assign n2848 = n2628 & n5570 ;
  assign n2849 = x34 | n2616 ;
  assign n2850 = n5570 & n2849 ;
  assign n5571 = ~n2850 ;
  assign n2851 = n2627 & n5571 ;
  assign n2852 = n2848 | n2851 ;
  assign n5572 = ~n2844 ;
  assign n2853 = n5572 & n2852 ;
  assign n5573 = ~n2853 ;
  assign n2854 = n2846 & n5573 ;
  assign n2855 = x36 & n2854 ;
  assign n2856 = x36 | n2854 ;
  assign n5574 = ~n2630 ;
  assign n2857 = n5574 & n2631 ;
  assign n2858 = n72 & n2857 ;
  assign n2859 = n2637 & n2858 ;
  assign n2860 = n2637 | n2858 ;
  assign n5575 = ~n2859 ;
  assign n2861 = n5575 & n2860 ;
  assign n5576 = ~n2861 ;
  assign n2862 = n2856 & n5576 ;
  assign n2863 = n2855 | n2862 ;
  assign n2864 = x37 & n2863 ;
  assign n2865 = x37 | n2863 ;
  assign n5577 = ~n2640 ;
  assign n2866 = n5577 & n2641 ;
  assign n2867 = n72 & n2866 ;
  assign n2868 = n5511 & n2867 ;
  assign n5578 = ~n2867 ;
  assign n2869 = n2646 & n5578 ;
  assign n2870 = n2868 | n2869 ;
  assign n5579 = ~n2870 ;
  assign n2871 = n2865 & n5579 ;
  assign n2872 = n2864 | n2871 ;
  assign n2873 = x38 & n2872 ;
  assign n2874 = x38 | n2872 ;
  assign n5580 = ~n2649 ;
  assign n2875 = n5580 & n2650 ;
  assign n2876 = n72 & n2875 ;
  assign n2877 = n2655 & n2876 ;
  assign n2878 = n2655 | n2876 ;
  assign n5581 = ~n2877 ;
  assign n2879 = n5581 & n2878 ;
  assign n5582 = ~n2879 ;
  assign n2880 = n2874 & n5582 ;
  assign n2881 = n2873 | n2880 ;
  assign n2882 = x39 & n2881 ;
  assign n2883 = x39 | n2881 ;
  assign n5583 = ~n2658 ;
  assign n2884 = n5583 & n2659 ;
  assign n2885 = n72 & n2884 ;
  assign n2886 = n2664 & n2885 ;
  assign n2887 = n2664 | n2885 ;
  assign n5584 = ~n2886 ;
  assign n2888 = n5584 & n2887 ;
  assign n5585 = ~n2888 ;
  assign n2889 = n2883 & n5585 ;
  assign n2890 = n2882 | n2889 ;
  assign n2891 = x40 & n2890 ;
  assign n2892 = x40 | n2890 ;
  assign n5586 = ~n2667 ;
  assign n2893 = n5586 & n2668 ;
  assign n2894 = n72 & n2893 ;
  assign n2895 = n2673 & n2894 ;
  assign n2896 = n2673 | n2894 ;
  assign n5587 = ~n2895 ;
  assign n2897 = n5587 & n2896 ;
  assign n5588 = ~n2897 ;
  assign n2898 = n2892 & n5588 ;
  assign n2899 = n2891 | n2898 ;
  assign n2900 = x41 & n2899 ;
  assign n5589 = ~n2676 ;
  assign n2901 = n5589 & n2682 ;
  assign n2902 = n72 & n2901 ;
  assign n2903 = n2681 & n2902 ;
  assign n2904 = n2681 | n2902 ;
  assign n5590 = ~n2903 ;
  assign n2905 = n5590 & n2904 ;
  assign n2906 = x41 | n2899 ;
  assign n5591 = ~n2905 ;
  assign n2907 = n5591 & n2906 ;
  assign n2908 = n2900 | n2907 ;
  assign n2909 = x42 & n2908 ;
  assign n5592 = ~n2685 ;
  assign n2910 = n5592 & n2691 ;
  assign n2911 = n72 & n2910 ;
  assign n2912 = n5523 & n2911 ;
  assign n5593 = ~n2911 ;
  assign n2913 = n2690 & n5593 ;
  assign n2914 = n2912 | n2913 ;
  assign n2915 = x42 | n2908 ;
  assign n5594 = ~n2914 ;
  assign n2916 = n5594 & n2915 ;
  assign n2917 = n2909 | n2916 ;
  assign n2918 = x43 & n2917 ;
  assign n2919 = x43 | n2917 ;
  assign n5595 = ~n2694 ;
  assign n2920 = n5595 & n2695 ;
  assign n2921 = n72 & n2920 ;
  assign n2922 = n5526 & n2921 ;
  assign n5596 = ~n2921 ;
  assign n2923 = n2700 & n5596 ;
  assign n2924 = n2922 | n2923 ;
  assign n5597 = ~n2924 ;
  assign n2925 = n2919 & n5597 ;
  assign n2926 = n2918 | n2925 ;
  assign n2927 = x44 & n2926 ;
  assign n2928 = x44 | n2926 ;
  assign n5598 = ~n2703 ;
  assign n2929 = n5598 & n2704 ;
  assign n2930 = n72 & n2929 ;
  assign n2931 = n5529 & n2930 ;
  assign n5599 = ~n2930 ;
  assign n2932 = n2709 & n5599 ;
  assign n2933 = n2931 | n2932 ;
  assign n5600 = ~n2933 ;
  assign n2934 = n2928 & n5600 ;
  assign n2935 = n2927 | n2934 ;
  assign n2936 = x45 & n2935 ;
  assign n2937 = x45 | n2935 ;
  assign n5601 = ~n2712 ;
  assign n2938 = n5601 & n2713 ;
  assign n2939 = n72 & n2938 ;
  assign n2940 = n2718 & n2939 ;
  assign n2941 = n2718 | n2939 ;
  assign n5602 = ~n2940 ;
  assign n2942 = n5602 & n2941 ;
  assign n5603 = ~n2942 ;
  assign n2943 = n2937 & n5603 ;
  assign n2944 = n2936 | n2943 ;
  assign n2945 = x46 & n2944 ;
  assign n2946 = x46 | n2944 ;
  assign n5604 = ~n2721 ;
  assign n2947 = n5604 & n2722 ;
  assign n2948 = n72 & n2947 ;
  assign n2949 = n2727 & n2948 ;
  assign n2950 = n2727 | n2948 ;
  assign n5605 = ~n2949 ;
  assign n2951 = n5605 & n2950 ;
  assign n5606 = ~n2951 ;
  assign n2952 = n2946 & n5606 ;
  assign n2953 = n2945 | n2952 ;
  assign n2954 = x47 & n2953 ;
  assign n2955 = x47 | n2953 ;
  assign n5607 = ~n2730 ;
  assign n2956 = n5607 & n2731 ;
  assign n2957 = n72 & n2956 ;
  assign n2958 = n5536 & n2957 ;
  assign n5608 = ~n2957 ;
  assign n2959 = n2736 & n5608 ;
  assign n2960 = n2958 | n2959 ;
  assign n5609 = ~n2960 ;
  assign n2961 = n2955 & n5609 ;
  assign n2962 = n2954 | n2961 ;
  assign n2963 = x48 & n2962 ;
  assign n2964 = x48 | n2962 ;
  assign n5610 = ~n2739 ;
  assign n2965 = n5610 & n2740 ;
  assign n2966 = n72 & n2965 ;
  assign n2967 = n2745 & n2966 ;
  assign n2968 = n2745 | n2966 ;
  assign n5611 = ~n2967 ;
  assign n2969 = n5611 & n2968 ;
  assign n5612 = ~n2969 ;
  assign n2970 = n2964 & n5612 ;
  assign n2971 = n2963 | n2970 ;
  assign n2972 = x49 & n2971 ;
  assign n2973 = x49 | n2971 ;
  assign n5613 = ~n2748 ;
  assign n2974 = n5613 & n2749 ;
  assign n2975 = n72 & n2974 ;
  assign n2976 = n2754 & n2975 ;
  assign n2977 = n2754 | n2975 ;
  assign n5614 = ~n2976 ;
  assign n2978 = n5614 & n2977 ;
  assign n5615 = ~n2978 ;
  assign n2979 = n2973 & n5615 ;
  assign n2980 = n2972 | n2979 ;
  assign n2981 = x50 & n2980 ;
  assign n2982 = x50 | n2980 ;
  assign n5616 = ~n2757 ;
  assign n2983 = n5616 & n2758 ;
  assign n2984 = n72 & n2983 ;
  assign n2985 = n5544 & n2984 ;
  assign n5617 = ~n2984 ;
  assign n2986 = n2763 & n5617 ;
  assign n2987 = n2985 | n2986 ;
  assign n5618 = ~n2987 ;
  assign n2988 = n2982 & n5618 ;
  assign n2989 = n2981 | n2988 ;
  assign n2990 = x51 & n2989 ;
  assign n2991 = x51 | n2989 ;
  assign n5619 = ~n2766 ;
  assign n2992 = n5619 & n2767 ;
  assign n2993 = n72 & n2992 ;
  assign n2994 = n5547 & n2993 ;
  assign n5620 = ~n2993 ;
  assign n2995 = n2772 & n5620 ;
  assign n2996 = n2994 | n2995 ;
  assign n5621 = ~n2996 ;
  assign n2997 = n2991 & n5621 ;
  assign n2998 = n2990 | n2997 ;
  assign n2999 = x52 & n2998 ;
  assign n3000 = x52 | n2998 ;
  assign n5622 = ~n2775 ;
  assign n3001 = n5622 & n2776 ;
  assign n3002 = n72 & n3001 ;
  assign n3003 = n2781 & n3002 ;
  assign n3004 = n2781 | n3002 ;
  assign n5623 = ~n3003 ;
  assign n3005 = n5623 & n3004 ;
  assign n5624 = ~n3005 ;
  assign n3006 = n3000 & n5624 ;
  assign n3007 = n2999 | n3006 ;
  assign n3008 = x53 & n3007 ;
  assign n3009 = x53 | n3007 ;
  assign n5625 = ~n2784 ;
  assign n3010 = n5625 & n2785 ;
  assign n3011 = n72 & n3010 ;
  assign n3012 = n2790 & n3011 ;
  assign n3013 = n2790 | n3011 ;
  assign n5626 = ~n3012 ;
  assign n3014 = n5626 & n3013 ;
  assign n5627 = ~n3014 ;
  assign n3015 = n3009 & n5627 ;
  assign n3016 = n3008 | n3015 ;
  assign n3017 = x54 & n3016 ;
  assign n3018 = x54 | n3016 ;
  assign n5628 = ~n2793 ;
  assign n3019 = n5628 & n2794 ;
  assign n3020 = n72 & n3019 ;
  assign n3021 = n2799 & n3020 ;
  assign n3022 = n2799 | n3020 ;
  assign n5629 = ~n3021 ;
  assign n3023 = n5629 & n3022 ;
  assign n5630 = ~n3023 ;
  assign n3024 = n3018 & n5630 ;
  assign n3025 = n3017 | n3024 ;
  assign n3026 = x55 & n3025 ;
  assign n3027 = x55 | n3025 ;
  assign n5631 = ~n2802 ;
  assign n3028 = n5631 & n2803 ;
  assign n3029 = n72 & n3028 ;
  assign n3030 = n2808 & n3029 ;
  assign n3031 = n2808 | n3029 ;
  assign n5632 = ~n3030 ;
  assign n3032 = n5632 & n3031 ;
  assign n5633 = ~n3032 ;
  assign n3033 = n3027 & n5633 ;
  assign n3034 = n3026 | n3033 ;
  assign n3035 = x56 & n3034 ;
  assign n3036 = x56 | n3034 ;
  assign n5634 = ~n2811 ;
  assign n3037 = n5634 & n2812 ;
  assign n3038 = n72 & n3037 ;
  assign n3039 = n5559 & n3038 ;
  assign n5635 = ~n3038 ;
  assign n3040 = n2817 & n5635 ;
  assign n3041 = n3039 | n3040 ;
  assign n5636 = ~n3041 ;
  assign n3042 = n3036 & n5636 ;
  assign n3043 = n3035 | n3042 ;
  assign n3044 = x57 | n3043 ;
  assign n3045 = x57 & n3043 ;
  assign n3046 = n116 | n3045 ;
  assign n5637 = ~n3046 ;
  assign n3048 = n3044 & n5637 ;
  assign n5638 = ~n3048 ;
  assign n3049 = n2825 & n5638 ;
  assign n5639 = ~x5 ;
  assign n102 = n5639 & n4602 ;
  assign n5640 = ~n2825 ;
  assign n3047 = n5640 & n3044 ;
  assign n3050 = n3046 | n3047 ;
  assign n71 = ~n3050 ;
  assign n3051 = x32 & n71 ;
  assign n3052 = x6 & n3051 ;
  assign n3054 = x6 | n3051 ;
  assign n5642 = ~n3052 ;
  assign n3055 = n5642 & n3054 ;
  assign n101 = n5639 & x32 ;
  assign n3056 = x33 | n101 ;
  assign n5643 = ~n3055 ;
  assign n3057 = n5643 & n3056 ;
  assign n3058 = n102 | n3057 ;
  assign n3059 = x34 & n3058 ;
  assign n3053 = n5562 & n3051 ;
  assign n5644 = ~n3051 ;
  assign n3060 = x6 & n5644 ;
  assign n3061 = n3053 | n3060 ;
  assign n5645 = ~n3061 ;
  assign n3062 = n3056 & n5645 ;
  assign n3063 = n102 | n3062 ;
  assign n3064 = x34 | n3063 ;
  assign n5646 = ~n100 ;
  assign n3065 = n5646 & n2832 ;
  assign n3066 = n71 & n3065 ;
  assign n3067 = n5566 & n3066 ;
  assign n5647 = ~n3066 ;
  assign n3068 = n2830 & n5647 ;
  assign n3069 = n3067 | n3068 ;
  assign n5648 = ~n3069 ;
  assign n3070 = n3064 & n5648 ;
  assign n3071 = n3059 | n3070 ;
  assign n3072 = x35 & n3071 ;
  assign n3073 = x35 | n3071 ;
  assign n5649 = ~n2835 ;
  assign n3074 = n5649 & n2841 ;
  assign n3075 = n71 & n3074 ;
  assign n3076 = n2840 & n3075 ;
  assign n3077 = n2840 | n3075 ;
  assign n5650 = ~n3076 ;
  assign n3078 = n5650 & n3077 ;
  assign n5651 = ~n3078 ;
  assign n3079 = n3073 & n5651 ;
  assign n3080 = n3072 | n3079 ;
  assign n3081 = x36 & n3080 ;
  assign n3082 = x36 | n3080 ;
  assign n2845 = n5416 & n2843 ;
  assign n5652 = ~n2843 ;
  assign n3083 = x35 & n5652 ;
  assign n3084 = n2845 | n3083 ;
  assign n3085 = n71 & n3084 ;
  assign n5653 = ~n2852 ;
  assign n3086 = n5653 & n3085 ;
  assign n5654 = ~n3085 ;
  assign n3087 = n2852 & n5654 ;
  assign n3088 = n3086 | n3087 ;
  assign n5655 = ~n3088 ;
  assign n3089 = n3082 & n5655 ;
  assign n3090 = n3081 | n3089 ;
  assign n3091 = x37 & n3090 ;
  assign n3092 = x37 | n3090 ;
  assign n5656 = ~n2855 ;
  assign n3093 = n5656 & n2856 ;
  assign n3094 = n71 & n3093 ;
  assign n3095 = n2861 & n3094 ;
  assign n3096 = n2861 | n3094 ;
  assign n5657 = ~n3095 ;
  assign n3097 = n5657 & n3096 ;
  assign n5658 = ~n3097 ;
  assign n3098 = n3092 & n5658 ;
  assign n3099 = n3091 | n3098 ;
  assign n3100 = x38 & n3099 ;
  assign n3101 = x38 | n3099 ;
  assign n5659 = ~n2864 ;
  assign n3102 = n5659 & n2865 ;
  assign n3103 = n71 & n3102 ;
  assign n3104 = n2870 & n3103 ;
  assign n3105 = n2870 | n3103 ;
  assign n5660 = ~n3104 ;
  assign n3106 = n5660 & n3105 ;
  assign n5661 = ~n3106 ;
  assign n3107 = n3101 & n5661 ;
  assign n3108 = n3100 | n3107 ;
  assign n3109 = x39 & n3108 ;
  assign n3110 = x39 | n3108 ;
  assign n5662 = ~n2873 ;
  assign n3111 = n5662 & n2874 ;
  assign n3112 = n71 & n3111 ;
  assign n3113 = n2879 & n3112 ;
  assign n3114 = n2879 | n3112 ;
  assign n5663 = ~n3113 ;
  assign n3115 = n5663 & n3114 ;
  assign n5664 = ~n3115 ;
  assign n3116 = n3110 & n5664 ;
  assign n3117 = n3109 | n3116 ;
  assign n3118 = x40 & n3117 ;
  assign n3119 = x40 | n3117 ;
  assign n5665 = ~n2882 ;
  assign n3120 = n5665 & n2883 ;
  assign n3121 = n71 & n3120 ;
  assign n3122 = n5585 & n3121 ;
  assign n5666 = ~n3121 ;
  assign n3123 = n2888 & n5666 ;
  assign n3124 = n3122 | n3123 ;
  assign n5667 = ~n3124 ;
  assign n3125 = n3119 & n5667 ;
  assign n3126 = n3118 | n3125 ;
  assign n3127 = x41 & n3126 ;
  assign n3128 = x41 | n3126 ;
  assign n5668 = ~n2891 ;
  assign n3129 = n5668 & n2892 ;
  assign n3130 = n71 & n3129 ;
  assign n3131 = n2897 & n3130 ;
  assign n3132 = n2897 | n3130 ;
  assign n5669 = ~n3131 ;
  assign n3133 = n5669 & n3132 ;
  assign n5670 = ~n3133 ;
  assign n3134 = n3128 & n5670 ;
  assign n3135 = n3127 | n3134 ;
  assign n3136 = x42 & n3135 ;
  assign n5671 = ~n2900 ;
  assign n3137 = n5671 & n2906 ;
  assign n3138 = n71 & n3137 ;
  assign n3139 = n2905 & n3138 ;
  assign n3140 = n2905 | n3138 ;
  assign n5672 = ~n3139 ;
  assign n3141 = n5672 & n3140 ;
  assign n3142 = x42 | n3135 ;
  assign n5673 = ~n3141 ;
  assign n3143 = n5673 & n3142 ;
  assign n3144 = n3136 | n3143 ;
  assign n3145 = x43 & n3144 ;
  assign n3146 = x43 | n3144 ;
  assign n5674 = ~n2909 ;
  assign n3147 = n5674 & n2915 ;
  assign n3148 = n71 & n3147 ;
  assign n3149 = n5594 & n3148 ;
  assign n5675 = ~n3148 ;
  assign n3150 = n2914 & n5675 ;
  assign n3151 = n3149 | n3150 ;
  assign n5676 = ~n3151 ;
  assign n3152 = n3146 & n5676 ;
  assign n3153 = n3145 | n3152 ;
  assign n3154 = x44 & n3153 ;
  assign n3155 = x44 | n3153 ;
  assign n5677 = ~n2918 ;
  assign n3156 = n5677 & n2919 ;
  assign n3157 = n71 & n3156 ;
  assign n3158 = n2924 & n3157 ;
  assign n3159 = n2924 | n3157 ;
  assign n5678 = ~n3158 ;
  assign n3160 = n5678 & n3159 ;
  assign n5679 = ~n3160 ;
  assign n3161 = n3155 & n5679 ;
  assign n3162 = n3154 | n3161 ;
  assign n3163 = x45 & n3162 ;
  assign n3164 = x45 | n3162 ;
  assign n5680 = ~n2927 ;
  assign n3165 = n5680 & n2928 ;
  assign n3166 = n71 & n3165 ;
  assign n3167 = n5600 & n3166 ;
  assign n5681 = ~n3166 ;
  assign n3168 = n2933 & n5681 ;
  assign n3169 = n3167 | n3168 ;
  assign n5682 = ~n3169 ;
  assign n3170 = n3164 & n5682 ;
  assign n3171 = n3163 | n3170 ;
  assign n3172 = x46 & n3171 ;
  assign n3173 = x46 | n3171 ;
  assign n5683 = ~n2936 ;
  assign n3174 = n5683 & n2937 ;
  assign n3175 = n71 & n3174 ;
  assign n3176 = n2942 & n3175 ;
  assign n3177 = n2942 | n3175 ;
  assign n5684 = ~n3176 ;
  assign n3178 = n5684 & n3177 ;
  assign n5685 = ~n3178 ;
  assign n3179 = n3173 & n5685 ;
  assign n3180 = n3172 | n3179 ;
  assign n3181 = x47 & n3180 ;
  assign n3182 = x47 | n3180 ;
  assign n5686 = ~n2945 ;
  assign n3183 = n5686 & n2946 ;
  assign n3184 = n71 & n3183 ;
  assign n3185 = n2951 & n3184 ;
  assign n3186 = n2951 | n3184 ;
  assign n5687 = ~n3185 ;
  assign n3187 = n5687 & n3186 ;
  assign n5688 = ~n3187 ;
  assign n3188 = n3182 & n5688 ;
  assign n3189 = n3181 | n3188 ;
  assign n3190 = x48 & n3189 ;
  assign n3191 = x48 | n3189 ;
  assign n5689 = ~n2954 ;
  assign n3192 = n5689 & n2955 ;
  assign n3193 = n71 & n3192 ;
  assign n3194 = n5609 & n3193 ;
  assign n5690 = ~n3193 ;
  assign n3195 = n2960 & n5690 ;
  assign n3196 = n3194 | n3195 ;
  assign n5691 = ~n3196 ;
  assign n3197 = n3191 & n5691 ;
  assign n3198 = n3190 | n3197 ;
  assign n3199 = x49 & n3198 ;
  assign n3200 = x49 | n3198 ;
  assign n5692 = ~n2963 ;
  assign n3201 = n5692 & n2964 ;
  assign n3202 = n71 & n3201 ;
  assign n3203 = n2969 & n3202 ;
  assign n3204 = n2969 | n3202 ;
  assign n5693 = ~n3203 ;
  assign n3205 = n5693 & n3204 ;
  assign n5694 = ~n3205 ;
  assign n3206 = n3200 & n5694 ;
  assign n3207 = n3199 | n3206 ;
  assign n3208 = x50 & n3207 ;
  assign n3209 = x50 | n3207 ;
  assign n5695 = ~n2972 ;
  assign n3210 = n5695 & n2973 ;
  assign n3211 = n71 & n3210 ;
  assign n3212 = n2978 & n3211 ;
  assign n3213 = n2978 | n3211 ;
  assign n5696 = ~n3212 ;
  assign n3214 = n5696 & n3213 ;
  assign n5697 = ~n3214 ;
  assign n3215 = n3209 & n5697 ;
  assign n3216 = n3208 | n3215 ;
  assign n3217 = x51 & n3216 ;
  assign n3218 = x51 | n3216 ;
  assign n5698 = ~n2981 ;
  assign n3219 = n5698 & n2982 ;
  assign n3220 = n71 & n3219 ;
  assign n3221 = n2987 & n3220 ;
  assign n3222 = n2987 | n3220 ;
  assign n5699 = ~n3221 ;
  assign n3223 = n5699 & n3222 ;
  assign n5700 = ~n3223 ;
  assign n3224 = n3218 & n5700 ;
  assign n3225 = n3217 | n3224 ;
  assign n3226 = x52 & n3225 ;
  assign n3227 = x52 | n3225 ;
  assign n5701 = ~n2990 ;
  assign n3228 = n5701 & n2991 ;
  assign n3229 = n71 & n3228 ;
  assign n3230 = n5621 & n3229 ;
  assign n5702 = ~n3229 ;
  assign n3231 = n2996 & n5702 ;
  assign n3232 = n3230 | n3231 ;
  assign n5703 = ~n3232 ;
  assign n3233 = n3227 & n5703 ;
  assign n3234 = n3226 | n3233 ;
  assign n3235 = x53 & n3234 ;
  assign n3236 = x53 | n3234 ;
  assign n5704 = ~n2999 ;
  assign n3237 = n5704 & n3000 ;
  assign n3238 = n71 & n3237 ;
  assign n3239 = n3005 & n3238 ;
  assign n3240 = n3005 | n3238 ;
  assign n5705 = ~n3239 ;
  assign n3241 = n5705 & n3240 ;
  assign n5706 = ~n3241 ;
  assign n3242 = n3236 & n5706 ;
  assign n3243 = n3235 | n3242 ;
  assign n3244 = x54 & n3243 ;
  assign n3245 = x54 | n3243 ;
  assign n5707 = ~n3008 ;
  assign n3246 = n5707 & n3009 ;
  assign n3247 = n71 & n3246 ;
  assign n3248 = n3014 & n3247 ;
  assign n3249 = n3014 | n3247 ;
  assign n5708 = ~n3248 ;
  assign n3250 = n5708 & n3249 ;
  assign n5709 = ~n3250 ;
  assign n3251 = n3245 & n5709 ;
  assign n3252 = n3244 | n3251 ;
  assign n3253 = x55 & n3252 ;
  assign n3254 = x55 | n3252 ;
  assign n5710 = ~n3017 ;
  assign n3255 = n5710 & n3018 ;
  assign n3256 = n71 & n3255 ;
  assign n3257 = n3023 & n3256 ;
  assign n3258 = n3023 | n3256 ;
  assign n5711 = ~n3257 ;
  assign n3259 = n5711 & n3258 ;
  assign n5712 = ~n3259 ;
  assign n3260 = n3254 & n5712 ;
  assign n3261 = n3253 | n3260 ;
  assign n3262 = x56 & n3261 ;
  assign n3263 = x56 | n3261 ;
  assign n5713 = ~n3026 ;
  assign n3264 = n5713 & n3027 ;
  assign n3265 = n71 & n3264 ;
  assign n3266 = n3032 & n3265 ;
  assign n3267 = n3032 | n3265 ;
  assign n5714 = ~n3266 ;
  assign n3268 = n5714 & n3267 ;
  assign n5715 = ~n3268 ;
  assign n3269 = n3263 & n5715 ;
  assign n3270 = n3262 | n3269 ;
  assign n3271 = x57 & n3270 ;
  assign n3272 = x57 | n3270 ;
  assign n5716 = ~n3035 ;
  assign n3273 = n5716 & n3036 ;
  assign n3274 = n71 & n3273 ;
  assign n3275 = n5636 & n3274 ;
  assign n5717 = ~n3274 ;
  assign n3276 = n3041 & n5717 ;
  assign n3277 = n3275 | n3276 ;
  assign n5718 = ~n3277 ;
  assign n3278 = n3272 & n5718 ;
  assign n3279 = n3271 | n3278 ;
  assign n3280 = x58 | n3279 ;
  assign n3281 = x58 & n3279 ;
  assign n3282 = n115 | n3281 ;
  assign n5719 = ~n3282 ;
  assign n3284 = n3280 & n5719 ;
  assign n5720 = ~n3284 ;
  assign n3285 = n3049 & n5720 ;
  assign n5721 = ~x4 ;
  assign n104 = n5721 & n4602 ;
  assign n5722 = ~n3049 ;
  assign n3283 = n5722 & n3280 ;
  assign n3286 = n3282 | n3283 ;
  assign n70 = ~n3286 ;
  assign n3287 = x32 & n70 ;
  assign n3288 = x5 & n3287 ;
  assign n3290 = x5 | n3287 ;
  assign n5724 = ~n3288 ;
  assign n3291 = n5724 & n3290 ;
  assign n103 = n5721 & x32 ;
  assign n3292 = x33 | n103 ;
  assign n5725 = ~n3291 ;
  assign n3293 = n5725 & n3292 ;
  assign n3294 = n104 | n3293 ;
  assign n3295 = x34 & n3294 ;
  assign n3289 = n5639 & n3287 ;
  assign n5726 = ~n3287 ;
  assign n3296 = x5 & n5726 ;
  assign n3297 = n3289 | n3296 ;
  assign n5727 = ~n3297 ;
  assign n3298 = n3292 & n5727 ;
  assign n3299 = n104 | n3298 ;
  assign n3300 = x34 | n3299 ;
  assign n5728 = ~n102 ;
  assign n3301 = n5728 & n3056 ;
  assign n3302 = n70 & n3301 ;
  assign n3303 = n3055 & n3302 ;
  assign n3304 = n3055 | n3302 ;
  assign n5729 = ~n3303 ;
  assign n3305 = n5729 & n3304 ;
  assign n5730 = ~n3305 ;
  assign n3306 = n3300 & n5730 ;
  assign n3307 = n3295 | n3306 ;
  assign n3308 = x35 & n3307 ;
  assign n3309 = x35 | n3307 ;
  assign n3310 = x34 | n3058 ;
  assign n3311 = n3059 | n3286 ;
  assign n5731 = ~n3311 ;
  assign n3312 = n3310 & n5731 ;
  assign n5732 = ~n3312 ;
  assign n3313 = n3069 & n5732 ;
  assign n3314 = n3070 & n5731 ;
  assign n3315 = n3313 | n3314 ;
  assign n5733 = ~n3315 ;
  assign n3316 = n3309 & n5733 ;
  assign n3317 = n3308 | n3316 ;
  assign n3318 = x36 & n3317 ;
  assign n3319 = x36 | n3317 ;
  assign n5734 = ~n3072 ;
  assign n3320 = n5734 & n3073 ;
  assign n3321 = n70 & n3320 ;
  assign n3322 = n3078 & n3321 ;
  assign n3323 = n3078 | n3321 ;
  assign n5735 = ~n3322 ;
  assign n3324 = n5735 & n3323 ;
  assign n5736 = ~n3324 ;
  assign n3325 = n3319 & n5736 ;
  assign n3326 = n3318 | n3325 ;
  assign n3327 = x37 & n3326 ;
  assign n3328 = x37 | n3326 ;
  assign n5737 = ~n3081 ;
  assign n3329 = n5737 & n3082 ;
  assign n3330 = n70 & n3329 ;
  assign n3331 = n3088 & n3330 ;
  assign n3332 = n3088 | n3330 ;
  assign n5738 = ~n3331 ;
  assign n3333 = n5738 & n3332 ;
  assign n5739 = ~n3333 ;
  assign n3334 = n3328 & n5739 ;
  assign n3335 = n3327 | n3334 ;
  assign n3336 = x38 & n3335 ;
  assign n3337 = x38 | n3335 ;
  assign n5740 = ~n3091 ;
  assign n3338 = n5740 & n3092 ;
  assign n3339 = n70 & n3338 ;
  assign n3340 = n3097 & n3339 ;
  assign n3341 = n3097 | n3339 ;
  assign n5741 = ~n3340 ;
  assign n3342 = n5741 & n3341 ;
  assign n5742 = ~n3342 ;
  assign n3343 = n3337 & n5742 ;
  assign n3344 = n3336 | n3343 ;
  assign n3345 = x39 & n3344 ;
  assign n3346 = x39 | n3344 ;
  assign n5743 = ~n3100 ;
  assign n3347 = n5743 & n3101 ;
  assign n3348 = n70 & n3347 ;
  assign n3349 = n3106 & n3348 ;
  assign n3350 = n3106 | n3348 ;
  assign n5744 = ~n3349 ;
  assign n3351 = n5744 & n3350 ;
  assign n5745 = ~n3351 ;
  assign n3352 = n3346 & n5745 ;
  assign n3353 = n3345 | n3352 ;
  assign n3354 = x40 & n3353 ;
  assign n3355 = x40 | n3353 ;
  assign n5746 = ~n3109 ;
  assign n3356 = n5746 & n3110 ;
  assign n3357 = n70 & n3356 ;
  assign n3358 = n3115 & n3357 ;
  assign n3359 = n3115 | n3357 ;
  assign n5747 = ~n3358 ;
  assign n3360 = n5747 & n3359 ;
  assign n5748 = ~n3360 ;
  assign n3361 = n3355 & n5748 ;
  assign n3362 = n3354 | n3361 ;
  assign n3363 = x41 & n3362 ;
  assign n3364 = x41 | n3362 ;
  assign n5749 = ~n3118 ;
  assign n3365 = n5749 & n3119 ;
  assign n3366 = n70 & n3365 ;
  assign n3367 = n5667 & n3366 ;
  assign n5750 = ~n3366 ;
  assign n3368 = n3124 & n5750 ;
  assign n3369 = n3367 | n3368 ;
  assign n5751 = ~n3369 ;
  assign n3370 = n3364 & n5751 ;
  assign n3371 = n3363 | n3370 ;
  assign n3372 = x42 & n3371 ;
  assign n3373 = x42 | n3371 ;
  assign n5752 = ~n3127 ;
  assign n3374 = n5752 & n3128 ;
  assign n3375 = n70 & n3374 ;
  assign n3376 = n3133 & n3375 ;
  assign n3377 = n3133 | n3375 ;
  assign n5753 = ~n3376 ;
  assign n3378 = n5753 & n3377 ;
  assign n5754 = ~n3378 ;
  assign n3379 = n3373 & n5754 ;
  assign n3380 = n3372 | n3379 ;
  assign n3381 = x43 & n3380 ;
  assign n5755 = ~n3136 ;
  assign n3382 = n5755 & n3142 ;
  assign n3383 = n70 & n3382 ;
  assign n3384 = n3141 & n3383 ;
  assign n3385 = n3141 | n3383 ;
  assign n5756 = ~n3384 ;
  assign n3386 = n5756 & n3385 ;
  assign n3387 = x43 | n3380 ;
  assign n5757 = ~n3386 ;
  assign n3388 = n5757 & n3387 ;
  assign n3389 = n3381 | n3388 ;
  assign n3390 = x44 & n3389 ;
  assign n5758 = ~n3145 ;
  assign n3391 = n5758 & n3146 ;
  assign n3392 = n70 & n3391 ;
  assign n3393 = n3151 & n3392 ;
  assign n3394 = n3151 | n3392 ;
  assign n5759 = ~n3393 ;
  assign n3395 = n5759 & n3394 ;
  assign n3396 = x44 | n3389 ;
  assign n5760 = ~n3395 ;
  assign n3397 = n5760 & n3396 ;
  assign n3398 = n3390 | n3397 ;
  assign n3399 = x45 & n3398 ;
  assign n3400 = x45 | n3398 ;
  assign n5761 = ~n3154 ;
  assign n3401 = n5761 & n3155 ;
  assign n3402 = n70 & n3401 ;
  assign n3403 = n3160 & n3402 ;
  assign n3404 = n3160 | n3402 ;
  assign n5762 = ~n3403 ;
  assign n3405 = n5762 & n3404 ;
  assign n5763 = ~n3405 ;
  assign n3406 = n3400 & n5763 ;
  assign n3407 = n3399 | n3406 ;
  assign n3408 = x46 & n3407 ;
  assign n3409 = x46 | n3407 ;
  assign n5764 = ~n3163 ;
  assign n3410 = n5764 & n3164 ;
  assign n3411 = n70 & n3410 ;
  assign n3412 = n3169 & n3411 ;
  assign n3413 = n3169 | n3411 ;
  assign n5765 = ~n3412 ;
  assign n3414 = n5765 & n3413 ;
  assign n5766 = ~n3414 ;
  assign n3415 = n3409 & n5766 ;
  assign n3416 = n3408 | n3415 ;
  assign n3417 = x47 & n3416 ;
  assign n3418 = x47 | n3416 ;
  assign n5767 = ~n3172 ;
  assign n3419 = n5767 & n3173 ;
  assign n3420 = n70 & n3419 ;
  assign n3421 = n3178 & n3420 ;
  assign n3422 = n3178 | n3420 ;
  assign n5768 = ~n3421 ;
  assign n3423 = n5768 & n3422 ;
  assign n5769 = ~n3423 ;
  assign n3424 = n3418 & n5769 ;
  assign n3425 = n3417 | n3424 ;
  assign n3426 = x48 & n3425 ;
  assign n3427 = x48 | n3425 ;
  assign n5770 = ~n3181 ;
  assign n3428 = n5770 & n3182 ;
  assign n3429 = n70 & n3428 ;
  assign n3430 = n5688 & n3429 ;
  assign n5771 = ~n3429 ;
  assign n3431 = n3187 & n5771 ;
  assign n3432 = n3430 | n3431 ;
  assign n5772 = ~n3432 ;
  assign n3433 = n3427 & n5772 ;
  assign n3434 = n3426 | n3433 ;
  assign n3435 = x49 & n3434 ;
  assign n3436 = x49 | n3434 ;
  assign n5773 = ~n3190 ;
  assign n3437 = n5773 & n3191 ;
  assign n3438 = n70 & n3437 ;
  assign n3439 = n5691 & n3438 ;
  assign n5774 = ~n3438 ;
  assign n3440 = n3196 & n5774 ;
  assign n3441 = n3439 | n3440 ;
  assign n5775 = ~n3441 ;
  assign n3442 = n3436 & n5775 ;
  assign n3443 = n3435 | n3442 ;
  assign n3444 = x50 & n3443 ;
  assign n3445 = x50 | n3443 ;
  assign n5776 = ~n3199 ;
  assign n3446 = n5776 & n3200 ;
  assign n3447 = n70 & n3446 ;
  assign n3448 = n3205 & n3447 ;
  assign n3449 = n3205 | n3447 ;
  assign n5777 = ~n3448 ;
  assign n3450 = n5777 & n3449 ;
  assign n5778 = ~n3450 ;
  assign n3451 = n3445 & n5778 ;
  assign n3452 = n3444 | n3451 ;
  assign n3453 = x51 & n3452 ;
  assign n3454 = x51 | n3452 ;
  assign n5779 = ~n3208 ;
  assign n3455 = n5779 & n3209 ;
  assign n3456 = n70 & n3455 ;
  assign n3457 = n3214 & n3456 ;
  assign n3458 = n3214 | n3456 ;
  assign n5780 = ~n3457 ;
  assign n3459 = n5780 & n3458 ;
  assign n5781 = ~n3459 ;
  assign n3460 = n3454 & n5781 ;
  assign n3461 = n3453 | n3460 ;
  assign n3462 = x52 & n3461 ;
  assign n3463 = x52 | n3461 ;
  assign n5782 = ~n3217 ;
  assign n3464 = n5782 & n3218 ;
  assign n3465 = n70 & n3464 ;
  assign n3466 = n3223 & n3465 ;
  assign n3467 = n3223 | n3465 ;
  assign n5783 = ~n3466 ;
  assign n3468 = n5783 & n3467 ;
  assign n5784 = ~n3468 ;
  assign n3469 = n3463 & n5784 ;
  assign n3470 = n3462 | n3469 ;
  assign n3471 = x53 & n3470 ;
  assign n3472 = x53 | n3470 ;
  assign n5785 = ~n3226 ;
  assign n3473 = n5785 & n3227 ;
  assign n3474 = n70 & n3473 ;
  assign n3475 = n3232 & n3474 ;
  assign n3476 = n3232 | n3474 ;
  assign n5786 = ~n3475 ;
  assign n3477 = n5786 & n3476 ;
  assign n5787 = ~n3477 ;
  assign n3478 = n3472 & n5787 ;
  assign n3479 = n3471 | n3478 ;
  assign n3480 = x54 & n3479 ;
  assign n3481 = x54 | n3479 ;
  assign n5788 = ~n3235 ;
  assign n3482 = n5788 & n3236 ;
  assign n3483 = n70 & n3482 ;
  assign n3484 = n3241 & n3483 ;
  assign n3485 = n3241 | n3483 ;
  assign n5789 = ~n3484 ;
  assign n3486 = n5789 & n3485 ;
  assign n5790 = ~n3486 ;
  assign n3487 = n3481 & n5790 ;
  assign n3488 = n3480 | n3487 ;
  assign n3489 = x55 & n3488 ;
  assign n3490 = x55 | n3488 ;
  assign n5791 = ~n3244 ;
  assign n3491 = n5791 & n3245 ;
  assign n3492 = n70 & n3491 ;
  assign n3493 = n3250 & n3492 ;
  assign n3494 = n3250 | n3492 ;
  assign n5792 = ~n3493 ;
  assign n3495 = n5792 & n3494 ;
  assign n5793 = ~n3495 ;
  assign n3496 = n3490 & n5793 ;
  assign n3497 = n3489 | n3496 ;
  assign n3498 = x56 & n3497 ;
  assign n3499 = x56 | n3497 ;
  assign n5794 = ~n3253 ;
  assign n3500 = n5794 & n3254 ;
  assign n3501 = n70 & n3500 ;
  assign n3502 = n3259 & n3501 ;
  assign n3503 = n3259 | n3501 ;
  assign n5795 = ~n3502 ;
  assign n3504 = n5795 & n3503 ;
  assign n5796 = ~n3504 ;
  assign n3505 = n3499 & n5796 ;
  assign n3506 = n3498 | n3505 ;
  assign n3507 = x57 & n3506 ;
  assign n3508 = x57 | n3506 ;
  assign n5797 = ~n3262 ;
  assign n3509 = n5797 & n3263 ;
  assign n3510 = n70 & n3509 ;
  assign n3511 = n3268 & n3510 ;
  assign n3512 = n3268 | n3510 ;
  assign n5798 = ~n3511 ;
  assign n3513 = n5798 & n3512 ;
  assign n5799 = ~n3513 ;
  assign n3514 = n3508 & n5799 ;
  assign n3515 = n3507 | n3514 ;
  assign n3516 = x58 & n3515 ;
  assign n3517 = x58 | n3515 ;
  assign n5800 = ~n3271 ;
  assign n3518 = n5800 & n3272 ;
  assign n3519 = n70 & n3518 ;
  assign n3520 = n5718 & n3519 ;
  assign n5801 = ~n3519 ;
  assign n3521 = n3277 & n5801 ;
  assign n3522 = n3520 | n3521 ;
  assign n5802 = ~n3522 ;
  assign n3523 = n3517 & n5802 ;
  assign n3524 = n3516 | n3523 ;
  assign n3525 = x59 & n3524 ;
  assign n3526 = n114 | n3525 ;
  assign n3527 = x59 | n3524 ;
  assign n5803 = ~n3526 ;
  assign n3528 = n5803 & n3527 ;
  assign n5804 = ~n3528 ;
  assign n3529 = n3285 & n5804 ;
  assign n5805 = ~x3 ;
  assign n105 = n5805 & n4602 ;
  assign n5806 = ~n3285 ;
  assign n3531 = n5806 & n3527 ;
  assign n3532 = n3526 | n3531 ;
  assign n69 = ~n3532 ;
  assign n3533 = x32 & n69 ;
  assign n3534 = n5721 & n3533 ;
  assign n5808 = ~n3533 ;
  assign n3535 = x4 & n5808 ;
  assign n3536 = n3534 | n3535 ;
  assign n3537 = n5805 & x32 ;
  assign n3538 = x33 | n3537 ;
  assign n5809 = ~n3536 ;
  assign n3539 = n5809 & n3538 ;
  assign n3540 = n105 | n3539 ;
  assign n3541 = x34 & n3540 ;
  assign n5810 = ~n104 ;
  assign n3542 = n5810 & n3292 ;
  assign n3543 = n69 & n3542 ;
  assign n3544 = n3291 & n3543 ;
  assign n3545 = n3291 | n3543 ;
  assign n5811 = ~n3544 ;
  assign n3546 = n5811 & n3545 ;
  assign n3547 = x34 | n3540 ;
  assign n5812 = ~n3546 ;
  assign n3548 = n5812 & n3547 ;
  assign n3549 = n3541 | n3548 ;
  assign n3552 = x35 | n3549 ;
  assign n3550 = x35 & n3549 ;
  assign n3553 = n3295 | n3532 ;
  assign n5813 = ~n3553 ;
  assign n3554 = n3306 & n5813 ;
  assign n3555 = x34 | n3294 ;
  assign n3556 = n5813 & n3555 ;
  assign n5814 = ~n3556 ;
  assign n3557 = n3305 & n5814 ;
  assign n3558 = n3554 | n3557 ;
  assign n5815 = ~n3550 ;
  assign n3559 = n5815 & n3558 ;
  assign n5816 = ~n3559 ;
  assign n3560 = n3552 & n5816 ;
  assign n3561 = x36 & n3560 ;
  assign n3562 = x36 | n3560 ;
  assign n5817 = ~n3308 ;
  assign n3563 = n5817 & n3309 ;
  assign n3564 = n69 & n3563 ;
  assign n3565 = n3315 & n3564 ;
  assign n3566 = n3315 | n3564 ;
  assign n5818 = ~n3565 ;
  assign n3567 = n5818 & n3566 ;
  assign n5819 = ~n3567 ;
  assign n3568 = n3562 & n5819 ;
  assign n3569 = n3561 | n3568 ;
  assign n3570 = x37 & n3569 ;
  assign n3571 = x37 | n3569 ;
  assign n5820 = ~n3318 ;
  assign n3572 = n5820 & n3319 ;
  assign n3573 = n69 & n3572 ;
  assign n3574 = n3324 & n3573 ;
  assign n3575 = n3324 | n3573 ;
  assign n5821 = ~n3574 ;
  assign n3576 = n5821 & n3575 ;
  assign n5822 = ~n3576 ;
  assign n3577 = n3571 & n5822 ;
  assign n3578 = n3570 | n3577 ;
  assign n3579 = x38 & n3578 ;
  assign n3580 = x38 | n3578 ;
  assign n5823 = ~n3327 ;
  assign n3581 = n5823 & n3328 ;
  assign n3582 = n69 & n3581 ;
  assign n3583 = n3333 & n3582 ;
  assign n3584 = n3333 | n3582 ;
  assign n5824 = ~n3583 ;
  assign n3585 = n5824 & n3584 ;
  assign n5825 = ~n3585 ;
  assign n3586 = n3580 & n5825 ;
  assign n3587 = n3579 | n3586 ;
  assign n3588 = x39 & n3587 ;
  assign n3589 = x39 | n3587 ;
  assign n5826 = ~n3336 ;
  assign n3590 = n5826 & n3337 ;
  assign n3591 = n69 & n3590 ;
  assign n3592 = n3342 & n3591 ;
  assign n3593 = n3342 | n3591 ;
  assign n5827 = ~n3592 ;
  assign n3594 = n5827 & n3593 ;
  assign n5828 = ~n3594 ;
  assign n3595 = n3589 & n5828 ;
  assign n3596 = n3588 | n3595 ;
  assign n3597 = x40 & n3596 ;
  assign n3598 = x40 | n3596 ;
  assign n5829 = ~n3345 ;
  assign n3599 = n5829 & n3346 ;
  assign n3600 = n69 & n3599 ;
  assign n3601 = n3351 & n3600 ;
  assign n3602 = n3351 | n3600 ;
  assign n5830 = ~n3601 ;
  assign n3603 = n5830 & n3602 ;
  assign n5831 = ~n3603 ;
  assign n3604 = n3598 & n5831 ;
  assign n3605 = n3597 | n3604 ;
  assign n3606 = x41 & n3605 ;
  assign n3607 = x41 | n3605 ;
  assign n5832 = ~n3354 ;
  assign n3608 = n5832 & n3355 ;
  assign n3609 = n69 & n3608 ;
  assign n3610 = n3360 & n3609 ;
  assign n3611 = n3360 | n3609 ;
  assign n5833 = ~n3610 ;
  assign n3612 = n5833 & n3611 ;
  assign n5834 = ~n3612 ;
  assign n3613 = n3607 & n5834 ;
  assign n3614 = n3606 | n3613 ;
  assign n3615 = x42 & n3614 ;
  assign n3616 = x42 | n3614 ;
  assign n5835 = ~n3363 ;
  assign n3617 = n5835 & n3364 ;
  assign n3618 = n69 & n3617 ;
  assign n3619 = n5751 & n3618 ;
  assign n5836 = ~n3618 ;
  assign n3620 = n3369 & n5836 ;
  assign n3621 = n3619 | n3620 ;
  assign n5837 = ~n3621 ;
  assign n3622 = n3616 & n5837 ;
  assign n3623 = n3615 | n3622 ;
  assign n3624 = x43 & n3623 ;
  assign n3625 = x43 | n3623 ;
  assign n5838 = ~n3372 ;
  assign n3626 = n5838 & n3373 ;
  assign n3627 = n69 & n3626 ;
  assign n3628 = n3378 & n3627 ;
  assign n3629 = n3378 | n3627 ;
  assign n5839 = ~n3628 ;
  assign n3630 = n5839 & n3629 ;
  assign n5840 = ~n3630 ;
  assign n3631 = n3625 & n5840 ;
  assign n3632 = n3624 | n3631 ;
  assign n3633 = x44 & n3632 ;
  assign n5841 = ~n3381 ;
  assign n3634 = n5841 & n3387 ;
  assign n3635 = n69 & n3634 ;
  assign n3636 = n3386 & n3635 ;
  assign n3637 = n3386 | n3635 ;
  assign n5842 = ~n3636 ;
  assign n3638 = n5842 & n3637 ;
  assign n3639 = x44 | n3632 ;
  assign n5843 = ~n3638 ;
  assign n3640 = n5843 & n3639 ;
  assign n3641 = n3633 | n3640 ;
  assign n3642 = x45 & n3641 ;
  assign n5844 = ~n3390 ;
  assign n3643 = n5844 & n3396 ;
  assign n3644 = n69 & n3643 ;
  assign n3645 = n3395 & n3644 ;
  assign n3646 = n3395 | n3644 ;
  assign n5845 = ~n3645 ;
  assign n3647 = n5845 & n3646 ;
  assign n3648 = x45 | n3641 ;
  assign n5846 = ~n3647 ;
  assign n3649 = n5846 & n3648 ;
  assign n3650 = n3642 | n3649 ;
  assign n3651 = x46 & n3650 ;
  assign n3652 = x46 | n3650 ;
  assign n5847 = ~n3399 ;
  assign n3653 = n5847 & n3400 ;
  assign n3654 = n69 & n3653 ;
  assign n3655 = n3405 & n3654 ;
  assign n3656 = n3405 | n3654 ;
  assign n5848 = ~n3655 ;
  assign n3657 = n5848 & n3656 ;
  assign n5849 = ~n3657 ;
  assign n3658 = n3652 & n5849 ;
  assign n3659 = n3651 | n3658 ;
  assign n3660 = x47 & n3659 ;
  assign n3661 = x47 | n3659 ;
  assign n5850 = ~n3408 ;
  assign n3662 = n5850 & n3409 ;
  assign n3663 = n69 & n3662 ;
  assign n3664 = n3414 & n3663 ;
  assign n3665 = n3414 | n3663 ;
  assign n5851 = ~n3664 ;
  assign n3666 = n5851 & n3665 ;
  assign n5852 = ~n3666 ;
  assign n3667 = n3661 & n5852 ;
  assign n3668 = n3660 | n3667 ;
  assign n3669 = x48 & n3668 ;
  assign n3670 = x48 | n3668 ;
  assign n5853 = ~n3417 ;
  assign n3671 = n5853 & n3418 ;
  assign n3672 = n69 & n3671 ;
  assign n3673 = n3423 & n3672 ;
  assign n3674 = n3423 | n3672 ;
  assign n5854 = ~n3673 ;
  assign n3675 = n5854 & n3674 ;
  assign n5855 = ~n3675 ;
  assign n3676 = n3670 & n5855 ;
  assign n3677 = n3669 | n3676 ;
  assign n3678 = x49 & n3677 ;
  assign n3679 = x49 | n3677 ;
  assign n5856 = ~n3426 ;
  assign n3680 = n5856 & n3427 ;
  assign n3681 = n69 & n3680 ;
  assign n3682 = n5772 & n3681 ;
  assign n5857 = ~n3681 ;
  assign n3683 = n3432 & n5857 ;
  assign n3684 = n3682 | n3683 ;
  assign n5858 = ~n3684 ;
  assign n3685 = n3679 & n5858 ;
  assign n3686 = n3678 | n3685 ;
  assign n3687 = x50 & n3686 ;
  assign n3688 = x50 | n3686 ;
  assign n5859 = ~n3435 ;
  assign n3689 = n5859 & n3436 ;
  assign n3690 = n69 & n3689 ;
  assign n3691 = n3441 & n3690 ;
  assign n3692 = n3441 | n3690 ;
  assign n5860 = ~n3691 ;
  assign n3693 = n5860 & n3692 ;
  assign n5861 = ~n3693 ;
  assign n3694 = n3688 & n5861 ;
  assign n3695 = n3687 | n3694 ;
  assign n3696 = x51 & n3695 ;
  assign n3697 = x51 | n3695 ;
  assign n5862 = ~n3444 ;
  assign n3698 = n5862 & n3445 ;
  assign n3699 = n69 & n3698 ;
  assign n3700 = n3450 & n3699 ;
  assign n3701 = n3450 | n3699 ;
  assign n5863 = ~n3700 ;
  assign n3702 = n5863 & n3701 ;
  assign n5864 = ~n3702 ;
  assign n3703 = n3697 & n5864 ;
  assign n3704 = n3696 | n3703 ;
  assign n3705 = x52 & n3704 ;
  assign n3706 = x52 | n3704 ;
  assign n5865 = ~n3453 ;
  assign n3707 = n5865 & n3454 ;
  assign n3708 = n69 & n3707 ;
  assign n3709 = n3459 & n3708 ;
  assign n3710 = n3459 | n3708 ;
  assign n5866 = ~n3709 ;
  assign n3711 = n5866 & n3710 ;
  assign n5867 = ~n3711 ;
  assign n3712 = n3706 & n5867 ;
  assign n3713 = n3705 | n3712 ;
  assign n3714 = x53 & n3713 ;
  assign n3715 = x53 | n3713 ;
  assign n5868 = ~n3462 ;
  assign n3716 = n5868 & n3463 ;
  assign n3717 = n69 & n3716 ;
  assign n3718 = n3468 & n3717 ;
  assign n3719 = n3468 | n3717 ;
  assign n5869 = ~n3718 ;
  assign n3720 = n5869 & n3719 ;
  assign n5870 = ~n3720 ;
  assign n3721 = n3715 & n5870 ;
  assign n3722 = n3714 | n3721 ;
  assign n3723 = x54 & n3722 ;
  assign n3724 = x54 | n3722 ;
  assign n5871 = ~n3471 ;
  assign n3725 = n5871 & n3472 ;
  assign n3726 = n69 & n3725 ;
  assign n3727 = n3477 & n3726 ;
  assign n3728 = n3477 | n3726 ;
  assign n5872 = ~n3727 ;
  assign n3729 = n5872 & n3728 ;
  assign n5873 = ~n3729 ;
  assign n3730 = n3724 & n5873 ;
  assign n3731 = n3723 | n3730 ;
  assign n3732 = x55 & n3731 ;
  assign n3733 = x55 | n3731 ;
  assign n5874 = ~n3480 ;
  assign n3734 = n5874 & n3481 ;
  assign n3735 = n69 & n3734 ;
  assign n3736 = n3486 & n3735 ;
  assign n3737 = n3486 | n3735 ;
  assign n5875 = ~n3736 ;
  assign n3738 = n5875 & n3737 ;
  assign n5876 = ~n3738 ;
  assign n3739 = n3733 & n5876 ;
  assign n3740 = n3732 | n3739 ;
  assign n3741 = x56 & n3740 ;
  assign n3742 = x56 | n3740 ;
  assign n5877 = ~n3489 ;
  assign n3743 = n5877 & n3490 ;
  assign n3744 = n69 & n3743 ;
  assign n3745 = n3495 & n3744 ;
  assign n3746 = n3495 | n3744 ;
  assign n5878 = ~n3745 ;
  assign n3747 = n5878 & n3746 ;
  assign n5879 = ~n3747 ;
  assign n3748 = n3742 & n5879 ;
  assign n3749 = n3741 | n3748 ;
  assign n3750 = x57 & n3749 ;
  assign n3751 = x57 | n3749 ;
  assign n5880 = ~n3498 ;
  assign n3752 = n5880 & n3499 ;
  assign n3753 = n69 & n3752 ;
  assign n3754 = n3504 & n3753 ;
  assign n3755 = n3504 | n3753 ;
  assign n5881 = ~n3754 ;
  assign n3756 = n5881 & n3755 ;
  assign n5882 = ~n3756 ;
  assign n3757 = n3751 & n5882 ;
  assign n3758 = n3750 | n3757 ;
  assign n3759 = x58 & n3758 ;
  assign n3760 = x58 | n3758 ;
  assign n5883 = ~n3507 ;
  assign n3761 = n5883 & n3508 ;
  assign n3762 = n69 & n3761 ;
  assign n3763 = n5799 & n3762 ;
  assign n5884 = ~n3762 ;
  assign n3764 = n3513 & n5884 ;
  assign n3765 = n3763 | n3764 ;
  assign n5885 = ~n3765 ;
  assign n3766 = n3760 & n5885 ;
  assign n3767 = n3759 | n3766 ;
  assign n3768 = x59 & n3767 ;
  assign n3769 = x59 | n3767 ;
  assign n5886 = ~n3516 ;
  assign n3770 = n5886 & n3517 ;
  assign n3771 = n69 & n3770 ;
  assign n3772 = n5802 & n3771 ;
  assign n5887 = ~n3771 ;
  assign n3773 = n3522 & n5887 ;
  assign n3774 = n3772 | n3773 ;
  assign n5888 = ~n3774 ;
  assign n3775 = n3769 & n5888 ;
  assign n3776 = n3768 | n3775 ;
  assign n3777 = x60 & n3776 ;
  assign n3778 = x60 | n3776 ;
  assign n5889 = ~n113 ;
  assign n3779 = n5889 & n3778 ;
  assign n5890 = ~n3777 ;
  assign n3780 = n5890 & n3779 ;
  assign n5891 = ~n3780 ;
  assign n3781 = n3529 & n5891 ;
  assign n5892 = ~x2 ;
  assign n107 = n5892 & n4602 ;
  assign n5893 = ~x60 ;
  assign n3530 = n5893 & n3529 ;
  assign n5894 = ~n3530 ;
  assign n3782 = n5894 & n3776 ;
  assign n5895 = ~n3529 ;
  assign n3783 = x60 & n5895 ;
  assign n3784 = n113 | n3783 ;
  assign n3785 = n3782 | n3784 ;
  assign n68 = ~n3785 ;
  assign n3786 = x32 & n68 ;
  assign n3787 = x3 & n3786 ;
  assign n3789 = x3 | n3786 ;
  assign n5897 = ~n3787 ;
  assign n3790 = n5897 & n3789 ;
  assign n106 = n5892 & x32 ;
  assign n3791 = x33 | n106 ;
  assign n5898 = ~n3790 ;
  assign n3792 = n5898 & n3791 ;
  assign n3793 = n107 | n3792 ;
  assign n3794 = x34 & n3793 ;
  assign n3788 = n5805 & n3786 ;
  assign n5899 = ~n3786 ;
  assign n3795 = x3 & n5899 ;
  assign n3796 = n3788 | n3795 ;
  assign n5900 = ~n3796 ;
  assign n3797 = n3791 & n5900 ;
  assign n3798 = n107 | n3797 ;
  assign n3799 = x34 | n3798 ;
  assign n5901 = ~n105 ;
  assign n3800 = n5901 & n3538 ;
  assign n3801 = n68 & n3800 ;
  assign n3802 = n5809 & n3801 ;
  assign n5902 = ~n3801 ;
  assign n3803 = n3536 & n5902 ;
  assign n3804 = n3802 | n3803 ;
  assign n5903 = ~n3804 ;
  assign n3805 = n3799 & n5903 ;
  assign n3806 = n3794 | n3805 ;
  assign n3807 = x35 & n3806 ;
  assign n3808 = x35 | n3806 ;
  assign n5904 = ~n3541 ;
  assign n3809 = n5904 & n3547 ;
  assign n3810 = n68 & n3809 ;
  assign n3811 = n3546 & n3810 ;
  assign n3812 = n3546 | n3810 ;
  assign n5905 = ~n3811 ;
  assign n3813 = n5905 & n3812 ;
  assign n5906 = ~n3813 ;
  assign n3814 = n3808 & n5906 ;
  assign n3815 = n3807 | n3814 ;
  assign n3816 = x36 & n3815 ;
  assign n3817 = x36 | n3815 ;
  assign n3551 = n5416 & n3549 ;
  assign n5907 = ~n3549 ;
  assign n3818 = x35 & n5907 ;
  assign n3819 = n3551 | n3818 ;
  assign n3820 = n68 & n3819 ;
  assign n5908 = ~n3558 ;
  assign n3821 = n5908 & n3820 ;
  assign n5909 = ~n3820 ;
  assign n3822 = n3558 & n5909 ;
  assign n3823 = n3821 | n3822 ;
  assign n5910 = ~n3823 ;
  assign n3824 = n3817 & n5910 ;
  assign n3825 = n3816 | n3824 ;
  assign n3826 = x37 & n3825 ;
  assign n3827 = x37 | n3825 ;
  assign n5911 = ~n3561 ;
  assign n3828 = n5911 & n3562 ;
  assign n3829 = n68 & n3828 ;
  assign n3830 = n3567 & n3829 ;
  assign n3831 = n3567 | n3829 ;
  assign n5912 = ~n3830 ;
  assign n3832 = n5912 & n3831 ;
  assign n5913 = ~n3832 ;
  assign n3833 = n3827 & n5913 ;
  assign n3834 = n3826 | n3833 ;
  assign n3835 = x38 & n3834 ;
  assign n3836 = x38 | n3834 ;
  assign n5914 = ~n3570 ;
  assign n3837 = n5914 & n3571 ;
  assign n3838 = n68 & n3837 ;
  assign n3839 = n3576 & n3838 ;
  assign n3840 = n3576 | n3838 ;
  assign n5915 = ~n3839 ;
  assign n3841 = n5915 & n3840 ;
  assign n5916 = ~n3841 ;
  assign n3842 = n3836 & n5916 ;
  assign n3843 = n3835 | n3842 ;
  assign n3844 = x39 & n3843 ;
  assign n3845 = x39 | n3843 ;
  assign n5917 = ~n3579 ;
  assign n3846 = n5917 & n3580 ;
  assign n3847 = n68 & n3846 ;
  assign n3848 = n3585 & n3847 ;
  assign n3849 = n3585 | n3847 ;
  assign n5918 = ~n3848 ;
  assign n3850 = n5918 & n3849 ;
  assign n5919 = ~n3850 ;
  assign n3851 = n3845 & n5919 ;
  assign n3852 = n3844 | n3851 ;
  assign n3853 = x40 & n3852 ;
  assign n3854 = x40 | n3852 ;
  assign n5920 = ~n3588 ;
  assign n3855 = n5920 & n3589 ;
  assign n3856 = n68 & n3855 ;
  assign n3857 = n3594 & n3856 ;
  assign n3858 = n3594 | n3856 ;
  assign n5921 = ~n3857 ;
  assign n3859 = n5921 & n3858 ;
  assign n5922 = ~n3859 ;
  assign n3860 = n3854 & n5922 ;
  assign n3861 = n3853 | n3860 ;
  assign n3862 = x41 & n3861 ;
  assign n3863 = x41 | n3861 ;
  assign n5923 = ~n3597 ;
  assign n3864 = n5923 & n3598 ;
  assign n3865 = n68 & n3864 ;
  assign n3866 = n3603 & n3865 ;
  assign n3867 = n3603 | n3865 ;
  assign n5924 = ~n3866 ;
  assign n3868 = n5924 & n3867 ;
  assign n5925 = ~n3868 ;
  assign n3869 = n3863 & n5925 ;
  assign n3870 = n3862 | n3869 ;
  assign n3871 = x42 & n3870 ;
  assign n3872 = x42 | n3870 ;
  assign n5926 = ~n3606 ;
  assign n3873 = n5926 & n3607 ;
  assign n3874 = n68 & n3873 ;
  assign n3875 = n3612 & n3874 ;
  assign n3876 = n3612 | n3874 ;
  assign n5927 = ~n3875 ;
  assign n3877 = n5927 & n3876 ;
  assign n5928 = ~n3877 ;
  assign n3878 = n3872 & n5928 ;
  assign n3879 = n3871 | n3878 ;
  assign n3880 = x43 & n3879 ;
  assign n3881 = x43 | n3879 ;
  assign n5929 = ~n3615 ;
  assign n3882 = n5929 & n3616 ;
  assign n3883 = n68 & n3882 ;
  assign n3884 = n3621 & n3883 ;
  assign n3885 = n3621 | n3883 ;
  assign n5930 = ~n3884 ;
  assign n3886 = n5930 & n3885 ;
  assign n5931 = ~n3886 ;
  assign n3887 = n3881 & n5931 ;
  assign n3888 = n3880 | n3887 ;
  assign n3889 = x44 & n3888 ;
  assign n3890 = x44 | n3888 ;
  assign n5932 = ~n3624 ;
  assign n3891 = n5932 & n3625 ;
  assign n3892 = n68 & n3891 ;
  assign n3893 = n5840 & n3892 ;
  assign n5933 = ~n3892 ;
  assign n3894 = n3630 & n5933 ;
  assign n3895 = n3893 | n3894 ;
  assign n5934 = ~n3895 ;
  assign n3896 = n3890 & n5934 ;
  assign n3897 = n3889 | n3896 ;
  assign n3898 = x45 & n3897 ;
  assign n5935 = ~n3633 ;
  assign n3899 = n5935 & n3639 ;
  assign n3900 = n68 & n3899 ;
  assign n3901 = n3638 & n3900 ;
  assign n3902 = n3638 | n3900 ;
  assign n5936 = ~n3901 ;
  assign n3903 = n5936 & n3902 ;
  assign n3904 = x45 | n3897 ;
  assign n5937 = ~n3903 ;
  assign n3905 = n5937 & n3904 ;
  assign n3906 = n3898 | n3905 ;
  assign n3907 = x46 & n3906 ;
  assign n3908 = x46 | n3906 ;
  assign n5938 = ~n3642 ;
  assign n3909 = n5938 & n3648 ;
  assign n3910 = n68 & n3909 ;
  assign n3911 = n3647 & n3910 ;
  assign n3912 = n3647 | n3910 ;
  assign n5939 = ~n3911 ;
  assign n3913 = n5939 & n3912 ;
  assign n5940 = ~n3913 ;
  assign n3914 = n3908 & n5940 ;
  assign n3915 = n3907 | n3914 ;
  assign n3916 = x47 & n3915 ;
  assign n3917 = x47 | n3915 ;
  assign n5941 = ~n3651 ;
  assign n3918 = n5941 & n3652 ;
  assign n3919 = n68 & n3918 ;
  assign n3920 = n3657 & n3919 ;
  assign n3921 = n3657 | n3919 ;
  assign n5942 = ~n3920 ;
  assign n3922 = n5942 & n3921 ;
  assign n5943 = ~n3922 ;
  assign n3923 = n3917 & n5943 ;
  assign n3924 = n3916 | n3923 ;
  assign n3925 = x48 & n3924 ;
  assign n3926 = x48 | n3924 ;
  assign n5944 = ~n3660 ;
  assign n3927 = n5944 & n3661 ;
  assign n3928 = n68 & n3927 ;
  assign n3929 = n3666 & n3928 ;
  assign n3930 = n3666 | n3928 ;
  assign n5945 = ~n3929 ;
  assign n3931 = n5945 & n3930 ;
  assign n5946 = ~n3931 ;
  assign n3932 = n3926 & n5946 ;
  assign n3933 = n3925 | n3932 ;
  assign n3934 = x49 & n3933 ;
  assign n3935 = x49 | n3933 ;
  assign n5947 = ~n3669 ;
  assign n3936 = n5947 & n3670 ;
  assign n3937 = n68 & n3936 ;
  assign n3938 = n3675 & n3937 ;
  assign n3939 = n3675 | n3937 ;
  assign n5948 = ~n3938 ;
  assign n3940 = n5948 & n3939 ;
  assign n5949 = ~n3940 ;
  assign n3941 = n3935 & n5949 ;
  assign n3942 = n3934 | n3941 ;
  assign n3943 = x50 & n3942 ;
  assign n3944 = x50 | n3942 ;
  assign n5950 = ~n3678 ;
  assign n3945 = n5950 & n3679 ;
  assign n3946 = n68 & n3945 ;
  assign n3947 = n5858 & n3946 ;
  assign n5951 = ~n3946 ;
  assign n3948 = n3684 & n5951 ;
  assign n3949 = n3947 | n3948 ;
  assign n5952 = ~n3949 ;
  assign n3950 = n3944 & n5952 ;
  assign n3951 = n3943 | n3950 ;
  assign n3952 = x51 & n3951 ;
  assign n3953 = x51 | n3951 ;
  assign n5953 = ~n3687 ;
  assign n3954 = n5953 & n3688 ;
  assign n3955 = n68 & n3954 ;
  assign n3956 = n3693 & n3955 ;
  assign n3957 = n3693 | n3955 ;
  assign n5954 = ~n3956 ;
  assign n3958 = n5954 & n3957 ;
  assign n5955 = ~n3958 ;
  assign n3959 = n3953 & n5955 ;
  assign n3960 = n3952 | n3959 ;
  assign n3961 = x52 & n3960 ;
  assign n3962 = x52 | n3960 ;
  assign n5956 = ~n3696 ;
  assign n3963 = n5956 & n3697 ;
  assign n3964 = n68 & n3963 ;
  assign n3965 = n3702 & n3964 ;
  assign n3966 = n3702 | n3964 ;
  assign n5957 = ~n3965 ;
  assign n3967 = n5957 & n3966 ;
  assign n5958 = ~n3967 ;
  assign n3968 = n3962 & n5958 ;
  assign n3969 = n3961 | n3968 ;
  assign n3970 = x53 & n3969 ;
  assign n3971 = x53 | n3969 ;
  assign n5959 = ~n3705 ;
  assign n3972 = n5959 & n3706 ;
  assign n3973 = n68 & n3972 ;
  assign n3974 = n3711 & n3973 ;
  assign n3975 = n3711 | n3973 ;
  assign n5960 = ~n3974 ;
  assign n3976 = n5960 & n3975 ;
  assign n5961 = ~n3976 ;
  assign n3977 = n3971 & n5961 ;
  assign n3978 = n3970 | n3977 ;
  assign n3979 = x54 & n3978 ;
  assign n3980 = x54 | n3978 ;
  assign n5962 = ~n3714 ;
  assign n3981 = n5962 & n3715 ;
  assign n3982 = n68 & n3981 ;
  assign n3983 = n3720 & n3982 ;
  assign n3984 = n3720 | n3982 ;
  assign n5963 = ~n3983 ;
  assign n3985 = n5963 & n3984 ;
  assign n5964 = ~n3985 ;
  assign n3986 = n3980 & n5964 ;
  assign n3987 = n3979 | n3986 ;
  assign n3988 = x55 & n3987 ;
  assign n3989 = x55 | n3987 ;
  assign n5965 = ~n3723 ;
  assign n3990 = n5965 & n3724 ;
  assign n3991 = n68 & n3990 ;
  assign n3992 = n3729 & n3991 ;
  assign n3993 = n3729 | n3991 ;
  assign n5966 = ~n3992 ;
  assign n3994 = n5966 & n3993 ;
  assign n5967 = ~n3994 ;
  assign n3995 = n3989 & n5967 ;
  assign n3996 = n3988 | n3995 ;
  assign n3997 = x56 & n3996 ;
  assign n3998 = x56 | n3996 ;
  assign n5968 = ~n3732 ;
  assign n3999 = n5968 & n3733 ;
  assign n4000 = n68 & n3999 ;
  assign n4001 = n5876 & n4000 ;
  assign n5969 = ~n4000 ;
  assign n4002 = n3738 & n5969 ;
  assign n4003 = n4001 | n4002 ;
  assign n5970 = ~n4003 ;
  assign n4004 = n3998 & n5970 ;
  assign n4005 = n3997 | n4004 ;
  assign n4006 = x57 & n4005 ;
  assign n4007 = x57 | n4005 ;
  assign n5971 = ~n3741 ;
  assign n4008 = n5971 & n3742 ;
  assign n4009 = n68 & n4008 ;
  assign n4010 = n3747 & n4009 ;
  assign n4011 = n3747 | n4009 ;
  assign n5972 = ~n4010 ;
  assign n4012 = n5972 & n4011 ;
  assign n5973 = ~n4012 ;
  assign n4013 = n4007 & n5973 ;
  assign n4014 = n4006 | n4013 ;
  assign n4015 = x58 & n4014 ;
  assign n4016 = x58 | n4014 ;
  assign n5974 = ~n3750 ;
  assign n4017 = n5974 & n3751 ;
  assign n4018 = n68 & n4017 ;
  assign n4019 = n3756 & n4018 ;
  assign n4020 = n3756 | n4018 ;
  assign n5975 = ~n4019 ;
  assign n4021 = n5975 & n4020 ;
  assign n5976 = ~n4021 ;
  assign n4022 = n4016 & n5976 ;
  assign n4023 = n4015 | n4022 ;
  assign n4024 = x59 & n4023 ;
  assign n4025 = x59 | n4023 ;
  assign n5977 = ~n3759 ;
  assign n4026 = n5977 & n3760 ;
  assign n4027 = n68 & n4026 ;
  assign n4028 = n5885 & n4027 ;
  assign n5978 = ~n4027 ;
  assign n4029 = n3765 & n5978 ;
  assign n4030 = n4028 | n4029 ;
  assign n5979 = ~n4030 ;
  assign n4031 = n4025 & n5979 ;
  assign n4032 = n4024 | n4031 ;
  assign n4033 = x60 & n4032 ;
  assign n5980 = ~n3768 ;
  assign n4034 = n5980 & n3769 ;
  assign n4035 = n68 & n4034 ;
  assign n4036 = n3774 & n4035 ;
  assign n4037 = n3774 | n4035 ;
  assign n5981 = ~n4036 ;
  assign n4038 = n5981 & n4037 ;
  assign n4039 = x60 | n4032 ;
  assign n5982 = ~n4038 ;
  assign n4040 = n5982 & n4039 ;
  assign n4041 = n4033 | n4040 ;
  assign n5983 = ~n3781 ;
  assign n4042 = n5983 & n4041 ;
  assign n4043 = x61 | n4042 ;
  assign n5984 = ~n4041 ;
  assign n4044 = n3529 & n5984 ;
  assign n5985 = ~n4044 ;
  assign n4045 = n4043 & n5985 ;
  assign n4046 = n112 | n4045 ;
  assign n67 = ~n4046 ;
  assign n4047 = x32 & n67 ;
  assign n4048 = x2 & n4047 ;
  assign n4050 = x2 | n4047 ;
  assign n5987 = ~n4048 ;
  assign n4051 = n5987 & n4050 ;
  assign n108 = n4597 & x32 ;
  assign n4052 = x33 | n108 ;
  assign n5988 = ~n4051 ;
  assign n4053 = n5988 & n4052 ;
  assign n4054 = n109 | n4053 ;
  assign n4055 = x34 & n4054 ;
  assign n4049 = n5892 & n4047 ;
  assign n5989 = ~n4047 ;
  assign n4056 = x2 & n5989 ;
  assign n4057 = n4049 | n4056 ;
  assign n5990 = ~n4057 ;
  assign n4058 = n4052 & n5990 ;
  assign n4059 = n109 | n4058 ;
  assign n4060 = x34 | n4059 ;
  assign n5991 = ~n107 ;
  assign n4061 = n5991 & n3791 ;
  assign n4062 = n67 & n4061 ;
  assign n4063 = n3790 & n4062 ;
  assign n4064 = n3790 | n4062 ;
  assign n5992 = ~n4063 ;
  assign n4065 = n5992 & n4064 ;
  assign n5993 = ~n4065 ;
  assign n4066 = n4060 & n5993 ;
  assign n4067 = n4055 | n4066 ;
  assign n4068 = x35 | n4067 ;
  assign n4069 = x35 & n4067 ;
  assign n4070 = n3794 | n4046 ;
  assign n5994 = ~n4070 ;
  assign n4071 = n3805 & n5994 ;
  assign n4072 = x34 | n3793 ;
  assign n4073 = n5994 & n4072 ;
  assign n5995 = ~n4073 ;
  assign n4074 = n3804 & n5995 ;
  assign n4075 = n4071 | n4074 ;
  assign n5996 = ~n4069 ;
  assign n4076 = n5996 & n4075 ;
  assign n5997 = ~n4076 ;
  assign n4077 = n4068 & n5997 ;
  assign n4078 = x36 & n4077 ;
  assign n4079 = x36 | n4077 ;
  assign n5998 = ~n3807 ;
  assign n4080 = n5998 & n3808 ;
  assign n4081 = n67 & n4080 ;
  assign n4082 = n3813 & n4081 ;
  assign n4083 = n3813 | n4081 ;
  assign n5999 = ~n4082 ;
  assign n4084 = n5999 & n4083 ;
  assign n6000 = ~n4084 ;
  assign n4085 = n4079 & n6000 ;
  assign n4086 = n4078 | n4085 ;
  assign n4087 = x37 & n4086 ;
  assign n4088 = x37 | n4086 ;
  assign n6001 = ~n3816 ;
  assign n4089 = n6001 & n3817 ;
  assign n4090 = n67 & n4089 ;
  assign n4091 = n3823 & n4090 ;
  assign n4092 = n3823 | n4090 ;
  assign n6002 = ~n4091 ;
  assign n4093 = n6002 & n4092 ;
  assign n6003 = ~n4093 ;
  assign n4094 = n4088 & n6003 ;
  assign n4095 = n4087 | n4094 ;
  assign n4096 = x38 & n4095 ;
  assign n4097 = x38 | n4095 ;
  assign n6004 = ~n3826 ;
  assign n4098 = n6004 & n3827 ;
  assign n4099 = n67 & n4098 ;
  assign n4100 = n3832 & n4099 ;
  assign n4101 = n3832 | n4099 ;
  assign n6005 = ~n4100 ;
  assign n4102 = n6005 & n4101 ;
  assign n6006 = ~n4102 ;
  assign n4103 = n4097 & n6006 ;
  assign n4104 = n4096 | n4103 ;
  assign n4105 = x39 & n4104 ;
  assign n4106 = x39 | n4104 ;
  assign n6007 = ~n3835 ;
  assign n4107 = n6007 & n3836 ;
  assign n4108 = n67 & n4107 ;
  assign n4109 = n3841 & n4108 ;
  assign n4110 = n3841 | n4108 ;
  assign n6008 = ~n4109 ;
  assign n4111 = n6008 & n4110 ;
  assign n6009 = ~n4111 ;
  assign n4112 = n4106 & n6009 ;
  assign n4113 = n4105 | n4112 ;
  assign n4114 = x40 & n4113 ;
  assign n4115 = x40 | n4113 ;
  assign n6010 = ~n3844 ;
  assign n4116 = n6010 & n3845 ;
  assign n4117 = n67 & n4116 ;
  assign n4118 = n5919 & n4117 ;
  assign n6011 = ~n4117 ;
  assign n4119 = n3850 & n6011 ;
  assign n4120 = n4118 | n4119 ;
  assign n6012 = ~n4120 ;
  assign n4121 = n4115 & n6012 ;
  assign n4122 = n4114 | n4121 ;
  assign n4123 = x41 & n4122 ;
  assign n4124 = x41 | n4122 ;
  assign n6013 = ~n3853 ;
  assign n4125 = n6013 & n3854 ;
  assign n4126 = n67 & n4125 ;
  assign n4127 = n5922 & n4126 ;
  assign n6014 = ~n4126 ;
  assign n4128 = n3859 & n6014 ;
  assign n4129 = n4127 | n4128 ;
  assign n6015 = ~n4129 ;
  assign n4130 = n4124 & n6015 ;
  assign n4131 = n4123 | n4130 ;
  assign n4132 = x42 & n4131 ;
  assign n4133 = x42 | n4131 ;
  assign n6016 = ~n3862 ;
  assign n4134 = n6016 & n3863 ;
  assign n4135 = n67 & n4134 ;
  assign n4136 = n3868 & n4135 ;
  assign n4137 = n3868 | n4135 ;
  assign n6017 = ~n4136 ;
  assign n4138 = n6017 & n4137 ;
  assign n6018 = ~n4138 ;
  assign n4139 = n4133 & n6018 ;
  assign n4140 = n4132 | n4139 ;
  assign n4141 = x43 & n4140 ;
  assign n4142 = x43 | n4140 ;
  assign n6019 = ~n3871 ;
  assign n4143 = n6019 & n3872 ;
  assign n4144 = n67 & n4143 ;
  assign n4145 = n3877 & n4144 ;
  assign n4146 = n3877 | n4144 ;
  assign n6020 = ~n4145 ;
  assign n4147 = n6020 & n4146 ;
  assign n6021 = ~n4147 ;
  assign n4148 = n4142 & n6021 ;
  assign n4149 = n4141 | n4148 ;
  assign n4150 = x44 & n4149 ;
  assign n4151 = x44 | n4149 ;
  assign n6022 = ~n3880 ;
  assign n4152 = n6022 & n3881 ;
  assign n4153 = n67 & n4152 ;
  assign n4154 = n3886 & n4153 ;
  assign n4155 = n3886 | n4153 ;
  assign n6023 = ~n4154 ;
  assign n4156 = n6023 & n4155 ;
  assign n6024 = ~n4156 ;
  assign n4157 = n4151 & n6024 ;
  assign n4158 = n4150 | n4157 ;
  assign n4159 = x45 & n4158 ;
  assign n4160 = x45 | n4158 ;
  assign n6025 = ~n3889 ;
  assign n4161 = n6025 & n3890 ;
  assign n4162 = n67 & n4161 ;
  assign n4163 = n5934 & n4162 ;
  assign n6026 = ~n4162 ;
  assign n4164 = n3895 & n6026 ;
  assign n4165 = n4163 | n4164 ;
  assign n6027 = ~n4165 ;
  assign n4166 = n4160 & n6027 ;
  assign n4167 = n4159 | n4166 ;
  assign n4168 = x46 & n4167 ;
  assign n6028 = ~n3898 ;
  assign n4169 = n6028 & n3904 ;
  assign n4170 = n67 & n4169 ;
  assign n4171 = n3903 & n4170 ;
  assign n4172 = n3903 | n4170 ;
  assign n6029 = ~n4171 ;
  assign n4173 = n6029 & n4172 ;
  assign n4174 = x46 | n4167 ;
  assign n6030 = ~n4173 ;
  assign n4175 = n6030 & n4174 ;
  assign n4176 = n4168 | n4175 ;
  assign n4177 = x47 & n4176 ;
  assign n6031 = ~n3907 ;
  assign n4178 = n6031 & n3908 ;
  assign n4179 = n67 & n4178 ;
  assign n4180 = n3913 & n4179 ;
  assign n4181 = n3913 | n4179 ;
  assign n6032 = ~n4180 ;
  assign n4182 = n6032 & n4181 ;
  assign n4183 = x47 | n4176 ;
  assign n6033 = ~n4182 ;
  assign n4184 = n6033 & n4183 ;
  assign n4185 = n4177 | n4184 ;
  assign n4186 = x48 & n4185 ;
  assign n4187 = x48 | n4185 ;
  assign n6034 = ~n3916 ;
  assign n4188 = n6034 & n3917 ;
  assign n4189 = n67 & n4188 ;
  assign n4190 = n5943 & n4189 ;
  assign n6035 = ~n4189 ;
  assign n4191 = n3922 & n6035 ;
  assign n4192 = n4190 | n4191 ;
  assign n6036 = ~n4192 ;
  assign n4193 = n4187 & n6036 ;
  assign n4194 = n4186 | n4193 ;
  assign n4195 = x49 & n4194 ;
  assign n4196 = x49 | n4194 ;
  assign n6037 = ~n3925 ;
  assign n4197 = n6037 & n3926 ;
  assign n4198 = n67 & n4197 ;
  assign n4199 = n3931 & n4198 ;
  assign n4200 = n3931 | n4198 ;
  assign n6038 = ~n4199 ;
  assign n4201 = n6038 & n4200 ;
  assign n6039 = ~n4201 ;
  assign n4202 = n4196 & n6039 ;
  assign n4203 = n4195 | n4202 ;
  assign n4204 = x50 & n4203 ;
  assign n4205 = x50 | n4203 ;
  assign n6040 = ~n3934 ;
  assign n4206 = n6040 & n3935 ;
  assign n4207 = n67 & n4206 ;
  assign n4208 = n3940 & n4207 ;
  assign n4209 = n3940 | n4207 ;
  assign n6041 = ~n4208 ;
  assign n4210 = n6041 & n4209 ;
  assign n6042 = ~n4210 ;
  assign n4211 = n4205 & n6042 ;
  assign n4212 = n4204 | n4211 ;
  assign n4213 = x51 & n4212 ;
  assign n4214 = x51 | n4212 ;
  assign n6043 = ~n3943 ;
  assign n4215 = n6043 & n3944 ;
  assign n4216 = n67 & n4215 ;
  assign n4217 = n3949 & n4216 ;
  assign n4218 = n3949 | n4216 ;
  assign n6044 = ~n4217 ;
  assign n4219 = n6044 & n4218 ;
  assign n6045 = ~n4219 ;
  assign n4220 = n4214 & n6045 ;
  assign n4221 = n4213 | n4220 ;
  assign n4222 = x52 & n4221 ;
  assign n4223 = x52 | n4221 ;
  assign n6046 = ~n3952 ;
  assign n4224 = n6046 & n3953 ;
  assign n4225 = n67 & n4224 ;
  assign n4226 = n3958 & n4225 ;
  assign n4227 = n3958 | n4225 ;
  assign n6047 = ~n4226 ;
  assign n4228 = n6047 & n4227 ;
  assign n6048 = ~n4228 ;
  assign n4229 = n4223 & n6048 ;
  assign n4230 = n4222 | n4229 ;
  assign n4231 = x53 & n4230 ;
  assign n4232 = x53 | n4230 ;
  assign n6049 = ~n3961 ;
  assign n4233 = n6049 & n3962 ;
  assign n4234 = n67 & n4233 ;
  assign n4235 = n3967 & n4234 ;
  assign n4236 = n3967 | n4234 ;
  assign n6050 = ~n4235 ;
  assign n4237 = n6050 & n4236 ;
  assign n6051 = ~n4237 ;
  assign n4238 = n4232 & n6051 ;
  assign n4239 = n4231 | n4238 ;
  assign n4240 = x54 & n4239 ;
  assign n4241 = x54 | n4239 ;
  assign n6052 = ~n3970 ;
  assign n4242 = n6052 & n3971 ;
  assign n4243 = n67 & n4242 ;
  assign n4244 = n3976 & n4243 ;
  assign n4245 = n3976 | n4243 ;
  assign n6053 = ~n4244 ;
  assign n4246 = n6053 & n4245 ;
  assign n6054 = ~n4246 ;
  assign n4247 = n4241 & n6054 ;
  assign n4248 = n4240 | n4247 ;
  assign n4249 = x55 & n4248 ;
  assign n4250 = x55 | n4248 ;
  assign n6055 = ~n3979 ;
  assign n4251 = n6055 & n3980 ;
  assign n4252 = n67 & n4251 ;
  assign n4253 = n3985 & n4252 ;
  assign n4254 = n3985 | n4252 ;
  assign n6056 = ~n4253 ;
  assign n4255 = n6056 & n4254 ;
  assign n6057 = ~n4255 ;
  assign n4256 = n4250 & n6057 ;
  assign n4257 = n4249 | n4256 ;
  assign n4258 = x56 & n4257 ;
  assign n4259 = x56 | n4257 ;
  assign n6058 = ~n3988 ;
  assign n4260 = n6058 & n3989 ;
  assign n4261 = n67 & n4260 ;
  assign n4262 = n3994 & n4261 ;
  assign n4263 = n3994 | n4261 ;
  assign n6059 = ~n4262 ;
  assign n4264 = n6059 & n4263 ;
  assign n6060 = ~n4264 ;
  assign n4265 = n4259 & n6060 ;
  assign n4266 = n4258 | n4265 ;
  assign n4267 = x57 & n4266 ;
  assign n4268 = x57 | n4266 ;
  assign n6061 = ~n3997 ;
  assign n4269 = n6061 & n3998 ;
  assign n4270 = n67 & n4269 ;
  assign n4271 = n5970 & n4270 ;
  assign n6062 = ~n4270 ;
  assign n4272 = n4003 & n6062 ;
  assign n4273 = n4271 | n4272 ;
  assign n6063 = ~n4273 ;
  assign n4274 = n4268 & n6063 ;
  assign n4275 = n4267 | n4274 ;
  assign n4276 = x58 & n4275 ;
  assign n4277 = x58 | n4275 ;
  assign n6064 = ~n4006 ;
  assign n4278 = n6064 & n4007 ;
  assign n4279 = n67 & n4278 ;
  assign n4280 = n4012 & n4279 ;
  assign n4281 = n4012 | n4279 ;
  assign n6065 = ~n4280 ;
  assign n4282 = n6065 & n4281 ;
  assign n6066 = ~n4282 ;
  assign n4283 = n4277 & n6066 ;
  assign n4284 = n4276 | n4283 ;
  assign n4285 = x59 & n4284 ;
  assign n4286 = x59 | n4284 ;
  assign n6067 = ~n4015 ;
  assign n4287 = n6067 & n4016 ;
  assign n4288 = n67 & n4287 ;
  assign n4289 = n5976 & n4288 ;
  assign n6068 = ~n4288 ;
  assign n4290 = n4021 & n6068 ;
  assign n4291 = n4289 | n4290 ;
  assign n6069 = ~n4291 ;
  assign n4292 = n4286 & n6069 ;
  assign n4293 = n4285 | n4292 ;
  assign n4294 = x60 & n4293 ;
  assign n4295 = x60 | n4293 ;
  assign n6070 = ~n4024 ;
  assign n4296 = n6070 & n4025 ;
  assign n4297 = n67 & n4296 ;
  assign n4298 = n4030 & n4297 ;
  assign n4299 = n4030 | n4297 ;
  assign n6071 = ~n4298 ;
  assign n4300 = n6071 & n4299 ;
  assign n6072 = ~n4300 ;
  assign n4301 = n4295 & n6072 ;
  assign n4302 = n4294 | n4301 ;
  assign n4303 = x61 & n4302 ;
  assign n6073 = ~n4033 ;
  assign n4304 = n6073 & n4039 ;
  assign n4305 = n67 & n4304 ;
  assign n4306 = n4038 & n4305 ;
  assign n4307 = n4038 | n4305 ;
  assign n6074 = ~n4306 ;
  assign n4308 = n6074 & n4307 ;
  assign n4309 = x61 | n4302 ;
  assign n6075 = ~n4308 ;
  assign n4310 = n6075 & n4309 ;
  assign n4311 = n4303 | n4310 ;
  assign n4312 = x62 & n4311 ;
  assign n4313 = x62 | n4311 ;
  assign n6076 = ~n4312 ;
  assign n4322 = n6076 & n4313 ;
  assign n4314 = x61 & n4041 ;
  assign n4315 = x61 | n4041 ;
  assign n6077 = ~n112 ;
  assign n4316 = n6077 & n4315 ;
  assign n6078 = ~n4314 ;
  assign n4317 = n6078 & n4316 ;
  assign n6079 = ~n4317 ;
  assign n4318 = n3781 & n6079 ;
  assign n6080 = ~x63 ;
  assign n4323 = n6080 & n4318 ;
  assign n6081 = ~n4322 ;
  assign n4594 = n6081 & n4323 ;
  assign n6082 = ~n4318 ;
  assign n4319 = n4313 & n6082 ;
  assign n4320 = x63 | n4312 ;
  assign n4321 = n4319 | n4320 ;
  assign n6083 = ~n4276 ;
  assign n4555 = n6083 & n4277 ;
  assign n66 = ~n4321 ;
  assign n4556 = n66 & n4555 ;
  assign n4557 = n4282 & n4556 ;
  assign n4558 = n4282 | n4556 ;
  assign n6085 = ~n4557 ;
  assign n4559 = n6085 & n4558 ;
  assign n6086 = ~x59 ;
  assign n4560 = n6086 & n4559 ;
  assign n6087 = ~n4285 ;
  assign n4564 = n6087 & n4286 ;
  assign n4565 = n66 & n4564 ;
  assign n4566 = n6069 & n4565 ;
  assign n6088 = ~n4565 ;
  assign n4567 = n4291 & n6088 ;
  assign n4568 = n4566 | n4567 ;
  assign n4570 = n5893 & n4568 ;
  assign n4571 = n4560 | n4570 ;
  assign n6089 = ~n4240 ;
  assign n4520 = n6089 & n4241 ;
  assign n4521 = n66 & n4520 ;
  assign n4522 = n4246 & n4521 ;
  assign n4523 = n4246 | n4521 ;
  assign n6090 = ~n4522 ;
  assign n4524 = n6090 & n4523 ;
  assign n6091 = ~x55 ;
  assign n4525 = n6091 & n4524 ;
  assign n6092 = ~n4249 ;
  assign n4528 = n6092 & n4250 ;
  assign n4529 = n66 & n4528 ;
  assign n4530 = n6057 & n4529 ;
  assign n6093 = ~n4529 ;
  assign n4531 = n4255 & n6093 ;
  assign n4532 = n4530 | n4531 ;
  assign n6094 = ~x56 ;
  assign n4534 = n6094 & n4532 ;
  assign n4535 = n4525 | n4534 ;
  assign n6095 = ~n4204 ;
  assign n4484 = n6095 & n4205 ;
  assign n4485 = n66 & n4484 ;
  assign n4486 = n4210 & n4485 ;
  assign n4487 = n4210 | n4485 ;
  assign n6096 = ~n4486 ;
  assign n4488 = n6096 & n4487 ;
  assign n6097 = ~x51 ;
  assign n4489 = n6097 & n4488 ;
  assign n6098 = ~n4213 ;
  assign n4492 = n6098 & n4214 ;
  assign n4493 = n66 & n4492 ;
  assign n4494 = n4219 & n4493 ;
  assign n4495 = n4219 | n4493 ;
  assign n6099 = ~n4494 ;
  assign n4496 = n6099 & n4495 ;
  assign n6100 = ~x52 ;
  assign n4497 = n6100 & n4496 ;
  assign n4498 = n4489 | n4497 ;
  assign n6101 = ~n4168 ;
  assign n4324 = n6101 & n4174 ;
  assign n4325 = n66 & n4324 ;
  assign n4326 = n4173 & n4325 ;
  assign n4327 = n4173 | n4325 ;
  assign n6102 = ~n4326 ;
  assign n4328 = n6102 & n4327 ;
  assign n6103 = ~x47 ;
  assign n4329 = n6103 & n4328 ;
  assign n6104 = ~n4177 ;
  assign n4456 = n6104 & n4183 ;
  assign n4457 = n66 & n4456 ;
  assign n4458 = n6033 & n4457 ;
  assign n6105 = ~n4457 ;
  assign n4459 = n4182 & n6105 ;
  assign n4460 = n4458 | n4459 ;
  assign n6106 = ~x48 ;
  assign n4462 = n6106 & n4460 ;
  assign n4463 = n4329 | n4462 ;
  assign n6107 = ~n4328 ;
  assign n4330 = x47 & n6107 ;
  assign n6108 = ~n4159 ;
  assign n4331 = n6108 & n4160 ;
  assign n4332 = n66 & n4331 ;
  assign n4333 = n6027 & n4332 ;
  assign n6109 = ~n4332 ;
  assign n4334 = n4165 & n6109 ;
  assign n4335 = n4333 | n4334 ;
  assign n6110 = ~x46 ;
  assign n4337 = n6110 & n4335 ;
  assign n6111 = ~n4141 ;
  assign n4435 = n6111 & n4142 ;
  assign n4436 = n66 & n4435 ;
  assign n4437 = n4147 & n4436 ;
  assign n4438 = n4147 | n4436 ;
  assign n6112 = ~n4437 ;
  assign n4439 = n6112 & n4438 ;
  assign n6113 = ~x44 ;
  assign n4440 = n6113 & n4439 ;
  assign n6114 = ~n4150 ;
  assign n4443 = n6114 & n4151 ;
  assign n4444 = n66 & n4443 ;
  assign n4445 = n4156 & n4444 ;
  assign n4446 = n4156 | n4444 ;
  assign n6115 = ~n4445 ;
  assign n4447 = n6115 & n4446 ;
  assign n6116 = ~x45 ;
  assign n4448 = n6116 & n4447 ;
  assign n4449 = n4440 | n4448 ;
  assign n6117 = ~n4105 ;
  assign n4399 = n6117 & n4106 ;
  assign n4400 = n66 & n4399 ;
  assign n4401 = n4111 & n4400 ;
  assign n4402 = n4111 | n4400 ;
  assign n6118 = ~n4401 ;
  assign n4403 = n6118 & n4402 ;
  assign n6119 = ~x40 ;
  assign n4404 = n6119 & n4403 ;
  assign n6120 = ~n4114 ;
  assign n4407 = n6120 & n4115 ;
  assign n4408 = n66 & n4407 ;
  assign n4409 = n6012 & n4408 ;
  assign n6121 = ~n4408 ;
  assign n4410 = n4120 & n6121 ;
  assign n4411 = n4409 | n4410 ;
  assign n6122 = ~x41 ;
  assign n4413 = n6122 & n4411 ;
  assign n4414 = n4404 | n4413 ;
  assign n6123 = ~n4078 ;
  assign n4374 = n6123 & n4079 ;
  assign n4375 = n66 & n4374 ;
  assign n4376 = n4084 & n4375 ;
  assign n4377 = n4084 | n4375 ;
  assign n6124 = ~n4376 ;
  assign n4378 = n6124 & n4377 ;
  assign n4338 = n4068 & n5996 ;
  assign n4339 = n66 & n4338 ;
  assign n6125 = ~n4075 ;
  assign n4340 = n6125 & n4339 ;
  assign n6126 = ~n4339 ;
  assign n4341 = n4075 & n6126 ;
  assign n4342 = n4340 | n4341 ;
  assign n6127 = ~x36 ;
  assign n4343 = n6127 & n4342 ;
  assign n6128 = ~n4342 ;
  assign n4344 = x36 & n6128 ;
  assign n4345 = x34 | n4054 ;
  assign n4346 = n4055 | n4321 ;
  assign n6129 = ~n4346 ;
  assign n4347 = n4345 & n6129 ;
  assign n6130 = ~n4347 ;
  assign n4348 = n4065 & n6130 ;
  assign n4349 = n4066 & n6129 ;
  assign n4350 = n4348 | n4349 ;
  assign n4351 = n5416 & n4350 ;
  assign n6131 = ~n4350 ;
  assign n4352 = x35 & n6131 ;
  assign n6132 = ~n109 ;
  assign n4353 = n6132 & n4052 ;
  assign n4354 = n66 & n4353 ;
  assign n4355 = n4051 & n4354 ;
  assign n4356 = n4051 | n4354 ;
  assign n6133 = ~n4355 ;
  assign n4357 = n6133 & n4356 ;
  assign n6134 = ~x34 ;
  assign n4358 = n6134 & n4357 ;
  assign n6135 = ~n4357 ;
  assign n4359 = x34 & n6135 ;
  assign n6136 = ~x0 ;
  assign n111 = n6136 & n4602 ;
  assign n4360 = x32 & n66 ;
  assign n6137 = ~n4360 ;
  assign n4362 = x1 & n6137 ;
  assign n4361 = n4597 & n4360 ;
  assign n110 = n6136 & x32 ;
  assign n4363 = x33 | n110 ;
  assign n6138 = ~n4361 ;
  assign n4364 = n6138 & n4363 ;
  assign n6139 = ~n4362 ;
  assign n4365 = n6139 & n4364 ;
  assign n4366 = n111 | n4365 ;
  assign n4367 = n4359 | n4366 ;
  assign n6140 = ~n4358 ;
  assign n4368 = n6140 & n4367 ;
  assign n4369 = n4352 | n4368 ;
  assign n6141 = ~n4351 ;
  assign n4370 = n6141 & n4369 ;
  assign n4371 = n4344 | n4370 ;
  assign n6142 = ~n4343 ;
  assign n4372 = n6142 & n4371 ;
  assign n4379 = x37 | n4372 ;
  assign n6143 = ~n4378 ;
  assign n4380 = n6143 & n4379 ;
  assign n4373 = x37 & n4372 ;
  assign n6144 = ~n4087 ;
  assign n4381 = n6144 & n4088 ;
  assign n4382 = n66 & n4381 ;
  assign n6145 = ~n4382 ;
  assign n4383 = n4093 & n6145 ;
  assign n4384 = n6003 & n4382 ;
  assign n4385 = n4383 | n4384 ;
  assign n6146 = ~n4385 ;
  assign n4386 = x38 & n6146 ;
  assign n4387 = n4373 | n4386 ;
  assign n4388 = n4380 | n4387 ;
  assign n6147 = ~x38 ;
  assign n4395 = n6147 & n4385 ;
  assign n6148 = ~n4096 ;
  assign n4389 = n6148 & n4097 ;
  assign n4390 = n66 & n4389 ;
  assign n4391 = n4102 & n4390 ;
  assign n4392 = n4102 | n4390 ;
  assign n6149 = ~n4391 ;
  assign n4393 = n6149 & n4392 ;
  assign n6150 = ~x39 ;
  assign n4396 = n6150 & n4393 ;
  assign n4397 = n4395 | n4396 ;
  assign n6151 = ~n4397 ;
  assign n4398 = n4388 & n6151 ;
  assign n6152 = ~n4393 ;
  assign n4394 = x39 & n6152 ;
  assign n6153 = ~n4403 ;
  assign n4405 = x40 & n6153 ;
  assign n4406 = n4394 | n4405 ;
  assign n4415 = n4398 | n4406 ;
  assign n6154 = ~n4414 ;
  assign n4416 = n6154 & n4415 ;
  assign n6155 = ~n4411 ;
  assign n4412 = x41 & n6155 ;
  assign n6156 = ~n4123 ;
  assign n4417 = n6156 & n4124 ;
  assign n4418 = n66 & n4417 ;
  assign n4419 = n6015 & n4418 ;
  assign n6157 = ~n4418 ;
  assign n4420 = n4129 & n6157 ;
  assign n4421 = n4419 | n4420 ;
  assign n6158 = ~n4421 ;
  assign n4422 = x42 & n6158 ;
  assign n4423 = n4412 | n4422 ;
  assign n4424 = n4416 | n4423 ;
  assign n6159 = ~x42 ;
  assign n4431 = n6159 & n4421 ;
  assign n6160 = ~n4132 ;
  assign n4425 = n6160 & n4133 ;
  assign n4426 = n66 & n4425 ;
  assign n4427 = n6018 & n4426 ;
  assign n6161 = ~n4426 ;
  assign n4428 = n4138 & n6161 ;
  assign n4429 = n4427 | n4428 ;
  assign n6162 = ~x43 ;
  assign n4432 = n6162 & n4429 ;
  assign n4433 = n4431 | n4432 ;
  assign n6163 = ~n4433 ;
  assign n4434 = n4424 & n6163 ;
  assign n6164 = ~n4429 ;
  assign n4430 = x43 & n6164 ;
  assign n6165 = ~n4439 ;
  assign n4441 = x44 & n6165 ;
  assign n4442 = n4430 | n4441 ;
  assign n4450 = n4434 | n4442 ;
  assign n6166 = ~n4449 ;
  assign n4451 = n6166 & n4450 ;
  assign n6167 = ~n4335 ;
  assign n4336 = x46 & n6167 ;
  assign n6168 = ~n4447 ;
  assign n4452 = x45 & n6168 ;
  assign n4453 = n4336 | n4452 ;
  assign n4454 = n4451 | n4453 ;
  assign n6169 = ~n4337 ;
  assign n4455 = n6169 & n4454 ;
  assign n4464 = n4330 | n4455 ;
  assign n6170 = ~n4463 ;
  assign n4465 = n6170 & n4464 ;
  assign n6171 = ~n4460 ;
  assign n4461 = x48 & n6171 ;
  assign n6172 = ~n4186 ;
  assign n4466 = n6172 & n4187 ;
  assign n4467 = n66 & n4466 ;
  assign n4468 = n6036 & n4467 ;
  assign n6173 = ~n4467 ;
  assign n4469 = n4192 & n6173 ;
  assign n4470 = n4468 | n4469 ;
  assign n6174 = ~n4470 ;
  assign n4471 = x49 & n6174 ;
  assign n4472 = n4461 | n4471 ;
  assign n4473 = n4465 | n4472 ;
  assign n6175 = ~x49 ;
  assign n4480 = n6175 & n4470 ;
  assign n6176 = ~n4195 ;
  assign n4474 = n6176 & n4196 ;
  assign n4475 = n66 & n4474 ;
  assign n4476 = n6039 & n4475 ;
  assign n6177 = ~n4475 ;
  assign n4477 = n4201 & n6177 ;
  assign n4478 = n4476 | n4477 ;
  assign n6178 = ~x50 ;
  assign n4481 = n6178 & n4478 ;
  assign n4482 = n4480 | n4481 ;
  assign n6179 = ~n4482 ;
  assign n4483 = n4473 & n6179 ;
  assign n6180 = ~n4478 ;
  assign n4479 = x50 & n6180 ;
  assign n6181 = ~n4488 ;
  assign n4490 = x51 & n6181 ;
  assign n4491 = n4479 | n4490 ;
  assign n4499 = n4483 | n4491 ;
  assign n6182 = ~n4498 ;
  assign n4500 = n6182 & n4499 ;
  assign n6183 = ~n4496 ;
  assign n4501 = x52 & n6183 ;
  assign n6184 = ~n4222 ;
  assign n4502 = n6184 & n4223 ;
  assign n4503 = n66 & n4502 ;
  assign n6185 = ~n4503 ;
  assign n4504 = n4228 & n6185 ;
  assign n4505 = n6048 & n4503 ;
  assign n4506 = n4504 | n4505 ;
  assign n6186 = ~n4506 ;
  assign n4507 = x53 & n6186 ;
  assign n4508 = n4501 | n4507 ;
  assign n4509 = n4500 | n4508 ;
  assign n6187 = ~x53 ;
  assign n4516 = n6187 & n4506 ;
  assign n6188 = ~n4231 ;
  assign n4510 = n6188 & n4232 ;
  assign n4511 = n66 & n4510 ;
  assign n4512 = n6051 & n4511 ;
  assign n6189 = ~n4511 ;
  assign n4513 = n4237 & n6189 ;
  assign n4514 = n4512 | n4513 ;
  assign n6190 = ~x54 ;
  assign n4517 = n6190 & n4514 ;
  assign n4518 = n4516 | n4517 ;
  assign n6191 = ~n4518 ;
  assign n4519 = n4509 & n6191 ;
  assign n6192 = ~n4514 ;
  assign n4515 = x54 & n6192 ;
  assign n6193 = ~n4524 ;
  assign n4526 = x55 & n6193 ;
  assign n4527 = n4515 | n4526 ;
  assign n4536 = n4519 | n4527 ;
  assign n6194 = ~n4535 ;
  assign n4537 = n6194 & n4536 ;
  assign n6195 = ~n4532 ;
  assign n4533 = x56 & n6195 ;
  assign n6196 = ~n4258 ;
  assign n4538 = n6196 & n4259 ;
  assign n4539 = n66 & n4538 ;
  assign n6197 = ~n4539 ;
  assign n4540 = n4264 & n6197 ;
  assign n4541 = n6060 & n4539 ;
  assign n4542 = n4540 | n4541 ;
  assign n6198 = ~n4542 ;
  assign n4543 = x57 & n6198 ;
  assign n4544 = n4533 | n4543 ;
  assign n4545 = n4537 | n4544 ;
  assign n6199 = ~n4267 ;
  assign n4546 = n6199 & n4268 ;
  assign n4547 = n66 & n4546 ;
  assign n4548 = n4273 & n4547 ;
  assign n4549 = n4273 | n4547 ;
  assign n6200 = ~n4548 ;
  assign n4550 = n6200 & n4549 ;
  assign n6201 = ~x58 ;
  assign n4551 = n6201 & n4550 ;
  assign n6202 = ~x57 ;
  assign n4552 = n6202 & n4542 ;
  assign n4553 = n4551 | n4552 ;
  assign n6203 = ~n4553 ;
  assign n4554 = n4545 & n6203 ;
  assign n6204 = ~n4550 ;
  assign n4561 = x58 & n6204 ;
  assign n6205 = ~n4559 ;
  assign n4562 = x59 & n6205 ;
  assign n4563 = n4561 | n4562 ;
  assign n4572 = n4554 | n4563 ;
  assign n6206 = ~n4571 ;
  assign n4573 = n6206 & n4572 ;
  assign n6207 = ~n4568 ;
  assign n4569 = x60 & n6207 ;
  assign n6208 = ~n4294 ;
  assign n4574 = n6208 & n4295 ;
  assign n4575 = n66 & n4574 ;
  assign n6209 = ~n4575 ;
  assign n4576 = n4300 & n6209 ;
  assign n4577 = n6072 & n4575 ;
  assign n4578 = n4576 | n4577 ;
  assign n6210 = ~n4578 ;
  assign n4579 = x61 & n6210 ;
  assign n4580 = n4569 | n4579 ;
  assign n4581 = n4573 | n4580 ;
  assign n6211 = ~n4303 ;
  assign n4582 = n6211 & n4309 ;
  assign n4583 = n66 & n4582 ;
  assign n4584 = n4308 & n4583 ;
  assign n4585 = n4308 | n4583 ;
  assign n6212 = ~n4584 ;
  assign n4586 = n6212 & n4585 ;
  assign n6213 = ~x62 ;
  assign n4587 = n6213 & n4586 ;
  assign n6214 = ~x61 ;
  assign n4588 = n6214 & n4578 ;
  assign n4589 = n4587 | n4588 ;
  assign n6215 = ~n4589 ;
  assign n4590 = n4581 & n6215 ;
  assign n4591 = x63 & n5983 ;
  assign n6216 = ~n4586 ;
  assign n4592 = x62 & n6216 ;
  assign n4593 = n4591 | n4592 ;
  assign n4595 = n4590 | n4593 ;
  assign n6217 = ~n4594 ;
  assign n4596 = n6217 & n4595 ;
  assign n65 = ~n4596 ;
  assign y0 = n65 ;
  assign y1 = n66 ;
  assign y2 = n67 ;
  assign y3 = n68 ;
  assign y4 = n69 ;
  assign y5 = n70 ;
  assign y6 = n71 ;
  assign y7 = n72 ;
  assign y8 = n73 ;
  assign y9 = n74 ;
  assign y10 = n75 ;
  assign y11 = n76 ;
  assign y12 = n77 ;
  assign y13 = n78 ;
  assign y14 = n79 ;
  assign y15 = n80 ;
  assign y16 = n81 ;
  assign y17 = n82 ;
  assign y18 = n83 ;
  assign y19 = n84 ;
  assign y20 = n85 ;
  assign y21 = n86 ;
  assign y22 = n87 ;
  assign y23 = n88 ;
  assign y24 = n89 ;
  assign y25 = n90 ;
  assign y26 = n91 ;
  assign y27 = n92 ;
  assign y28 = n93 ;
  assign y29 = n94 ;
  assign y30 = n95 ;
  assign y31 = n96 ;
endmodule
