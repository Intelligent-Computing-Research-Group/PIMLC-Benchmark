module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 ;
  assign n17 = x0 & x8 ;
  assign n42 = x1 & x9 ;
  assign n57 = n17 & n42 ;
  assign n45 = x0 & x9 ;
  assign n46 = x1 & x8 ;
  assign n78 = n45 | n46 ;
  assign n222 = ~n57 ;
  assign n18 = n222 & n78 ;
  assign n75 = x0 & x10 ;
  assign n77 = x2 & x8 ;
  assign n58 = n75 | n77 ;
  assign n79 = n75 & n77 ;
  assign n223 = ~n17 ;
  assign n59 = n223 & n42 ;
  assign n60 = n79 | n59 ;
  assign n61 = n58 & n60 ;
  assign n76 = n58 | n59 ;
  assign n224 = ~n61 ;
  assign n19 = n224 & n76 ;
  assign n41 = x1 & x10 ;
  assign n62 = n57 | n61 ;
  assign n63 = n41 | n62 ;
  assign n64 = n41 & n62 ;
  assign n43 = x2 & x9 ;
  assign n65 = n17 & n43 ;
  assign n225 = ~n65 ;
  assign n66 = n64 & n225 ;
  assign n226 = ~n66 ;
  assign n67 = n63 & n226 ;
  assign n214 = x3 & x8 ;
  assign n215 = x0 & x11 ;
  assign n44 = n214 & n215 ;
  assign n68 = n214 | n215 ;
  assign n227 = ~n44 ;
  assign n69 = n227 & n68 ;
  assign n228 = ~n43 ;
  assign n70 = n228 & n69 ;
  assign n229 = ~n69 ;
  assign n71 = n43 & n229 ;
  assign n72 = n70 | n71 ;
  assign n73 = n67 | n72 ;
  assign n74 = n67 & n72 ;
  assign n230 = ~n74 ;
  assign n20 = n73 & n230 ;
  assign n25 = x4 & x8 ;
  assign n217 = x1 & x11 ;
  assign n221 = x3 & x9 ;
  assign n47 = n217 & n221 ;
  assign n83 = n217 | n221 ;
  assign n231 = ~n47 ;
  assign n84 = n231 & n83 ;
  assign n85 = n25 & n84 ;
  assign n86 = n25 | n84 ;
  assign n232 = ~n85 ;
  assign n87 = n232 & n86 ;
  assign n233 = ~n70 ;
  assign n88 = n68 & n233 ;
  assign n89 = n87 & n88 ;
  assign n90 = n87 | n88 ;
  assign n234 = ~n89 ;
  assign n91 = n234 & n90 ;
  assign n26 = x2 & x10 ;
  assign n27 = x0 & x12 ;
  assign n92 = n26 | n27 ;
  assign n48 = x2 & x12 ;
  assign n95 = n75 & n48 ;
  assign n235 = ~n95 ;
  assign n97 = n92 & n235 ;
  assign n98 = n91 & n97 ;
  assign n99 = n91 | n97 ;
  assign n236 = ~n98 ;
  assign n100 = n236 & n99 ;
  assign n80 = n64 | n74 ;
  assign n81 = n64 & n71 ;
  assign n82 = n67 & n81 ;
  assign n237 = ~n82 ;
  assign n218 = n80 & n237 ;
  assign n219 = n100 & n218 ;
  assign n220 = n100 | n218 ;
  assign n238 = ~n219 ;
  assign n21 = n238 & n220 ;
  assign n101 = n82 | n100 ;
  assign n102 = n80 & n101 ;
  assign n49 = x1 & x12 ;
  assign n28 = x3 & x10 ;
  assign n29 = x0 & x13 ;
  assign n50 = n28 & n29 ;
  assign n103 = n28 | n29 ;
  assign n239 = ~n50 ;
  assign n104 = n239 & n103 ;
  assign n240 = ~n49 ;
  assign n105 = n240 & n104 ;
  assign n241 = ~n104 ;
  assign n106 = n49 & n241 ;
  assign n107 = n105 | n106 ;
  assign n32 = x2 & x11 ;
  assign n30 = x5 & x8 ;
  assign n31 = x4 & x9 ;
  assign n51 = n30 & n31 ;
  assign n108 = n30 | n31 ;
  assign n242 = ~n51 ;
  assign n109 = n242 & n108 ;
  assign n110 = n32 & n109 ;
  assign n111 = n32 | n109 ;
  assign n243 = ~n110 ;
  assign n112 = n243 & n111 ;
  assign n244 = ~n25 ;
  assign n113 = n244 & n84 ;
  assign n245 = ~n113 ;
  assign n114 = n83 & n245 ;
  assign n115 = n112 & n114 ;
  assign n116 = n112 | n114 ;
  assign n246 = ~n115 ;
  assign n117 = n246 & n116 ;
  assign n247 = ~n107 ;
  assign n118 = n247 & n117 ;
  assign n248 = ~n117 ;
  assign n119 = n107 & n248 ;
  assign n120 = n118 | n119 ;
  assign n93 = n91 & n92 ;
  assign n96 = n89 & n95 ;
  assign n121 = n89 | n95 ;
  assign n249 = ~n96 ;
  assign n122 = n249 & n121 ;
  assign n123 = n93 | n122 ;
  assign n124 = n120 | n123 ;
  assign n125 = n120 & n123 ;
  assign n250 = ~n125 ;
  assign n126 = n124 & n250 ;
  assign n127 = n102 | n126 ;
  assign n128 = n102 & n126 ;
  assign n251 = ~n128 ;
  assign n22 = n127 & n251 ;
  assign n132 = n49 & n104 ;
  assign n133 = n50 | n132 ;
  assign n252 = ~n118 ;
  assign n134 = n116 & n252 ;
  assign n253 = ~n133 ;
  assign n135 = n253 & n134 ;
  assign n254 = ~n134 ;
  assign n136 = n133 & n254 ;
  assign n137 = n135 | n136 ;
  assign n37 = x0 & x14 ;
  assign n36 = x4 & x10 ;
  assign n33 = x3 & x11 ;
  assign n34 = x6 & x9 ;
  assign n255 = ~n31 ;
  assign n138 = n30 & n255 ;
  assign n139 = n34 & n138 ;
  assign n52 = x5 & x9 ;
  assign n53 = x6 & x8 ;
  assign n140 = n52 | n53 ;
  assign n256 = ~n139 ;
  assign n141 = n256 & n140 ;
  assign n142 = n110 & n141 ;
  assign n144 = n110 | n141 ;
  assign n257 = ~x6 ;
  assign n143 = n257 & n25 ;
  assign n145 = n52 & n143 ;
  assign n258 = ~n145 ;
  assign n146 = n144 & n258 ;
  assign n259 = ~n142 ;
  assign n147 = n259 & n146 ;
  assign n148 = n33 & n147 ;
  assign n149 = n33 | n147 ;
  assign n260 = ~n148 ;
  assign n150 = n260 & n149 ;
  assign n35 = x1 & x13 ;
  assign n261 = ~n48 ;
  assign n94 = n35 & n261 ;
  assign n262 = ~n35 ;
  assign n151 = n262 & n48 ;
  assign n152 = n94 | n151 ;
  assign n153 = n150 | n152 ;
  assign n154 = n150 & n152 ;
  assign n263 = ~n154 ;
  assign n155 = n153 & n263 ;
  assign n156 = n36 & n155 ;
  assign n157 = n36 | n155 ;
  assign n264 = ~n156 ;
  assign n158 = n264 & n157 ;
  assign n265 = ~n158 ;
  assign n159 = n37 & n265 ;
  assign n266 = ~n37 ;
  assign n160 = n266 & n158 ;
  assign n161 = n159 | n160 ;
  assign n162 = n137 | n161 ;
  assign n163 = n137 & n161 ;
  assign n267 = ~n163 ;
  assign n164 = n162 & n267 ;
  assign n129 = n96 | n125 ;
  assign n130 = n251 & n129 ;
  assign n165 = n249 & n128 ;
  assign n166 = n130 | n165 ;
  assign n268 = ~n164 ;
  assign n167 = n268 & n166 ;
  assign n269 = ~n166 ;
  assign n216 = n164 & n269 ;
  assign n23 = n167 | n216 ;
  assign n131 = n128 | n129 ;
  assign n270 = ~n167 ;
  assign n168 = n131 & n270 ;
  assign n54 = x2 & x13 ;
  assign n169 = n240 & n54 ;
  assign n170 = n168 & n169 ;
  assign n171 = n168 | n169 ;
  assign n271 = ~n170 ;
  assign n172 = n271 & n171 ;
  assign n55 = x4 & x11 ;
  assign n38 = x0 & x15 ;
  assign n272 = ~n30 ;
  assign n173 = n272 & n34 ;
  assign n273 = ~n173 ;
  assign n174 = n38 & n273 ;
  assign n274 = ~n38 ;
  assign n175 = n274 & n173 ;
  assign n176 = n174 | n175 ;
  assign n177 = n55 | n176 ;
  assign n178 = n55 & n176 ;
  assign n275 = ~n178 ;
  assign n179 = n177 & n275 ;
  assign n180 = n172 & n179 ;
  assign n181 = n172 | n179 ;
  assign n276 = ~n180 ;
  assign n182 = n276 & n181 ;
  assign n39 = x5 & x10 ;
  assign n277 = ~n36 ;
  assign n183 = n277 & n155 ;
  assign n278 = ~n183 ;
  assign n184 = n153 & n278 ;
  assign n185 = n39 & n184 ;
  assign n186 = n39 | n184 ;
  assign n279 = ~n185 ;
  assign n187 = n279 & n186 ;
  assign n188 = n133 & n134 ;
  assign n189 = n163 | n188 ;
  assign n40 = x7 & x8 ;
  assign n56 = x3 & x12 ;
  assign n280 = ~n56 ;
  assign n190 = n40 & n280 ;
  assign n281 = ~n40 ;
  assign n191 = n281 & n56 ;
  assign n192 = n190 | n191 ;
  assign n282 = ~n192 ;
  assign n193 = n189 & n282 ;
  assign n283 = ~n189 ;
  assign n194 = n283 & n192 ;
  assign n195 = n193 | n194 ;
  assign n284 = ~n195 ;
  assign n196 = n187 & n284 ;
  assign n285 = ~n187 ;
  assign n197 = n285 & n195 ;
  assign n198 = n196 | n197 ;
  assign n286 = ~n33 ;
  assign n199 = n286 & n147 ;
  assign n287 = ~n199 ;
  assign n200 = n144 & n287 ;
  assign n201 = x0 & n158 ;
  assign n202 = x1 & n201 ;
  assign n203 = x1 | n201 ;
  assign n204 = x14 & n203 ;
  assign n288 = ~n202 ;
  assign n205 = n288 & n204 ;
  assign n289 = ~n200 ;
  assign n206 = n289 & n205 ;
  assign n290 = ~n205 ;
  assign n207 = n200 & n290 ;
  assign n208 = n206 | n207 ;
  assign n209 = n198 | n208 ;
  assign n210 = n198 & n208 ;
  assign n291 = ~n210 ;
  assign n211 = n209 & n291 ;
  assign n212 = n182 & n211 ;
  assign n213 = n182 | n211 ;
  assign n292 = ~n212 ;
  assign n24 = n292 & n213 ;
  assign y0 = n17 ;
  assign y1 = n18 ;
  assign y2 = n19 ;
  assign y3 = n20 ;
  assign y4 = n21 ;
  assign y5 = n22 ;
  assign y6 = n23 ;
  assign y7 = n24 ;
endmodule
