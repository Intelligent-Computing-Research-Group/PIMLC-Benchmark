module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 ;
  assign n52 = x8 | x9 ;
  assign n25 = x4 | x7 ;
  assign n403 = ~x0 ;
  assign n39 = n403 & x1 ;
  assign n404 = ~x9 ;
  assign n117 = n404 & n39 ;
  assign n118 = x2 | n117 ;
  assign n405 = ~x1 ;
  assign n82 = n405 & x9 ;
  assign n119 = n403 & x8 ;
  assign n120 = n82 | n119 ;
  assign n121 = n118 | n120 ;
  assign n102 = n403 & x5 ;
  assign n515 = x2 & x8 ;
  assign n350 = x5 & x8 ;
  assign n303 = x2 & x9 ;
  assign n354 = x8 & x9 ;
  assign n122 = n303 | n354 ;
  assign n406 = ~n350 ;
  assign n123 = n406 & n122 ;
  assign n124 = n515 | n123 ;
  assign n407 = ~x6 ;
  assign n125 = n407 & n124 ;
  assign n126 = n102 | n125 ;
  assign n408 = ~n121 ;
  assign n127 = n408 & n126 ;
  assign n409 = ~x5 ;
  assign n68 = x1 & n409 ;
  assign n97 = n404 & n68 ;
  assign n410 = ~x8 ;
  assign n98 = x2 & n410 ;
  assign n99 = n97 & n98 ;
  assign n100 = x2 & n406 ;
  assign n45 = x3 | x9 ;
  assign n60 = x1 & n407 ;
  assign n101 = n45 & n60 ;
  assign n411 = ~n100 ;
  assign n104 = n411 & n101 ;
  assign n103 = x3 | x6 ;
  assign n412 = ~n102 ;
  assign n105 = n412 & n103 ;
  assign n106 = n104 | n105 ;
  assign n107 = n99 | n106 ;
  assign n29 = x1 | x5 ;
  assign n413 = ~n29 ;
  assign n129 = n354 & n413 ;
  assign n130 = n107 | n129 ;
  assign n131 = x0 | x1 ;
  assign n414 = ~n131 ;
  assign n132 = x2 & n414 ;
  assign n415 = ~x2 ;
  assign n135 = n415 & n117 ;
  assign n136 = n132 | n135 ;
  assign n137 = n130 & n136 ;
  assign n138 = n127 | n137 ;
  assign n416 = ~x3 ;
  assign n139 = n416 & n138 ;
  assign n140 = n403 & x2 ;
  assign n141 = n415 & n131 ;
  assign n142 = x1 | n141 ;
  assign n143 = x3 | n142 ;
  assign n144 = x5 & n143 ;
  assign n145 = n140 | n144 ;
  assign n146 = x6 | x9 ;
  assign n147 = n415 & x8 ;
  assign n360 = x1 & x3 ;
  assign n148 = x0 & n360 ;
  assign n417 = ~n147 ;
  assign n149 = n417 & n148 ;
  assign n150 = n146 | n149 ;
  assign n418 = ~n150 ;
  assign n151 = n145 & n418 ;
  assign n27 = x6 | x8 ;
  assign n28 = x3 & n407 ;
  assign n30 = x0 | n29 ;
  assign n31 = n28 | n30 ;
  assign n32 = n27 & n31 ;
  assign n33 = n303 & n360 ;
  assign n377 = x2 & x6 ;
  assign n35 = x2 | x9 ;
  assign n419 = ~n377 ;
  assign n36 = n419 & n35 ;
  assign n420 = ~n33 ;
  assign n37 = n420 & n36 ;
  assign n421 = ~n32 ;
  assign n38 = n421 & n37 ;
  assign n40 = n303 | n39 ;
  assign n41 = n360 | n40 ;
  assign n42 = x5 | x8 ;
  assign n422 = ~n42 ;
  assign n43 = n41 & n422 ;
  assign n44 = n38 | n43 ;
  assign n516 = x5 & x6 ;
  assign n423 = ~n516 ;
  assign n152 = x8 & n423 ;
  assign n386 = x0 & x1 ;
  assign n154 = x9 & n386 ;
  assign n77 = x2 | x3 ;
  assign n155 = x9 & n77 ;
  assign n156 = n154 | n155 ;
  assign n424 = ~n152 ;
  assign n157 = n424 & n156 ;
  assign n425 = ~n44 ;
  assign n158 = n425 & n157 ;
  assign n34 = x6 & n33 ;
  assign n51 = x5 | n354 ;
  assign n324 = x3 & x8 ;
  assign n426 = ~n324 ;
  assign n53 = n426 & n52 ;
  assign n54 = n51 | n53 ;
  assign n55 = x0 & n409 ;
  assign n427 = ~n35 ;
  assign n56 = n427 & n55 ;
  assign n428 = ~n56 ;
  assign n57 = n54 & n428 ;
  assign n58 = n415 & x3 ;
  assign n59 = n27 & n58 ;
  assign n61 = x3 & n410 ;
  assign n62 = n405 & x6 ;
  assign n429 = ~n61 ;
  assign n63 = n429 & n62 ;
  assign n64 = n60 | n63 ;
  assign n65 = n59 | n64 ;
  assign n430 = ~n57 ;
  assign n66 = n430 & n65 ;
  assign n173 = n34 | n66 ;
  assign n88 = x0 & n404 ;
  assign n159 = n413 & n88 ;
  assign n162 = n410 & n159 ;
  assign n46 = x6 & n410 ;
  assign n161 = x0 | n46 ;
  assign n431 = ~n161 ;
  assign n163 = n97 & n431 ;
  assign n164 = n162 | n163 ;
  assign n166 = x8 | n164 ;
  assign n432 = ~n68 ;
  assign n69 = x6 & n432 ;
  assign n70 = x9 | n69 ;
  assign n167 = x5 | x6 ;
  assign n168 = x0 & n82 ;
  assign n169 = n167 & n168 ;
  assign n433 = ~n169 ;
  assign n170 = n70 & n433 ;
  assign n171 = n426 & n77 ;
  assign n434 = ~n170 ;
  assign n172 = n434 & n171 ;
  assign n174 = n166 & n172 ;
  assign n175 = n173 | n174 ;
  assign n176 = n158 | n175 ;
  assign n177 = n151 | n176 ;
  assign n178 = n139 | n177 ;
  assign n435 = ~n25 ;
  assign n378 = n435 & n178 ;
  assign n436 = ~n52 ;
  assign n379 = n436 & n378 ;
  assign n288 = x2 & x3 ;
  assign n437 = ~n288 ;
  assign n83 = n437 & n77 ;
  assign n84 = n82 | n83 ;
  assign n438 = ~n386 ;
  assign n85 = x9 & n438 ;
  assign n86 = x9 | n39 ;
  assign n439 = ~n85 ;
  assign n87 = n439 & n86 ;
  assign n440 = ~n84 ;
  assign n90 = n440 & n87 ;
  assign n89 = n77 | n88 ;
  assign n91 = x6 & n89 ;
  assign n92 = n90 | n91 ;
  assign n93 = n435 & n92 ;
  assign n81 = x1 | n77 ;
  assign n277 = x7 | n81 ;
  assign n279 = n403 & x4 ;
  assign n441 = ~n277 ;
  assign n280 = n441 & n279 ;
  assign n353 = n516 & n280 ;
  assign n442 = ~n353 ;
  assign n387 = x8 & n442 ;
  assign n443 = ~n93 ;
  assign n388 = n443 & n387 ;
  assign n281 = n423 & n280 ;
  assign n390 = x8 | n281 ;
  assign n444 = ~n77 ;
  assign n80 = x6 & n444 ;
  assign n327 = n416 & x9 ;
  assign n328 = n80 | n327 ;
  assign n389 = n403 & n328 ;
  assign n391 = x5 | n389 ;
  assign n392 = n390 & n391 ;
  assign n445 = ~n388 ;
  assign n396 = n445 & n392 ;
  assign n76 = n288 & n55 ;
  assign n94 = n77 | n92 ;
  assign n446 = ~n76 ;
  assign n95 = n446 & n94 ;
  assign n447 = ~n95 ;
  assign n160 = n447 & n159 ;
  assign n393 = x1 | n155 ;
  assign n394 = n44 & n393 ;
  assign n395 = n160 | n394 ;
  assign n397 = n435 & n395 ;
  assign n398 = n396 | n397 ;
  assign n399 = n379 | n398 ;
  assign n197 = x2 | n68 ;
  assign n448 = ~n130 ;
  assign n198 = n448 & n197 ;
  assign n449 = ~n46 ;
  assign n47 = n45 & n449 ;
  assign n450 = ~n47 ;
  assign n48 = n39 & n450 ;
  assign n451 = ~n48 ;
  assign n49 = n44 & n451 ;
  assign n452 = ~n49 ;
  assign n50 = n288 & n452 ;
  assign n67 = x3 | n66 ;
  assign n71 = n350 | n70 ;
  assign n72 = n403 & n71 ;
  assign n73 = n67 & n72 ;
  assign n74 = n48 | n73 ;
  assign n453 = ~n50 ;
  assign n75 = n453 & n74 ;
  assign n229 = n57 & n75 ;
  assign n78 = n436 & n77 ;
  assign n216 = n419 & n52 ;
  assign n217 = n78 | n216 ;
  assign n454 = ~n217 ;
  assign n218 = x1 & n454 ;
  assign n219 = n92 & n218 ;
  assign n220 = n430 & n219 ;
  assign n221 = x2 | x6 ;
  assign n455 = ~n221 ;
  assign n224 = x8 & n455 ;
  assign n225 = n84 | n224 ;
  assign n226 = n426 & n225 ;
  assign n456 = ~n226 ;
  assign n227 = n55 & n456 ;
  assign n457 = ~n125 ;
  assign n228 = n457 & n227 ;
  assign n458 = ~n220 ;
  assign n230 = n458 & n228 ;
  assign n231 = n229 | n230 ;
  assign n368 = n198 | n231 ;
  assign n190 = x5 & n360 ;
  assign n191 = n416 & n68 ;
  assign n192 = n190 | n191 ;
  assign n459 = ~n354 ;
  assign n207 = n459 & n52 ;
  assign n369 = x0 & n407 ;
  assign n460 = ~n98 ;
  assign n370 = n460 & n369 ;
  assign n461 = ~n207 ;
  assign n371 = n461 & n370 ;
  assign n372 = n81 & n371 ;
  assign n373 = n75 | n372 ;
  assign n462 = ~n192 ;
  assign n374 = n462 & n373 ;
  assign n375 = n368 | n374 ;
  assign n376 = n435 & n375 ;
  assign n267 = x4 | x5 ;
  assign n268 = n103 | n267 ;
  assign n208 = n405 & n207 ;
  assign n299 = n140 & n208 ;
  assign n463 = ~n299 ;
  assign n318 = n121 & n463 ;
  assign n319 = n268 | n318 ;
  assign n400 = n157 | n319 ;
  assign n401 = n376 | n400 ;
  assign n464 = ~n399 ;
  assign n402 = n464 & n401 ;
  assign n23 = x6 & x9 ;
  assign n465 = ~n23 ;
  assign n248 = n465 & n146 ;
  assign n466 = ~n248 ;
  assign n380 = n57 & n466 ;
  assign n381 = n280 & n380 ;
  assign n382 = n378 | n381 ;
  assign n269 = x2 & n131 ;
  assign n270 = n268 | n269 ;
  assign n467 = ~n270 ;
  assign n383 = n25 & n467 ;
  assign n468 = ~n219 ;
  assign n384 = n468 & n383 ;
  assign n385 = n368 & n384 ;
  assign n12 = n382 | n385 ;
  assign n115 = x8 & n404 ;
  assign n469 = ~n115 ;
  assign n361 = n469 & n130 ;
  assign n470 = ~n361 ;
  assign n365 = n280 & n470 ;
  assign n128 = x7 & n127 ;
  assign n271 = n128 | n164 ;
  assign n362 = x2 & n25 ;
  assign n471 = ~n515 ;
  assign n363 = n471 & n268 ;
  assign n364 = n362 | n363 ;
  assign n472 = ~n364 ;
  assign n366 = n271 & n472 ;
  assign n367 = n365 | n366 ;
  assign n13 = n367 | n376 ;
  assign n153 = n516 | n125 ;
  assign n358 = n153 & n280 ;
  assign n96 = n75 | n95 ;
  assign n108 = n39 & n107 ;
  assign n109 = x3 & n459 ;
  assign n473 = ~n39 ;
  assign n110 = n473 & n109 ;
  assign n111 = x6 | n110 ;
  assign n112 = n108 | n111 ;
  assign n113 = n96 & n112 ;
  assign n116 = n288 & n469 ;
  assign n179 = n350 | n102 ;
  assign n180 = n35 | n119 ;
  assign n181 = n179 | n180 ;
  assign n474 = ~n181 ;
  assign n182 = n178 & n474 ;
  assign n183 = n116 | n182 ;
  assign n184 = n405 & n183 ;
  assign n185 = n113 | n184 ;
  assign n186 = n516 & n131 ;
  assign n475 = ~n186 ;
  assign n236 = n185 & n475 ;
  assign n187 = x8 & n87 ;
  assign n188 = x3 | n187 ;
  assign n189 = n141 & n188 ;
  assign n165 = x3 & n164 ;
  assign n193 = n459 & n360 ;
  assign n194 = n386 & n462 ;
  assign n195 = n193 | n194 ;
  assign n196 = n182 & n195 ;
  assign n199 = n182 | n195 ;
  assign n476 = ~n198 ;
  assign n200 = n476 & n199 ;
  assign n477 = ~n196 ;
  assign n201 = n477 & n200 ;
  assign n202 = n165 | n201 ;
  assign n203 = n386 & n436 ;
  assign n478 = ~n203 ;
  assign n204 = x2 & n478 ;
  assign n479 = ~n202 ;
  assign n205 = n479 & n204 ;
  assign n206 = n189 | n205 ;
  assign n212 = x5 & n407 ;
  assign n209 = x1 & n354 ;
  assign n210 = n77 & n209 ;
  assign n211 = n208 | n210 ;
  assign n213 = n437 & n211 ;
  assign n480 = ~n213 ;
  assign n214 = n212 & n480 ;
  assign n215 = n206 & n214 ;
  assign n481 = ~n103 ;
  assign n232 = n481 & n122 ;
  assign n482 = ~n232 ;
  assign n233 = n386 & n482 ;
  assign n483 = ~n231 ;
  assign n234 = n483 & n233 ;
  assign n484 = ~n182 ;
  assign n235 = n484 & n234 ;
  assign n485 = ~n215 ;
  assign n237 = n485 & n235 ;
  assign n238 = n236 | n237 ;
  assign n359 = n435 & n238 ;
  assign n14 = n358 | n359 ;
  assign n351 = n516 & n435 ;
  assign n134 = n58 | n131 ;
  assign n486 = ~n141 ;
  assign n355 = n134 & n486 ;
  assign n356 = n351 & n355 ;
  assign n15 = n353 | n356 ;
  assign n133 = x2 | n131 ;
  assign n244 = x3 & n133 ;
  assign n352 = n244 & n351 ;
  assign n16 = n352 | n353 ;
  assign n256 = x2 & n481 ;
  assign n487 = ~n119 ;
  assign n246 = n68 & n487 ;
  assign n257 = n80 & n246 ;
  assign n258 = n256 | n257 ;
  assign n259 = n72 & n258 ;
  assign n260 = n219 | n259 ;
  assign n114 = x0 & n113 ;
  assign n245 = n61 | n244 ;
  assign n249 = n103 & n248 ;
  assign n250 = n303 | n249 ;
  assign n251 = n409 & n250 ;
  assign n252 = n246 | n251 ;
  assign n253 = n245 | n252 ;
  assign n254 = n414 & n253 ;
  assign n255 = n114 | n254 ;
  assign n261 = n354 & n255 ;
  assign n262 = n260 | n261 ;
  assign n263 = n202 | n262 ;
  assign n22 = x2 & n350 ;
  assign n240 = n45 | n119 ;
  assign n241 = n22 | n240 ;
  assign n239 = n405 & n51 ;
  assign n242 = x8 | n239 ;
  assign n488 = ~n241 ;
  assign n243 = n488 & n242 ;
  assign n489 = ~n238 ;
  assign n264 = n489 & n243 ;
  assign n265 = n263 | n264 ;
  assign n266 = n435 & n265 ;
  assign n272 = x7 & n404 ;
  assign n273 = n417 & n272 ;
  assign n274 = n98 | n273 ;
  assign n275 = n271 | n274 ;
  assign n276 = n467 & n275 ;
  assign n490 = ~x7 ;
  assign n282 = n490 & n516 ;
  assign n283 = n280 | n282 ;
  assign n284 = n276 | n283 ;
  assign n285 = n266 | n284 ;
  assign n222 = n88 | n221 ;
  assign n491 = ~n222 ;
  assign n223 = n109 & n491 ;
  assign n329 = n98 & n327 ;
  assign n330 = n377 & n52 ;
  assign n331 = n329 | n330 ;
  assign n332 = n223 | n331 ;
  assign n357 = x3 & x6 ;
  assign n492 = ~n357 ;
  assign n325 = n492 & n35 ;
  assign n326 = x0 | n207 ;
  assign n333 = n325 | n326 ;
  assign n493 = ~n332 ;
  assign n334 = n493 & n333 ;
  assign n335 = n29 | n334 ;
  assign n336 = n459 & n146 ;
  assign n337 = x3 | n336 ;
  assign n79 = n52 | n77 ;
  assign n338 = n415 & x6 ;
  assign n339 = n79 & n338 ;
  assign n494 = ~n339 ;
  assign n340 = n337 & n494 ;
  assign n495 = ~n340 ;
  assign n341 = n142 & n495 ;
  assign n342 = n39 & n147 ;
  assign n343 = n341 | n342 ;
  assign n344 = n252 & n343 ;
  assign n496 = ~n344 ;
  assign n345 = n335 & n496 ;
  assign n346 = n485 & n345 ;
  assign n347 = n25 | n346 ;
  assign n26 = x2 & n435 ;
  assign n286 = n26 & n202 ;
  assign n287 = n280 | n286 ;
  assign n497 = ~n167 ;
  assign n21 = n497 & n287 ;
  assign n278 = n208 & n277 ;
  assign n498 = ~n319 ;
  assign n348 = n278 & n498 ;
  assign n349 = n21 | n348 ;
  assign n499 = ~n349 ;
  assign n18 = n347 & n499 ;
  assign n289 = n245 & n252 ;
  assign n500 = ~n289 ;
  assign n290 = x6 & n500 ;
  assign n501 = ~n253 ;
  assign n291 = n354 & n501 ;
  assign n292 = n25 | n291 ;
  assign n293 = n290 | n292 ;
  assign n502 = ~n45 ;
  assign n247 = n502 & n246 ;
  assign n304 = x2 & n28 ;
  assign n503 = ~n246 ;
  assign n305 = n503 & n304 ;
  assign n504 = ~n164 ;
  assign n306 = n504 & n305 ;
  assign n307 = n247 | n306 ;
  assign n24 = x5 & n354 ;
  assign n294 = n52 & n239 ;
  assign n295 = x3 & n294 ;
  assign n308 = n24 | n295 ;
  assign n505 = ~n294 ;
  assign n309 = n221 & n505 ;
  assign n310 = n308 | n309 ;
  assign n506 = ~n307 ;
  assign n311 = n506 & n310 ;
  assign n312 = n408 & n179 ;
  assign n507 = ~n195 ;
  assign n313 = n507 & n312 ;
  assign n314 = n311 | n313 ;
  assign n508 = ~n310 ;
  assign n315 = n307 & n508 ;
  assign n316 = n314 | n315 ;
  assign n509 = ~n293 ;
  assign n317 = n509 & n316 ;
  assign n510 = ~n208 ;
  assign n320 = x0 & n510 ;
  assign n321 = n319 | n320 ;
  assign n322 = n409 & n280 ;
  assign n511 = ~n322 ;
  assign n323 = n321 & n511 ;
  assign n512 = ~n317 ;
  assign n19 = n512 & n323 ;
  assign n296 = x2 & n505 ;
  assign n297 = n67 | n296 ;
  assign n298 = n509 & n297 ;
  assign n513 = ~n268 ;
  assign n300 = n513 & n299 ;
  assign n301 = n281 | n300 ;
  assign n302 = n298 | n301 ;
  assign n514 = ~n21 ;
  assign n20 = n514 & n302 ;
  assign n11 = ~n402 ;
  assign n17 = ~n285 ;
  assign y0 = n11 ;
  assign y1 = n12 ;
  assign y2 = n13 ;
  assign y3 = n14 ;
  assign y4 = n15 ;
  assign y5 = n16 ;
  assign y6 = n17 ;
  assign y7 = n18 ;
  assign y8 = n19 ;
  assign y9 = n20 ;
  assign y10 = n21 ;
endmodule
