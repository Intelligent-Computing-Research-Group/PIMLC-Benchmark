module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 ;
  assign n25 = x5 | x6 ;
  assign n128 = x5 & x6 ;
  assign n150 = ~n128 ;
  assign n26 = x9 & n150 ;
  assign n28 = n25 & n26 ;
  assign n146 = x1 & x2 ;
  assign n35 = x1 | x2 ;
  assign n151 = ~n146 ;
  assign n36 = n151 & n35 ;
  assign n38 = x6 | x7 ;
  assign n152 = ~x8 ;
  assign n41 = x5 & n152 ;
  assign n153 = ~n38 ;
  assign n43 = n153 & n41 ;
  assign n44 = n36 & n43 ;
  assign n45 = n28 | n44 ;
  assign n144 = x4 & x5 ;
  assign n31 = x4 | x5 ;
  assign n154 = ~n144 ;
  assign n32 = n154 & n31 ;
  assign n155 = ~n32 ;
  assign n33 = x8 & n155 ;
  assign n34 = x9 | n33 ;
  assign n40 = x3 & n38 ;
  assign n149 = x4 & x7 ;
  assign n156 = ~x7 ;
  assign n49 = x6 & n156 ;
  assign n50 = x2 & n49 ;
  assign n52 = n149 | n50 ;
  assign n157 = ~n52 ;
  assign n53 = n40 & n157 ;
  assign n158 = ~x3 ;
  assign n54 = n158 & n52 ;
  assign n55 = n53 | n54 ;
  assign n91 = x1 & x4 ;
  assign n159 = ~x0 ;
  assign n141 = n159 & n91 ;
  assign n160 = ~n91 ;
  assign n29 = x0 & n160 ;
  assign n30 = n141 | n29 ;
  assign n71 = x5 | n38 ;
  assign n161 = ~n71 ;
  assign n72 = n30 & n161 ;
  assign n73 = x8 | n72 ;
  assign n74 = n55 | n73 ;
  assign n162 = ~n34 ;
  assign n75 = n162 & n74 ;
  assign n76 = n45 | n75 ;
  assign n163 = ~x10 ;
  assign n77 = n163 & n76 ;
  assign n39 = x10 & n38 ;
  assign n134 = x8 & x9 ;
  assign n22 = x6 & x7 ;
  assign n164 = ~n134 ;
  assign n89 = n164 & n22 ;
  assign n165 = ~n89 ;
  assign n90 = n39 & n165 ;
  assign n12 = n77 | n90 ;
  assign n88 = x8 | n22 ;
  assign n92 = x8 & n22 ;
  assign n166 = ~n92 ;
  assign n93 = x10 & n166 ;
  assign n94 = n90 | n93 ;
  assign n95 = n88 & n94 ;
  assign n37 = x3 & n151 ;
  assign n167 = ~n37 ;
  assign n46 = n167 & n43 ;
  assign n47 = n158 & n146 ;
  assign n168 = ~n47 ;
  assign n48 = n46 & n168 ;
  assign n61 = x6 & n144 ;
  assign n169 = ~n61 ;
  assign n62 = x8 & n169 ;
  assign n63 = x6 | n144 ;
  assign n64 = n62 & n63 ;
  assign n56 = x3 & n52 ;
  assign n170 = ~x5 ;
  assign n19 = n170 & x7 ;
  assign n171 = ~x4 ;
  assign n51 = n171 & n49 ;
  assign n57 = n19 | n51 ;
  assign n172 = ~n57 ;
  assign n58 = n56 & n172 ;
  assign n173 = ~n56 ;
  assign n59 = n173 & n57 ;
  assign n60 = x8 | n59 ;
  assign n65 = n58 | n60 ;
  assign n174 = ~n64 ;
  assign n66 = n174 & n65 ;
  assign n67 = n48 | n66 ;
  assign n175 = ~x9 ;
  assign n68 = n175 & n67 ;
  assign n20 = x2 & x4 ;
  assign n21 = n159 & x4 ;
  assign n176 = ~n21 ;
  assign n78 = x1 & n176 ;
  assign n177 = ~n20 ;
  assign n79 = n177 & n78 ;
  assign n178 = ~n78 ;
  assign n80 = n20 & n178 ;
  assign n81 = n71 | n80 ;
  assign n82 = n79 | n81 ;
  assign n27 = n156 & n26 ;
  assign n23 = x5 & x9 ;
  assign n123 = n22 & n23 ;
  assign n124 = x10 | n123 ;
  assign n125 = n27 | n124 ;
  assign n179 = ~n125 ;
  assign n126 = n82 & n179 ;
  assign n180 = ~n68 ;
  assign n127 = n180 & n126 ;
  assign n13 = n95 | n127 ;
  assign n69 = x3 & n67 ;
  assign n70 = x4 & n69 ;
  assign n181 = ~n81 ;
  assign n83 = x2 & n181 ;
  assign n84 = n70 | n83 ;
  assign n85 = n152 & n84 ;
  assign n96 = n144 & n92 ;
  assign n86 = x6 | x8 ;
  assign n87 = x4 | n86 ;
  assign n97 = n69 | n87 ;
  assign n182 = ~n96 ;
  assign n98 = n182 & n97 ;
  assign n42 = x7 | n41 ;
  assign n99 = n42 | n61 ;
  assign n183 = ~n86 ;
  assign n100 = x3 & n183 ;
  assign n101 = n99 | n100 ;
  assign n102 = x7 & n183 ;
  assign n184 = ~n102 ;
  assign n103 = n101 & n184 ;
  assign n104 = n98 & n103 ;
  assign n105 = x10 | n104 ;
  assign n106 = n85 | n105 ;
  assign n185 = ~n93 ;
  assign n107 = n185 & n106 ;
  assign n108 = x9 | n107 ;
  assign n109 = n84 & n104 ;
  assign n119 = x9 | n109 ;
  assign n186 = ~n123 ;
  assign n129 = x8 & n186 ;
  assign n130 = n152 & n123 ;
  assign n131 = x10 | n130 ;
  assign n132 = n129 | n131 ;
  assign n187 = ~n132 ;
  assign n133 = n119 & n187 ;
  assign n188 = ~n133 ;
  assign n14 = n108 & n188 ;
  assign n136 = x2 | x3 ;
  assign n137 = n96 & n136 ;
  assign n138 = x9 | n137 ;
  assign n142 = x10 | n138 ;
  assign n189 = ~n142 ;
  assign n143 = n96 & n189 ;
  assign n145 = x9 | x10 ;
  assign n147 = n87 | n145 ;
  assign n148 = n101 | n147 ;
  assign n190 = ~n143 ;
  assign n15 = n190 & n148 ;
  assign n191 = ~x6 ;
  assign n114 = x5 & n191 ;
  assign n115 = x7 | n114 ;
  assign n192 = ~n115 ;
  assign n116 = n98 & n192 ;
  assign n193 = ~n109 ;
  assign n117 = n193 & n116 ;
  assign n118 = n109 & n115 ;
  assign n120 = x8 | x10 ;
  assign n121 = n118 | n120 ;
  assign n122 = n117 | n121 ;
  assign n135 = x7 & n187 ;
  assign n139 = n163 & n138 ;
  assign n194 = ~n135 ;
  assign n140 = n194 & n139 ;
  assign n195 = ~n140 ;
  assign n16 = n122 & n195 ;
  assign n110 = n25 | n109 ;
  assign n24 = x7 | x8 ;
  assign n111 = x6 & n109 ;
  assign n112 = n24 | n111 ;
  assign n196 = ~n112 ;
  assign n113 = n110 & n196 ;
  assign n17 = n113 | n142 ;
  assign n18 = n112 | n145 ;
  assign y0 = n12 ;
  assign y1 = n13 ;
  assign y2 = n14 ;
  assign y3 = n15 ;
  assign y4 = n16 ;
  assign y5 = n17 ;
  assign y6 = n18 ;
endmodule
