module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 ;
  assign n141 = x0 & x16 ;
  assign n56 = x0 | x16 ;
  assign n152 = ~n141 ;
  assign n33 = n152 & n56 ;
  assign n151 = x1 & x17 ;
  assign n79 = x1 | x17 ;
  assign n153 = ~n151 ;
  assign n80 = n153 & n79 ;
  assign n81 = n152 & n80 ;
  assign n154 = ~n80 ;
  assign n82 = n141 & n154 ;
  assign n34 = n81 | n82 ;
  assign n83 = x2 & x18 ;
  assign n77 = x2 | x18 ;
  assign n155 = ~n83 ;
  assign n78 = n155 & n77 ;
  assign n84 = n141 | n151 ;
  assign n85 = n79 & n84 ;
  assign n86 = n78 & n85 ;
  assign n150 = n78 | n85 ;
  assign n156 = ~n86 ;
  assign n35 = n156 & n150 ;
  assign n135 = x3 & x19 ;
  assign n75 = x3 | x19 ;
  assign n157 = ~n135 ;
  assign n76 = n157 & n75 ;
  assign n87 = n83 | n85 ;
  assign n88 = n77 & n87 ;
  assign n147 = n76 | n88 ;
  assign n148 = n76 & n88 ;
  assign n158 = ~n148 ;
  assign n36 = n147 & n158 ;
  assign n117 = x4 & x20 ;
  assign n73 = x4 | x20 ;
  assign n159 = ~n117 ;
  assign n74 = n159 & n73 ;
  assign n89 = n135 | n88 ;
  assign n90 = n75 & n89 ;
  assign n91 = n74 & n90 ;
  assign n145 = n74 | n90 ;
  assign n160 = ~n91 ;
  assign n37 = n160 & n145 ;
  assign n137 = x5 & x21 ;
  assign n71 = x5 | x21 ;
  assign n161 = ~n137 ;
  assign n72 = n161 & n71 ;
  assign n92 = n117 | n90 ;
  assign n93 = n73 & n92 ;
  assign n142 = n72 | n93 ;
  assign n143 = n72 & n93 ;
  assign n162 = ~n143 ;
  assign n38 = n142 & n162 ;
  assign n125 = x6 & x22 ;
  assign n69 = x6 | x22 ;
  assign n163 = ~n125 ;
  assign n70 = n163 & n69 ;
  assign n94 = n137 | n93 ;
  assign n95 = n71 & n94 ;
  assign n96 = n70 & n95 ;
  assign n140 = n70 | n95 ;
  assign n164 = ~n96 ;
  assign n39 = n164 & n140 ;
  assign n139 = x7 & x23 ;
  assign n49 = x7 | x23 ;
  assign n165 = ~n139 ;
  assign n50 = n165 & n49 ;
  assign n97 = n125 | n95 ;
  assign n98 = n69 & n97 ;
  assign n166 = ~n98 ;
  assign n99 = n50 & n166 ;
  assign n167 = ~n50 ;
  assign n138 = n167 & n98 ;
  assign n40 = n99 | n138 ;
  assign n127 = x8 & x24 ;
  assign n67 = x8 | x24 ;
  assign n168 = ~n127 ;
  assign n68 = n168 & n67 ;
  assign n169 = ~n99 ;
  assign n100 = n49 & n169 ;
  assign n101 = n68 & n100 ;
  assign n136 = n68 | n100 ;
  assign n170 = ~n101 ;
  assign n41 = n170 & n136 ;
  assign n57 = x9 & x25 ;
  assign n51 = x9 | x25 ;
  assign n171 = ~n57 ;
  assign n55 = n171 & n51 ;
  assign n102 = n127 | n100 ;
  assign n103 = n67 & n102 ;
  assign n104 = n55 | n103 ;
  assign n134 = n55 & n103 ;
  assign n172 = ~n134 ;
  assign n42 = n104 & n172 ;
  assign n129 = x10 & x26 ;
  assign n65 = x10 | x26 ;
  assign n173 = ~n129 ;
  assign n66 = n173 & n65 ;
  assign n105 = n51 & n103 ;
  assign n106 = n57 | n105 ;
  assign n107 = n66 & n106 ;
  assign n132 = n66 | n106 ;
  assign n174 = ~n107 ;
  assign n43 = n174 & n132 ;
  assign n149 = x11 & x27 ;
  assign n63 = x11 | x27 ;
  assign n175 = ~n149 ;
  assign n64 = n175 & n63 ;
  assign n108 = n129 | n106 ;
  assign n109 = n65 & n108 ;
  assign n176 = ~n109 ;
  assign n110 = n64 & n176 ;
  assign n177 = ~n64 ;
  assign n130 = n177 & n109 ;
  assign n44 = n110 | n130 ;
  assign n131 = x12 & x28 ;
  assign n61 = x12 | x28 ;
  assign n178 = ~n131 ;
  assign n62 = n178 & n61 ;
  assign n179 = ~n110 ;
  assign n111 = n63 & n179 ;
  assign n112 = n62 & n111 ;
  assign n128 = n62 | n111 ;
  assign n180 = ~n112 ;
  assign n45 = n180 & n128 ;
  assign n146 = x13 & x29 ;
  assign n52 = x13 | x29 ;
  assign n181 = ~n146 ;
  assign n60 = n181 & n52 ;
  assign n113 = n131 | n111 ;
  assign n114 = n61 & n113 ;
  assign n115 = n60 | n114 ;
  assign n116 = n60 & n114 ;
  assign n182 = ~n116 ;
  assign n46 = n115 & n182 ;
  assign n133 = x14 & x30 ;
  assign n53 = x14 | x30 ;
  assign n183 = ~n133 ;
  assign n54 = n183 & n53 ;
  assign n118 = n52 & n114 ;
  assign n119 = n146 | n118 ;
  assign n120 = n54 & n119 ;
  assign n126 = n54 | n119 ;
  assign n184 = ~n120 ;
  assign n47 = n184 & n126 ;
  assign n144 = x15 & x31 ;
  assign n58 = x15 | x31 ;
  assign n185 = ~n144 ;
  assign n59 = n185 & n58 ;
  assign n121 = n53 & n119 ;
  assign n122 = n133 | n121 ;
  assign n123 = n59 | n122 ;
  assign n124 = n59 & n122 ;
  assign n186 = ~n124 ;
  assign n48 = n123 & n186 ;
  assign y0 = n33 ;
  assign y1 = n34 ;
  assign y2 = n35 ;
  assign y3 = n36 ;
  assign y4 = n37 ;
  assign y5 = n38 ;
  assign y6 = n39 ;
  assign y7 = n40 ;
  assign y8 = n41 ;
  assign y9 = n42 ;
  assign y10 = n43 ;
  assign y11 = n44 ;
  assign y12 = n45 ;
  assign y13 = n46 ;
  assign y14 = n47 ;
  assign y15 = n48 ;
endmodule
