module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 ;
  assign n33 = x0 & x16 ;
  assign n128 = x0 & x17 ;
  assign n129 = x1 & x16 ;
  assign n141 = n128 & n129 ;
  assign n233 = n128 | n129 ;
  assign n1003 = ~n141 ;
  assign n34 = n1003 & n233 ;
  assign n170 = x2 & x18 ;
  assign n534 = x2 | x18 ;
  assign n1004 = ~n170 ;
  assign n535 = n1004 & n534 ;
  assign n1005 = ~n535 ;
  assign n536 = n33 & n1005 ;
  assign n80 = x1 & x17 ;
  assign n81 = x0 & x18 ;
  assign n173 = x2 & x16 ;
  assign n588 = n81 | n173 ;
  assign n1006 = ~n588 ;
  assign n589 = n80 & n1006 ;
  assign n1007 = ~n80 ;
  assign n590 = n1007 & n588 ;
  assign n591 = n33 | n590 ;
  assign n592 = n589 | n591 ;
  assign n1008 = ~n536 ;
  assign n35 = n1008 & n592 ;
  assign n79 = x3 & x16 ;
  assign n77 = x2 & x17 ;
  assign n78 = x0 & x19 ;
  assign n169 = n77 & n78 ;
  assign n504 = n77 | n78 ;
  assign n1009 = ~n169 ;
  assign n505 = n1009 & n504 ;
  assign n1010 = ~n505 ;
  assign n506 = n79 & n1010 ;
  assign n1011 = ~n79 ;
  assign n507 = n1011 & n505 ;
  assign n533 = n506 | n507 ;
  assign n537 = n81 | n536 ;
  assign n538 = n80 & n537 ;
  assign n539 = n170 & n33 ;
  assign n540 = n538 | n539 ;
  assign n541 = n533 | n540 ;
  assign n542 = n533 & n540 ;
  assign n1012 = ~n542 ;
  assign n553 = n541 & n1012 ;
  assign n550 = n80 & n173 ;
  assign n1013 = ~x18 ;
  assign n551 = n1013 & n550 ;
  assign n82 = x1 & x18 ;
  assign n1014 = ~n550 ;
  assign n554 = n82 & n1014 ;
  assign n555 = n551 | n554 ;
  assign n556 = n553 & n555 ;
  assign n557 = n553 | n555 ;
  assign n1015 = ~n556 ;
  assign n36 = n1015 & n557 ;
  assign n76 = x4 & x16 ;
  assign n74 = x3 & x17 ;
  assign n75 = x1 & x19 ;
  assign n168 = n74 & n75 ;
  assign n471 = n74 | n75 ;
  assign n1016 = ~n168 ;
  assign n472 = n1016 & n471 ;
  assign n473 = n76 & n472 ;
  assign n502 = n76 | n472 ;
  assign n1017 = ~n473 ;
  assign n503 = n1017 & n502 ;
  assign n1018 = ~n507 ;
  assign n508 = n504 & n1018 ;
  assign n1019 = ~n508 ;
  assign n509 = n503 & n1019 ;
  assign n1020 = ~n503 ;
  assign n525 = n1020 & n508 ;
  assign n526 = n509 | n525 ;
  assign n69 = x2 & x20 ;
  assign n511 = n69 & n81 ;
  assign n171 = x0 & x20 ;
  assign n527 = n170 | n171 ;
  assign n1021 = ~n511 ;
  assign n543 = n1021 & n527 ;
  assign n544 = n526 & n543 ;
  assign n545 = n526 | n543 ;
  assign n1022 = ~n544 ;
  assign n546 = n1022 & n545 ;
  assign n547 = n542 & n546 ;
  assign n548 = n542 | n546 ;
  assign n1023 = ~n547 ;
  assign n549 = n1023 & n548 ;
  assign n552 = n82 | n550 ;
  assign n1024 = ~n553 ;
  assign n559 = n1024 & n555 ;
  assign n1025 = ~n559 ;
  assign n560 = n552 & n1025 ;
  assign n1026 = ~n549 ;
  assign n561 = n1026 & n560 ;
  assign n1027 = ~n560 ;
  assign n562 = n549 & n1027 ;
  assign n37 = n561 | n562 ;
  assign n167 = x1 & x20 ;
  assign n72 = x0 & x21 ;
  assign n73 = x3 & x18 ;
  assign n463 = n72 | n73 ;
  assign n576 = x3 & x21 ;
  assign n464 = n576 & n81 ;
  assign n1028 = ~n464 ;
  assign n465 = n463 & n1028 ;
  assign n1029 = ~n167 ;
  assign n466 = n1029 & n465 ;
  assign n1030 = ~n465 ;
  assign n478 = n167 & n1030 ;
  assign n479 = n466 | n478 ;
  assign n165 = x2 & x19 ;
  assign n70 = x4 & x17 ;
  assign n71 = x5 & x16 ;
  assign n166 = n70 & n71 ;
  assign n431 = n70 | n71 ;
  assign n1031 = ~n166 ;
  assign n432 = n1031 & n431 ;
  assign n1032 = ~n165 ;
  assign n433 = n1032 & n432 ;
  assign n1033 = ~n432 ;
  assign n469 = n165 & n1033 ;
  assign n470 = n433 | n469 ;
  assign n1034 = ~n76 ;
  assign n474 = n1034 & n472 ;
  assign n1035 = ~n474 ;
  assign n475 = n471 & n1035 ;
  assign n476 = n470 & n475 ;
  assign n477 = n470 | n475 ;
  assign n1036 = ~n476 ;
  assign n480 = n1036 & n477 ;
  assign n1037 = ~n479 ;
  assign n481 = n1037 & n480 ;
  assign n1038 = ~n480 ;
  assign n521 = n479 & n1038 ;
  assign n522 = n481 | n521 ;
  assign n510 = n503 & n508 ;
  assign n512 = n510 & n511 ;
  assign n523 = n510 | n511 ;
  assign n1039 = ~n512 ;
  assign n524 = n1039 & n523 ;
  assign n528 = n526 & n527 ;
  assign n529 = n524 | n528 ;
  assign n530 = n522 | n529 ;
  assign n531 = n522 & n529 ;
  assign n1040 = ~n531 ;
  assign n532 = n530 & n1040 ;
  assign n1041 = ~n562 ;
  assign n564 = n548 & n1041 ;
  assign n1042 = ~n564 ;
  assign n565 = n532 & n1042 ;
  assign n1043 = ~n532 ;
  assign n566 = n1043 & n564 ;
  assign n38 = n565 | n566 ;
  assign n159 = x3 & x19 ;
  assign n64 = x5 & x17 ;
  assign n65 = x6 & x16 ;
  assign n160 = n64 & n65 ;
  assign n365 = n64 | n65 ;
  assign n1044 = ~n160 ;
  assign n366 = n1044 & n365 ;
  assign n1045 = ~n159 ;
  assign n367 = n1045 & n366 ;
  assign n1046 = ~n366 ;
  assign n429 = n159 & n1046 ;
  assign n430 = n367 | n429 ;
  assign n1047 = ~n433 ;
  assign n434 = n431 & n1047 ;
  assign n435 = n430 & n434 ;
  assign n436 = n430 | n434 ;
  assign n1048 = ~n435 ;
  assign n437 = n1048 & n436 ;
  assign n67 = x4 & x18 ;
  assign n68 = x1 & x21 ;
  assign n164 = n67 & n68 ;
  assign n418 = n67 | n68 ;
  assign n1049 = ~n164 ;
  assign n419 = n1049 & n418 ;
  assign n420 = n69 & n419 ;
  assign n438 = n69 | n419 ;
  assign n1050 = ~n420 ;
  assign n439 = n1050 & n438 ;
  assign n440 = n437 & n439 ;
  assign n461 = n437 | n439 ;
  assign n1051 = ~n440 ;
  assign n462 = n1051 & n461 ;
  assign n1052 = ~n466 ;
  assign n467 = n463 & n1052 ;
  assign n468 = n462 & n467 ;
  assign n487 = n462 | n467 ;
  assign n1053 = ~n468 ;
  assign n488 = n1053 & n487 ;
  assign n161 = x0 & x22 ;
  assign n1054 = ~n481 ;
  assign n482 = n477 & n1054 ;
  assign n1055 = ~n161 ;
  assign n483 = n1055 & n482 ;
  assign n1056 = ~n482 ;
  assign n513 = n161 & n1056 ;
  assign n514 = n483 | n513 ;
  assign n1057 = ~n514 ;
  assign n515 = n488 & n1057 ;
  assign n1058 = ~n488 ;
  assign n516 = n1058 & n514 ;
  assign n517 = n515 | n516 ;
  assign n518 = n512 | n517 ;
  assign n519 = n512 & n517 ;
  assign n1059 = ~n519 ;
  assign n520 = n518 & n1059 ;
  assign n1060 = ~n565 ;
  assign n568 = n530 & n1060 ;
  assign n569 = n520 & n568 ;
  assign n586 = n520 | n568 ;
  assign n1061 = ~n569 ;
  assign n39 = n1061 & n586 ;
  assign n60 = x6 & x17 ;
  assign n58 = x4 & x19 ;
  assign n59 = x7 & x16 ;
  assign n157 = n58 & n59 ;
  assign n338 = n58 | n59 ;
  assign n1062 = ~n157 ;
  assign n339 = n1062 & n338 ;
  assign n1063 = ~n60 ;
  assign n340 = n1063 & n339 ;
  assign n1064 = ~n339 ;
  assign n370 = n60 & n1064 ;
  assign n371 = n340 | n370 ;
  assign n61 = x5 & x18 ;
  assign n62 = x2 & x21 ;
  assign n63 = x3 & x20 ;
  assign n158 = n62 & n63 ;
  assign n360 = n62 | n63 ;
  assign n1065 = ~n158 ;
  assign n361 = n1065 & n360 ;
  assign n362 = n61 & n361 ;
  assign n363 = n61 | n361 ;
  assign n1066 = ~n362 ;
  assign n364 = n1066 & n363 ;
  assign n1067 = ~n367 ;
  assign n368 = n365 & n1067 ;
  assign n369 = n364 & n368 ;
  assign n372 = n364 | n368 ;
  assign n1068 = ~n369 ;
  assign n373 = n1068 & n372 ;
  assign n1069 = ~n371 ;
  assign n374 = n1069 & n373 ;
  assign n1070 = ~n373 ;
  assign n425 = n371 & n1070 ;
  assign n426 = n374 | n425 ;
  assign n584 = x1 & x22 ;
  assign n66 = x0 & x23 ;
  assign n163 = n584 & n66 ;
  assign n416 = n584 | n66 ;
  assign n1071 = ~n163 ;
  assign n417 = n1071 & n416 ;
  assign n1072 = ~n69 ;
  assign n421 = n1072 & n419 ;
  assign n1073 = ~n421 ;
  assign n422 = n418 & n1073 ;
  assign n1074 = ~n417 ;
  assign n423 = n1074 & n422 ;
  assign n1075 = ~n422 ;
  assign n427 = n417 & n1075 ;
  assign n428 = n423 | n427 ;
  assign n441 = n435 | n440 ;
  assign n442 = n428 | n441 ;
  assign n443 = n428 & n441 ;
  assign n1076 = ~n443 ;
  assign n444 = n442 & n1076 ;
  assign n1077 = ~n444 ;
  assign n445 = n426 & n1077 ;
  assign n1078 = ~n426 ;
  assign n492 = n1078 & n444 ;
  assign n493 = n445 | n492 ;
  assign n485 = n161 & n482 ;
  assign n486 = n468 & n485 ;
  assign n484 = n161 | n482 ;
  assign n489 = n485 | n488 ;
  assign n490 = n484 & n489 ;
  assign n491 = n468 | n490 ;
  assign n1079 = ~n486 ;
  assign n498 = n1079 & n491 ;
  assign n499 = n493 | n498 ;
  assign n500 = n493 & n498 ;
  assign n1080 = ~n500 ;
  assign n501 = n499 & n1080 ;
  assign n570 = n519 | n569 ;
  assign n571 = n501 | n570 ;
  assign n572 = n501 & n570 ;
  assign n1081 = ~n572 ;
  assign n40 = n571 & n1081 ;
  assign n155 = x7 & x17 ;
  assign n52 = x8 & x16 ;
  assign n53 = x5 & x19 ;
  assign n156 = n52 & n53 ;
  assign n291 = n52 | n53 ;
  assign n1082 = ~n156 ;
  assign n292 = n1082 & n291 ;
  assign n1083 = ~n155 ;
  assign n293 = n1083 & n292 ;
  assign n1084 = ~n292 ;
  assign n330 = n155 & n1084 ;
  assign n331 = n293 | n330 ;
  assign n563 = x4 & x20 ;
  assign n567 = x6 & x18 ;
  assign n145 = n563 & n567 ;
  assign n239 = n563 | n567 ;
  assign n1085 = ~n145 ;
  assign n240 = n1085 & n239 ;
  assign n241 = n576 & n240 ;
  assign n332 = n576 | n240 ;
  assign n1086 = ~n241 ;
  assign n333 = n1086 & n332 ;
  assign n1087 = ~n333 ;
  assign n334 = n331 & n1087 ;
  assign n1088 = ~n331 ;
  assign n336 = n1088 & n333 ;
  assign n337 = n334 | n336 ;
  assign n1089 = ~n340 ;
  assign n341 = n338 & n1089 ;
  assign n1090 = ~n337 ;
  assign n342 = n1090 & n341 ;
  assign n1091 = ~n341 ;
  assign n389 = n337 & n1091 ;
  assign n390 = n342 | n389 ;
  assign n1092 = ~n374 ;
  assign n375 = n372 & n1092 ;
  assign n558 = x1 & x23 ;
  assign n143 = x0 & x24 ;
  assign n144 = x2 & x22 ;
  assign n237 = n143 | n144 ;
  assign n238 = n558 & n237 ;
  assign n376 = n1055 & n238 ;
  assign n377 = n558 | n237 ;
  assign n1093 = ~n376 ;
  assign n378 = n1093 & n377 ;
  assign n55 = x2 & x24 ;
  assign n379 = x2 | x24 ;
  assign n1094 = ~n55 ;
  assign n380 = n1094 & n379 ;
  assign n1095 = ~n380 ;
  assign n381 = n161 & n1095 ;
  assign n1096 = ~n381 ;
  assign n382 = n378 & n1096 ;
  assign n1097 = ~n61 ;
  assign n383 = n1097 & n361 ;
  assign n1098 = ~n383 ;
  assign n384 = n360 & n1098 ;
  assign n1099 = ~n382 ;
  assign n385 = n1099 & n384 ;
  assign n1100 = ~n384 ;
  assign n386 = n382 & n1100 ;
  assign n387 = n385 | n386 ;
  assign n388 = n375 | n387 ;
  assign n391 = n375 & n387 ;
  assign n1101 = ~n391 ;
  assign n392 = n388 & n1101 ;
  assign n1102 = ~n390 ;
  assign n393 = n1102 & n392 ;
  assign n1103 = ~n392 ;
  assign n448 = n390 & n1103 ;
  assign n449 = n393 | n448 ;
  assign n424 = n417 & n422 ;
  assign n446 = n426 & n444 ;
  assign n447 = n424 & n446 ;
  assign n450 = n424 | n446 ;
  assign n1104 = ~n447 ;
  assign n451 = n1104 & n450 ;
  assign n452 = n443 | n451 ;
  assign n1105 = ~n452 ;
  assign n453 = n449 & n1105 ;
  assign n1106 = ~n449 ;
  assign n459 = n1106 & n452 ;
  assign n460 = n453 | n459 ;
  assign n494 = n486 | n493 ;
  assign n495 = n491 & n494 ;
  assign n496 = n460 & n495 ;
  assign n497 = n460 | n495 ;
  assign n1107 = ~n496 ;
  assign n573 = n1107 & n497 ;
  assign n574 = n1081 & n573 ;
  assign n1108 = ~n573 ;
  assign n575 = n572 & n1108 ;
  assign n41 = n574 | n575 ;
  assign n1109 = ~n393 ;
  assign n394 = n388 & n1109 ;
  assign n1110 = ~n386 ;
  assign n395 = n378 & n1110 ;
  assign n396 = n394 & n395 ;
  assign n402 = n394 | n395 ;
  assign n1111 = ~n396 ;
  assign n403 = n1111 & n402 ;
  assign n162 = x0 & x25 ;
  assign n582 = x2 & x23 ;
  assign n585 = x3 & x24 ;
  assign n148 = n584 & n585 ;
  assign n146 = x1 & x24 ;
  assign n147 = x3 & x22 ;
  assign n245 = n146 | n147 ;
  assign n1112 = ~n148 ;
  assign n246 = n1112 & n245 ;
  assign n247 = n582 & n246 ;
  assign n248 = n582 | n246 ;
  assign n1113 = ~n247 ;
  assign n249 = n1113 & n248 ;
  assign n1114 = ~n576 ;
  assign n242 = n1114 & n240 ;
  assign n1115 = ~n242 ;
  assign n243 = n239 & n1115 ;
  assign n244 = n238 & n243 ;
  assign n250 = n238 | n243 ;
  assign n1116 = ~n244 ;
  assign n251 = n1116 & n250 ;
  assign n252 = n249 & n251 ;
  assign n346 = n249 | n251 ;
  assign n1117 = ~n252 ;
  assign n347 = n1117 & n346 ;
  assign n49 = x7 & x18 ;
  assign n50 = x4 & x21 ;
  assign n51 = x5 & x20 ;
  assign n154 = n50 & n51 ;
  assign n280 = n50 | n51 ;
  assign n1118 = ~n154 ;
  assign n281 = n1118 & n280 ;
  assign n282 = n49 & n281 ;
  assign n283 = n49 | n281 ;
  assign n1119 = ~n282 ;
  assign n284 = n1119 & n283 ;
  assign n152 = x8 & x17 ;
  assign n1000 = x9 & x16 ;
  assign n1002 = x6 & x19 ;
  assign n153 = n1000 & n1002 ;
  assign n272 = n1000 | n1002 ;
  assign n1120 = ~n153 ;
  assign n273 = n1120 & n272 ;
  assign n1121 = ~n152 ;
  assign n274 = n1121 & n273 ;
  assign n1122 = ~n273 ;
  assign n285 = n152 & n1122 ;
  assign n286 = n274 | n285 ;
  assign n1123 = ~n286 ;
  assign n287 = n284 & n1123 ;
  assign n1124 = ~n284 ;
  assign n289 = n1124 & n286 ;
  assign n290 = n287 | n289 ;
  assign n1125 = ~n293 ;
  assign n294 = n291 & n1125 ;
  assign n295 = n290 & n294 ;
  assign n328 = n290 | n294 ;
  assign n1126 = ~n295 ;
  assign n329 = n1126 & n328 ;
  assign n335 = n331 & n333 ;
  assign n343 = n337 & n341 ;
  assign n344 = n335 | n343 ;
  assign n345 = n329 | n344 ;
  assign n348 = n329 & n344 ;
  assign n1127 = ~n348 ;
  assign n349 = n345 & n1127 ;
  assign n1128 = ~n349 ;
  assign n350 = n347 & n1128 ;
  assign n1129 = ~n347 ;
  assign n351 = n1129 & n349 ;
  assign n397 = n350 | n351 ;
  assign n398 = n162 & n397 ;
  assign n401 = n162 | n397 ;
  assign n1130 = ~n398 ;
  assign n412 = n1130 & n401 ;
  assign n413 = n403 & n412 ;
  assign n414 = n403 | n412 ;
  assign n1131 = ~n413 ;
  assign n415 = n1131 & n414 ;
  assign n454 = n449 & n452 ;
  assign n455 = n447 | n454 ;
  assign n456 = n415 | n455 ;
  assign n457 = n415 & n455 ;
  assign n1132 = ~n457 ;
  assign n458 = n456 & n1132 ;
  assign n1133 = ~n574 ;
  assign n577 = n497 & n1133 ;
  assign n578 = n458 & n577 ;
  assign n583 = n458 | n577 ;
  assign n1134 = ~n578 ;
  assign n42 = n1134 & n583 ;
  assign n172 = x1 & x25 ;
  assign n234 = x0 & x26 ;
  assign n142 = n172 & n234 ;
  assign n235 = n172 | n234 ;
  assign n1135 = ~n142 ;
  assign n236 = n1135 & n235 ;
  assign n253 = n244 | n252 ;
  assign n1136 = ~n253 ;
  assign n254 = n236 & n1136 ;
  assign n1137 = ~n236 ;
  assign n256 = n1137 & n253 ;
  assign n257 = n254 | n256 ;
  assign n587 = x7 & x19 ;
  assign n593 = x9 & x17 ;
  assign n944 = x10 & x16 ;
  assign n149 = n593 & n944 ;
  assign n258 = n593 | n944 ;
  assign n1138 = ~n149 ;
  assign n259 = n1138 & n258 ;
  assign n260 = n587 & n259 ;
  assign n261 = n587 | n259 ;
  assign n1139 = ~n260 ;
  assign n262 = n1139 & n261 ;
  assign n150 = x5 & x21 ;
  assign n996 = x6 & x20 ;
  assign n998 = x8 & x18 ;
  assign n151 = n996 & n998 ;
  assign n201 = n996 | n998 ;
  assign n1140 = ~n151 ;
  assign n263 = n1140 & n201 ;
  assign n1141 = ~n150 ;
  assign n264 = n1141 & n263 ;
  assign n1142 = ~n263 ;
  assign n266 = n150 & n1142 ;
  assign n267 = n264 | n266 ;
  assign n1143 = ~n267 ;
  assign n268 = n262 & n1143 ;
  assign n1144 = ~n262 ;
  assign n270 = n1144 & n267 ;
  assign n271 = n268 | n270 ;
  assign n1145 = ~n274 ;
  assign n275 = n272 & n1145 ;
  assign n276 = n271 & n275 ;
  assign n278 = n271 | n275 ;
  assign n1146 = ~n276 ;
  assign n279 = n1146 & n278 ;
  assign n288 = n284 & n286 ;
  assign n296 = n288 | n295 ;
  assign n297 = n279 | n296 ;
  assign n298 = n279 & n296 ;
  assign n1147 = ~n298 ;
  assign n299 = n297 & n1147 ;
  assign n54 = x4 & x22 ;
  assign n57 = n582 & n585 ;
  assign n56 = x3 & x23 ;
  assign n300 = n55 | n56 ;
  assign n1148 = ~n57 ;
  assign n301 = n1148 & n300 ;
  assign n307 = n54 & n301 ;
  assign n308 = n54 | n301 ;
  assign n1149 = ~n307 ;
  assign n309 = n1149 & n308 ;
  assign n1150 = ~n49 ;
  assign n310 = n1150 & n281 ;
  assign n1151 = ~n310 ;
  assign n311 = n280 & n1151 ;
  assign n1152 = ~n582 ;
  assign n312 = n1152 & n246 ;
  assign n1153 = ~n312 ;
  assign n313 = n245 & n1153 ;
  assign n314 = n311 & n313 ;
  assign n315 = n311 | n313 ;
  assign n1154 = ~n314 ;
  assign n316 = n1154 & n315 ;
  assign n317 = n309 & n316 ;
  assign n319 = n309 | n316 ;
  assign n1155 = ~n317 ;
  assign n320 = n1155 & n319 ;
  assign n1156 = ~n299 ;
  assign n321 = n1156 & n320 ;
  assign n1157 = ~n320 ;
  assign n322 = n299 & n1157 ;
  assign n324 = n321 | n322 ;
  assign n325 = n257 | n324 ;
  assign n326 = n257 & n324 ;
  assign n1158 = ~n326 ;
  assign n327 = n325 & n1158 ;
  assign n1159 = ~n351 ;
  assign n352 = n345 & n1159 ;
  assign n353 = n327 | n352 ;
  assign n354 = n327 & n352 ;
  assign n1160 = ~n354 ;
  assign n359 = n353 & n1160 ;
  assign n399 = n396 & n398 ;
  assign n404 = n398 | n403 ;
  assign n405 = n401 & n404 ;
  assign n406 = n396 | n405 ;
  assign n1161 = ~n399 ;
  assign n408 = n1161 & n406 ;
  assign n409 = n359 | n408 ;
  assign n410 = n359 & n408 ;
  assign n1162 = ~n410 ;
  assign n411 = n409 & n1162 ;
  assign n579 = n457 | n578 ;
  assign n580 = n411 | n579 ;
  assign n581 = n411 & n579 ;
  assign n1163 = ~n581 ;
  assign n43 = n580 & n1163 ;
  assign n400 = n359 | n399 ;
  assign n407 = n400 & n406 ;
  assign n255 = n236 & n253 ;
  assign n355 = n255 & n354 ;
  assign n356 = n255 | n354 ;
  assign n1164 = ~n355 ;
  assign n357 = n1164 & n356 ;
  assign n358 = n326 | n357 ;
  assign n1165 = ~n264 ;
  assign n265 = n201 & n1165 ;
  assign n1166 = ~n54 ;
  assign n302 = n1166 & n301 ;
  assign n1167 = ~n302 ;
  assign n303 = n300 & n1167 ;
  assign n304 = n265 & n303 ;
  assign n305 = n265 | n303 ;
  assign n1168 = ~n304 ;
  assign n306 = n1168 & n305 ;
  assign n88 = x5 & x23 ;
  assign n89 = n54 & n88 ;
  assign n86 = x5 & x22 ;
  assign n87 = x4 & x23 ;
  assign n600 = n86 | n87 ;
  assign n1169 = ~n89 ;
  assign n601 = n1169 & n600 ;
  assign n602 = n585 & n601 ;
  assign n603 = n585 | n601 ;
  assign n1170 = ~n602 ;
  assign n604 = n1170 & n603 ;
  assign n1171 = ~n604 ;
  assign n605 = n306 & n1171 ;
  assign n1172 = ~n306 ;
  assign n607 = n1172 & n604 ;
  assign n608 = n605 | n607 ;
  assign n269 = n262 & n267 ;
  assign n277 = n269 | n276 ;
  assign n111 = x11 & x16 ;
  assign n109 = x8 & x19 ;
  assign n110 = x10 & x17 ;
  assign n194 = n109 & n110 ;
  assign n704 = n109 | n110 ;
  assign n1173 = ~n194 ;
  assign n705 = n1173 & n704 ;
  assign n706 = n111 & n705 ;
  assign n730 = n111 | n705 ;
  assign n1174 = ~n706 ;
  assign n731 = n1174 & n730 ;
  assign n1175 = ~n587 ;
  assign n732 = n1175 & n259 ;
  assign n1176 = ~n732 ;
  assign n733 = n258 & n1176 ;
  assign n734 = n731 & n733 ;
  assign n735 = n731 | n733 ;
  assign n1177 = ~n734 ;
  assign n736 = n1177 & n735 ;
  assign n175 = x7 & x20 ;
  assign n84 = x6 & x21 ;
  assign n85 = x9 & x18 ;
  assign n176 = n84 & n85 ;
  assign n596 = n84 | n85 ;
  assign n1178 = ~n176 ;
  assign n597 = n1178 & n596 ;
  assign n1179 = ~n175 ;
  assign n598 = n1179 & n597 ;
  assign n1180 = ~n597 ;
  assign n737 = n175 & n1180 ;
  assign n738 = n598 | n737 ;
  assign n1181 = ~n738 ;
  assign n739 = n736 & n1181 ;
  assign n1182 = ~n736 ;
  assign n740 = n1182 & n738 ;
  assign n741 = n739 | n740 ;
  assign n742 = n277 | n741 ;
  assign n743 = n277 & n741 ;
  assign n1183 = ~n743 ;
  assign n744 = n742 & n1183 ;
  assign n745 = n608 & n744 ;
  assign n746 = n608 | n744 ;
  assign n1184 = ~n745 ;
  assign n747 = n1184 & n746 ;
  assign n1185 = ~n322 ;
  assign n323 = n297 & n1185 ;
  assign n318 = n314 | n317 ;
  assign n180 = x1 & x26 ;
  assign n178 = x0 & x27 ;
  assign n179 = x2 & x25 ;
  assign n622 = n178 | n179 ;
  assign n623 = n180 | n622 ;
  assign n624 = n180 & n622 ;
  assign n1186 = ~n624 ;
  assign n625 = n623 & n1186 ;
  assign n626 = n162 | n625 ;
  assign n181 = x2 & x27 ;
  assign n920 = x2 | x27 ;
  assign n1187 = ~n181 ;
  assign n921 = n1187 & n920 ;
  assign n1188 = ~n921 ;
  assign n922 = n162 & n1188 ;
  assign n1189 = ~n922 ;
  assign n923 = n626 & n1189 ;
  assign n924 = n318 | n923 ;
  assign n925 = n318 & n923 ;
  assign n1190 = ~n925 ;
  assign n926 = n924 & n1190 ;
  assign n927 = n323 & n926 ;
  assign n928 = n323 | n926 ;
  assign n1191 = ~n927 ;
  assign n929 = n1191 & n928 ;
  assign n1192 = ~n747 ;
  assign n930 = n1192 & n929 ;
  assign n1193 = ~n929 ;
  assign n931 = n747 & n1193 ;
  assign n932 = n930 | n931 ;
  assign n933 = n358 | n932 ;
  assign n934 = n358 & n932 ;
  assign n1194 = ~n934 ;
  assign n936 = n933 & n1194 ;
  assign n937 = n407 & n936 ;
  assign n938 = n407 | n936 ;
  assign n1195 = ~n937 ;
  assign n939 = n1195 & n938 ;
  assign n942 = n581 & n939 ;
  assign n943 = n581 | n939 ;
  assign n1196 = ~n942 ;
  assign n44 = n1196 & n943 ;
  assign n940 = n1163 & n939 ;
  assign n1197 = ~n940 ;
  assign n941 = n938 & n1197 ;
  assign n935 = n355 | n934 ;
  assign n1198 = ~n930 ;
  assign n945 = n928 & n1198 ;
  assign n1199 = ~n945 ;
  assign n946 = n925 & n1199 ;
  assign n948 = n1190 & n945 ;
  assign n949 = n946 | n948 ;
  assign n748 = n743 | n745 ;
  assign n107 = x12 & x16 ;
  assign n105 = x9 & x19 ;
  assign n106 = x11 & x17 ;
  assign n189 = n105 & n106 ;
  assign n686 = n105 | n106 ;
  assign n1200 = ~n189 ;
  assign n687 = n1200 & n686 ;
  assign n688 = n107 & n687 ;
  assign n710 = n107 | n687 ;
  assign n1201 = ~n688 ;
  assign n711 = n1201 & n710 ;
  assign n186 = x7 & x21 ;
  assign n100 = x8 & x20 ;
  assign n101 = x10 & x18 ;
  assign n187 = n100 & n101 ;
  assign n669 = n100 | n101 ;
  assign n1202 = ~n187 ;
  assign n670 = n1202 & n669 ;
  assign n1203 = ~n186 ;
  assign n671 = n1203 & n670 ;
  assign n1204 = ~n670 ;
  assign n702 = n186 & n1204 ;
  assign n703 = n671 | n702 ;
  assign n1205 = ~n111 ;
  assign n707 = n1205 & n705 ;
  assign n1206 = ~n707 ;
  assign n708 = n704 & n1206 ;
  assign n709 = n703 & n708 ;
  assign n712 = n703 | n708 ;
  assign n1207 = ~n709 ;
  assign n713 = n1207 & n712 ;
  assign n1208 = ~n711 ;
  assign n714 = n1208 & n713 ;
  assign n1209 = ~n713 ;
  assign n752 = n711 & n1209 ;
  assign n753 = n714 | n752 ;
  assign n1210 = ~n598 ;
  assign n599 = n596 & n1210 ;
  assign n1211 = ~n585 ;
  assign n609 = n1211 & n601 ;
  assign n1212 = ~n609 ;
  assign n610 = n600 & n1212 ;
  assign n611 = n599 & n610 ;
  assign n612 = n599 | n610 ;
  assign n1213 = ~n611 ;
  assign n613 = n1213 & n612 ;
  assign n90 = x4 & x24 ;
  assign n91 = x6 & x22 ;
  assign n177 = n90 & n91 ;
  assign n614 = n90 | n91 ;
  assign n1214 = ~n177 ;
  assign n615 = n1214 & n614 ;
  assign n616 = n88 & n615 ;
  assign n617 = n88 | n615 ;
  assign n1215 = ~n616 ;
  assign n618 = n1215 & n617 ;
  assign n1216 = ~n618 ;
  assign n619 = n613 & n1216 ;
  assign n1217 = ~n613 ;
  assign n728 = n1217 & n618 ;
  assign n729 = n619 | n728 ;
  assign n749 = n736 & n738 ;
  assign n750 = n734 | n749 ;
  assign n751 = n729 | n750 ;
  assign n754 = n729 & n750 ;
  assign n1218 = ~n754 ;
  assign n755 = n751 & n1218 ;
  assign n1219 = ~n753 ;
  assign n756 = n1219 & n755 ;
  assign n1220 = ~n755 ;
  assign n757 = n753 & n1220 ;
  assign n758 = n756 | n757 ;
  assign n759 = n748 | n758 ;
  assign n760 = n748 & n758 ;
  assign n1221 = ~n760 ;
  assign n761 = n759 & n1221 ;
  assign n1222 = ~n605 ;
  assign n606 = n305 & n1222 ;
  assign n92 = x3 & x25 ;
  assign n93 = x1 & x27 ;
  assign n94 = x2 & x26 ;
  assign n182 = n93 & n94 ;
  assign n630 = n93 | n94 ;
  assign n1223 = ~n182 ;
  assign n631 = n1223 & n630 ;
  assign n632 = n92 & n631 ;
  assign n633 = n92 | n631 ;
  assign n1224 = ~n632 ;
  assign n634 = n1224 & n633 ;
  assign n83 = x0 & x28 ;
  assign n627 = n162 & n181 ;
  assign n628 = n624 | n627 ;
  assign n629 = n83 & n628 ;
  assign n635 = n83 | n628 ;
  assign n1225 = ~n629 ;
  assign n636 = n1225 & n635 ;
  assign n637 = n634 & n636 ;
  assign n638 = n634 | n636 ;
  assign n1226 = ~n637 ;
  assign n639 = n1226 & n638 ;
  assign n950 = n180 & n922 ;
  assign n951 = n639 & n950 ;
  assign n952 = n639 | n950 ;
  assign n1227 = ~n951 ;
  assign n953 = n1227 & n952 ;
  assign n954 = n606 & n953 ;
  assign n956 = n606 | n953 ;
  assign n1228 = ~n954 ;
  assign n957 = n1228 & n956 ;
  assign n958 = n761 & n957 ;
  assign n970 = n761 | n957 ;
  assign n1229 = ~n958 ;
  assign n971 = n1229 & n970 ;
  assign n1230 = ~n949 ;
  assign n977 = n1230 & n971 ;
  assign n1231 = ~n971 ;
  assign n978 = n949 & n1231 ;
  assign n979 = n977 | n978 ;
  assign n1232 = ~n935 ;
  assign n980 = n1232 & n979 ;
  assign n1233 = ~n979 ;
  assign n982 = n935 & n1233 ;
  assign n983 = n980 | n982 ;
  assign n984 = n941 | n983 ;
  assign n1001 = n941 & n983 ;
  assign n1234 = ~n1001 ;
  assign n45 = n984 & n1234 ;
  assign n97 = x6 & x23 ;
  assign n98 = x7 & x22 ;
  assign n99 = x5 & x24 ;
  assign n185 = n98 & n99 ;
  assign n664 = n98 | n99 ;
  assign n1235 = ~n185 ;
  assign n665 = n1235 & n664 ;
  assign n666 = n97 & n665 ;
  assign n667 = n97 | n665 ;
  assign n1236 = ~n666 ;
  assign n668 = n1236 & n667 ;
  assign n1237 = ~n671 ;
  assign n672 = n669 & n1237 ;
  assign n1238 = ~n88 ;
  assign n673 = n1238 & n615 ;
  assign n1239 = ~n673 ;
  assign n674 = n614 & n1239 ;
  assign n675 = n672 & n674 ;
  assign n676 = n672 | n674 ;
  assign n1240 = ~n675 ;
  assign n677 = n1240 & n676 ;
  assign n678 = n668 & n677 ;
  assign n679 = n668 | n677 ;
  assign n1241 = ~n678 ;
  assign n680 = n1241 & n679 ;
  assign n102 = x8 & x21 ;
  assign n103 = x11 & x18 ;
  assign n104 = x9 & x20 ;
  assign n188 = n103 & n104 ;
  assign n681 = n103 | n104 ;
  assign n1242 = ~n188 ;
  assign n682 = n1242 & n681 ;
  assign n683 = n102 & n682 ;
  assign n684 = n102 | n682 ;
  assign n1243 = ~n683 ;
  assign n685 = n1243 & n684 ;
  assign n1244 = ~n107 ;
  assign n689 = n1244 & n687 ;
  assign n1245 = ~n689 ;
  assign n690 = n686 & n1245 ;
  assign n691 = n685 & n690 ;
  assign n692 = n685 | n690 ;
  assign n1246 = ~n691 ;
  assign n693 = n1246 & n692 ;
  assign n190 = x10 & x19 ;
  assign n108 = x13 & x17 ;
  assign n193 = n107 & n108 ;
  assign n191 = x13 & x16 ;
  assign n192 = x12 & x17 ;
  assign n694 = n191 | n192 ;
  assign n1247 = ~n193 ;
  assign n695 = n1247 & n694 ;
  assign n1248 = ~n190 ;
  assign n696 = n1248 & n695 ;
  assign n1249 = ~n695 ;
  assign n697 = n190 & n1249 ;
  assign n698 = n696 | n697 ;
  assign n1250 = ~n698 ;
  assign n699 = n693 & n1250 ;
  assign n1251 = ~n693 ;
  assign n700 = n1251 & n698 ;
  assign n701 = n699 | n700 ;
  assign n715 = n711 & n713 ;
  assign n716 = n709 | n715 ;
  assign n717 = n701 | n716 ;
  assign n718 = n701 & n716 ;
  assign n1252 = ~n718 ;
  assign n719 = n717 & n1252 ;
  assign n720 = n680 & n719 ;
  assign n721 = n680 | n719 ;
  assign n1253 = ~n720 ;
  assign n722 = n1253 & n721 ;
  assign n95 = x3 & x26 ;
  assign n96 = x4 & x25 ;
  assign n183 = n95 & n96 ;
  assign n643 = n95 | n96 ;
  assign n1254 = ~n183 ;
  assign n644 = n1254 & n643 ;
  assign n645 = n1187 & n644 ;
  assign n1255 = ~n644 ;
  assign n646 = n181 & n1255 ;
  assign n647 = n645 | n646 ;
  assign n1256 = ~n92 ;
  assign n648 = n1256 & n631 ;
  assign n1257 = ~n648 ;
  assign n649 = n630 & n1257 ;
  assign n174 = x1 & x29 ;
  assign n595 = n83 & n174 ;
  assign n135 = x0 & x29 ;
  assign n184 = x1 & x28 ;
  assign n650 = n135 | n184 ;
  assign n1258 = ~n595 ;
  assign n651 = n1258 & n650 ;
  assign n652 = n649 & n651 ;
  assign n653 = n649 | n651 ;
  assign n1259 = ~n652 ;
  assign n654 = n1259 & n653 ;
  assign n655 = n647 & n654 ;
  assign n656 = n647 | n654 ;
  assign n1260 = ~n655 ;
  assign n657 = n1260 & n656 ;
  assign n620 = n613 & n618 ;
  assign n621 = n611 | n620 ;
  assign n640 = n629 | n637 ;
  assign n641 = n621 | n640 ;
  assign n642 = n621 & n640 ;
  assign n1261 = ~n642 ;
  assign n658 = n641 & n1261 ;
  assign n659 = n657 & n658 ;
  assign n723 = n657 | n658 ;
  assign n1262 = ~n659 ;
  assign n724 = n1262 & n723 ;
  assign n725 = n722 & n724 ;
  assign n726 = n722 | n724 ;
  assign n1263 = ~n725 ;
  assign n727 = n1263 & n726 ;
  assign n1264 = ~n756 ;
  assign n762 = n751 & n1264 ;
  assign n763 = n727 & n762 ;
  assign n764 = n727 | n762 ;
  assign n1265 = ~n763 ;
  assign n765 = n1265 & n764 ;
  assign n955 = n951 | n954 ;
  assign n959 = n760 | n958 ;
  assign n960 = n955 | n959 ;
  assign n961 = n955 & n959 ;
  assign n1266 = ~n961 ;
  assign n962 = n960 & n1266 ;
  assign n1267 = ~n765 ;
  assign n963 = n1267 & n962 ;
  assign n1268 = ~n962 ;
  assign n968 = n765 & n1268 ;
  assign n969 = n963 | n968 ;
  assign n947 = n925 & n945 ;
  assign n972 = n949 & n971 ;
  assign n973 = n947 | n972 ;
  assign n974 = n969 & n973 ;
  assign n975 = n969 | n973 ;
  assign n1269 = ~n974 ;
  assign n976 = n1269 & n975 ;
  assign n981 = n935 | n979 ;
  assign n1270 = ~n941 ;
  assign n985 = n1270 & n983 ;
  assign n1271 = ~n985 ;
  assign n986 = n981 & n1271 ;
  assign n1272 = ~n986 ;
  assign n987 = n976 & n1272 ;
  assign n1273 = ~n976 ;
  assign n999 = n1273 & n986 ;
  assign n46 = n987 | n999 ;
  assign n660 = n642 | n659 ;
  assign n661 = n595 | n660 ;
  assign n662 = n595 & n660 ;
  assign n1274 = ~n662 ;
  assign n663 = n661 & n1274 ;
  assign n766 = n725 | n763 ;
  assign n1275 = ~n766 ;
  assign n767 = n663 & n1275 ;
  assign n1276 = ~n663 ;
  assign n769 = n1276 & n766 ;
  assign n770 = n767 | n769 ;
  assign n1277 = ~n97 ;
  assign n771 = n1277 & n665 ;
  assign n1278 = ~n771 ;
  assign n772 = n664 & n1278 ;
  assign n1279 = ~n102 ;
  assign n773 = n1279 & n682 ;
  assign n1280 = ~n773 ;
  assign n774 = n681 & n1280 ;
  assign n775 = n772 | n774 ;
  assign n776 = n772 & n774 ;
  assign n1281 = ~n776 ;
  assign n777 = n775 & n1281 ;
  assign n195 = x6 & x24 ;
  assign n112 = x8 & x22 ;
  assign n113 = x7 & x23 ;
  assign n196 = n112 & n113 ;
  assign n216 = n112 | n113 ;
  assign n1282 = ~n196 ;
  assign n778 = n1282 & n216 ;
  assign n1283 = ~n195 ;
  assign n779 = n1283 & n778 ;
  assign n1284 = ~n778 ;
  assign n784 = n195 & n1284 ;
  assign n785 = n779 | n784 ;
  assign n786 = n777 | n785 ;
  assign n787 = n777 & n785 ;
  assign n1285 = ~n787 ;
  assign n792 = n786 & n1285 ;
  assign n793 = n675 | n678 ;
  assign n794 = n792 | n793 ;
  assign n795 = n792 & n793 ;
  assign n1286 = ~n795 ;
  assign n796 = n794 & n1286 ;
  assign n797 = n693 & n698 ;
  assign n798 = n691 | n797 ;
  assign n1287 = ~n798 ;
  assign n799 = n796 & n1287 ;
  assign n1288 = ~n796 ;
  assign n802 = n1288 & n798 ;
  assign n803 = n799 | n802 ;
  assign n1289 = ~n647 ;
  assign n804 = n1289 & n654 ;
  assign n1290 = ~n804 ;
  assign n805 = n653 & n1290 ;
  assign n1291 = ~n803 ;
  assign n807 = n1291 & n805 ;
  assign n1292 = ~n805 ;
  assign n808 = n803 & n1292 ;
  assign n809 = n807 | n808 ;
  assign n1293 = ~n680 ;
  assign n810 = n1293 & n719 ;
  assign n1294 = ~n810 ;
  assign n811 = n717 & n1294 ;
  assign n114 = x12 & x18 ;
  assign n115 = x10 & x20 ;
  assign n197 = x9 & x21 ;
  assign n1295 = ~n197 ;
  assign n812 = n115 & n1295 ;
  assign n1296 = ~n115 ;
  assign n813 = n1296 & n197 ;
  assign n814 = n812 | n813 ;
  assign n1297 = ~n814 ;
  assign n815 = n114 & n1297 ;
  assign n1298 = ~n114 ;
  assign n820 = n1298 & n814 ;
  assign n821 = n815 | n820 ;
  assign n116 = x11 & x19 ;
  assign n117 = x14 & x16 ;
  assign n198 = n116 & n117 ;
  assign n205 = n116 | n117 ;
  assign n1299 = ~n198 ;
  assign n822 = n1299 & n205 ;
  assign n831 = n108 & n822 ;
  assign n832 = n108 | n822 ;
  assign n1300 = ~n831 ;
  assign n833 = n1300 & n832 ;
  assign n1301 = ~n696 ;
  assign n834 = n694 & n1301 ;
  assign n835 = n833 & n834 ;
  assign n836 = n833 | n834 ;
  assign n1302 = ~n835 ;
  assign n837 = n1302 & n836 ;
  assign n843 = n821 & n837 ;
  assign n844 = n821 | n837 ;
  assign n1303 = ~n843 ;
  assign n845 = n1303 & n844 ;
  assign n118 = x3 & x27 ;
  assign n119 = x4 & x26 ;
  assign n120 = x5 & x25 ;
  assign n199 = n119 & n120 ;
  assign n217 = n119 | n120 ;
  assign n1304 = ~n199 ;
  assign n846 = n1304 & n217 ;
  assign n858 = n118 & n846 ;
  assign n859 = n118 | n846 ;
  assign n1305 = ~n858 ;
  assign n860 = n1305 & n859 ;
  assign n1306 = ~n645 ;
  assign n861 = n643 & n1306 ;
  assign n1307 = ~n860 ;
  assign n862 = n1307 & n861 ;
  assign n1308 = ~n861 ;
  assign n864 = n860 & n1308 ;
  assign n865 = n862 | n864 ;
  assign n200 = x2 & x28 ;
  assign n121 = x0 & x30 ;
  assign n1309 = ~n174 ;
  assign n594 = n121 & n1309 ;
  assign n1310 = ~n121 ;
  assign n866 = n1310 & n174 ;
  assign n867 = n594 | n866 ;
  assign n868 = n200 | n867 ;
  assign n869 = n200 & n867 ;
  assign n1311 = ~n869 ;
  assign n883 = n868 & n1311 ;
  assign n884 = n865 & n883 ;
  assign n890 = n865 | n883 ;
  assign n1312 = ~n884 ;
  assign n891 = n1312 & n890 ;
  assign n892 = n845 | n891 ;
  assign n894 = n845 & n891 ;
  assign n1313 = ~n894 ;
  assign n896 = n892 & n1313 ;
  assign n1314 = ~n811 ;
  assign n897 = n1314 & n896 ;
  assign n1315 = ~n896 ;
  assign n898 = n811 & n1315 ;
  assign n899 = n897 | n898 ;
  assign n900 = n809 | n899 ;
  assign n901 = n809 & n899 ;
  assign n1316 = ~n901 ;
  assign n906 = n900 & n1316 ;
  assign n907 = n770 & n906 ;
  assign n918 = n770 | n906 ;
  assign n1317 = ~n907 ;
  assign n919 = n1317 & n918 ;
  assign n1318 = ~n963 ;
  assign n964 = n960 & n1318 ;
  assign n965 = n919 & n964 ;
  assign n966 = n919 | n964 ;
  assign n1319 = ~n965 ;
  assign n967 = n1319 & n966 ;
  assign n1320 = ~n987 ;
  assign n988 = n975 & n1320 ;
  assign n1321 = ~n988 ;
  assign n989 = n967 & n1321 ;
  assign n1322 = ~n967 ;
  assign n997 = n1322 & n988 ;
  assign n47 = n989 | n997 ;
  assign n137 = x12 & x19 ;
  assign n126 = x2 & x29 ;
  assign n138 = x11 & x20 ;
  assign n1323 = ~n138 ;
  assign n218 = n126 & n1323 ;
  assign n1324 = ~n126 ;
  assign n219 = n1324 & n138 ;
  assign n220 = n218 | n219 ;
  assign n139 = x13 & x18 ;
  assign n127 = x0 & x31 ;
  assign n140 = x7 & x24 ;
  assign n1325 = ~n140 ;
  assign n221 = n127 & n1325 ;
  assign n1326 = ~n127 ;
  assign n222 = n1326 & n140 ;
  assign n223 = n221 | n222 ;
  assign n224 = n139 | n223 ;
  assign n225 = n139 & n223 ;
  assign n1327 = ~n225 ;
  assign n226 = n224 & n1327 ;
  assign n1328 = ~n220 ;
  assign n227 = n1328 & n226 ;
  assign n1329 = ~n226 ;
  assign n228 = n220 & n1329 ;
  assign n229 = n227 | n228 ;
  assign n230 = n137 | n229 ;
  assign n231 = n137 & n229 ;
  assign n1330 = ~n231 ;
  assign n232 = n230 & n1330 ;
  assign n800 = n796 & n798 ;
  assign n801 = n795 | n800 ;
  assign n131 = x6 & x25 ;
  assign n132 = x5 & x26 ;
  assign n123 = x9 & x22 ;
  assign n133 = x4 & x27 ;
  assign n1331 = ~n133 ;
  assign n206 = n123 & n1331 ;
  assign n1332 = ~n123 ;
  assign n207 = n1332 & n133 ;
  assign n208 = n206 | n207 ;
  assign n209 = n132 | n208 ;
  assign n210 = n132 & n208 ;
  assign n1333 = ~n210 ;
  assign n211 = n209 & n1333 ;
  assign n1334 = ~n131 ;
  assign n212 = n1334 & n211 ;
  assign n1335 = ~n211 ;
  assign n213 = n131 & n1335 ;
  assign n214 = n212 | n213 ;
  assign n1336 = ~n108 ;
  assign n823 = n1336 & n822 ;
  assign n1337 = ~n823 ;
  assign n824 = n205 & n1337 ;
  assign n825 = n214 | n824 ;
  assign n826 = n214 & n824 ;
  assign n1338 = ~n826 ;
  assign n827 = n825 & n1338 ;
  assign n1339 = ~n801 ;
  assign n828 = n1339 & n827 ;
  assign n1340 = ~n827 ;
  assign n829 = n801 & n1340 ;
  assign n830 = n828 | n829 ;
  assign n136 = x10 & x21 ;
  assign n816 = n114 & n814 ;
  assign n1341 = ~n136 ;
  assign n817 = n1341 & n816 ;
  assign n1342 = ~n104 ;
  assign n215 = n1342 & n136 ;
  assign n1343 = ~n816 ;
  assign n818 = n215 & n1343 ;
  assign n819 = n817 | n818 ;
  assign n124 = x14 & x17 ;
  assign n1344 = ~n779 ;
  assign n780 = n216 & n1344 ;
  assign n781 = n124 & n780 ;
  assign n782 = n124 | n780 ;
  assign n1345 = ~n781 ;
  assign n783 = n1345 & n782 ;
  assign n125 = x15 & x16 ;
  assign n1346 = ~n118 ;
  assign n847 = n1346 & n846 ;
  assign n1347 = ~n847 ;
  assign n848 = n217 & n1347 ;
  assign n1348 = ~n848 ;
  assign n849 = n125 & n1348 ;
  assign n1349 = ~n125 ;
  assign n850 = n1349 & n848 ;
  assign n851 = n849 | n850 ;
  assign n1350 = ~n851 ;
  assign n852 = n783 & n1350 ;
  assign n1351 = ~n783 ;
  assign n853 = n1351 & n851 ;
  assign n854 = n852 | n853 ;
  assign n1352 = ~n854 ;
  assign n855 = n819 & n1352 ;
  assign n1353 = ~n819 ;
  assign n856 = n1353 & n854 ;
  assign n857 = n855 | n856 ;
  assign n134 = x1 & x30 ;
  assign n870 = n135 | n869 ;
  assign n871 = n134 & n870 ;
  assign n872 = n134 | n869 ;
  assign n1354 = ~n871 ;
  assign n873 = n1354 & n872 ;
  assign n874 = n857 | n873 ;
  assign n875 = n857 & n873 ;
  assign n1355 = ~n875 ;
  assign n876 = n874 & n1355 ;
  assign n1356 = ~n830 ;
  assign n877 = n1356 & n876 ;
  assign n1357 = ~n876 ;
  assign n878 = n830 & n1357 ;
  assign n879 = n877 | n878 ;
  assign n1358 = ~n879 ;
  assign n880 = n232 & n1358 ;
  assign n1359 = ~n232 ;
  assign n881 = n1359 & n879 ;
  assign n882 = n880 | n881 ;
  assign n863 = n860 | n861 ;
  assign n1360 = ~n883 ;
  assign n885 = n865 & n1360 ;
  assign n1361 = ~n885 ;
  assign n886 = n863 & n1361 ;
  assign n887 = n1274 & n886 ;
  assign n1362 = ~n886 ;
  assign n888 = n662 & n1362 ;
  assign n889 = n887 | n888 ;
  assign n806 = n803 & n805 ;
  assign n902 = n806 | n901 ;
  assign n1363 = ~n889 ;
  assign n903 = n1363 & n902 ;
  assign n1364 = ~n902 ;
  assign n904 = n889 & n1364 ;
  assign n905 = n903 | n904 ;
  assign n893 = n811 & n892 ;
  assign n895 = n893 | n894 ;
  assign n768 = n663 & n766 ;
  assign n908 = n768 | n907 ;
  assign n909 = n895 | n908 ;
  assign n910 = n895 & n908 ;
  assign n1365 = ~n910 ;
  assign n911 = n909 & n1365 ;
  assign n1366 = ~n905 ;
  assign n912 = n1366 & n911 ;
  assign n1367 = ~n911 ;
  assign n913 = n905 & n1367 ;
  assign n914 = n912 | n913 ;
  assign n915 = n882 | n914 ;
  assign n916 = n882 & n914 ;
  assign n1368 = ~n916 ;
  assign n917 = n915 & n1368 ;
  assign n122 = x3 & x28 ;
  assign n130 = x8 & x23 ;
  assign n1369 = ~n130 ;
  assign n202 = n122 & n1369 ;
  assign n1370 = ~n122 ;
  assign n203 = n1370 & n130 ;
  assign n204 = n202 | n203 ;
  assign n788 = n776 | n787 ;
  assign n1371 = ~n204 ;
  assign n789 = n1371 & n788 ;
  assign n1372 = ~n788 ;
  assign n790 = n204 & n1372 ;
  assign n791 = n789 | n790 ;
  assign n1373 = ~n821 ;
  assign n838 = n1373 & n837 ;
  assign n1374 = ~n838 ;
  assign n839 = n836 & n1374 ;
  assign n840 = n791 | n839 ;
  assign n841 = n791 & n839 ;
  assign n1375 = ~n841 ;
  assign n842 = n840 & n1375 ;
  assign n1376 = ~n989 ;
  assign n990 = n966 & n1376 ;
  assign n991 = n842 & n990 ;
  assign n992 = n842 | n990 ;
  assign n1377 = ~n991 ;
  assign n993 = n1377 & n992 ;
  assign n994 = n917 & n993 ;
  assign n995 = n917 | n993 ;
  assign n1378 = ~n994 ;
  assign n48 = n1378 & n995 ;
  assign y0 = n33 ;
  assign y1 = n34 ;
  assign y2 = n35 ;
  assign y3 = n36 ;
  assign y4 = n37 ;
  assign y5 = n38 ;
  assign y6 = n39 ;
  assign y7 = n40 ;
  assign y8 = n41 ;
  assign y9 = n42 ;
  assign y10 = n43 ;
  assign y11 = n44 ;
  assign y12 = n45 ;
  assign y13 = n46 ;
  assign y14 = n47 ;
  assign y15 = n48 ;
endmodule
