module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 ;
  assign n190 = x64 | x66 ;
  assign n498 = ~x2 ;
  assign n274 = x1 & n498 ;
  assign n381 = x3 | n274 ;
  assign n499 = ~x4 ;
  assign n425 = n499 & n381 ;
  assign n458 = x5 | n425 ;
  assign n500 = ~x6 ;
  assign n477 = n500 & n458 ;
  assign n479 = x7 | n477 ;
  assign n501 = ~x8 ;
  assign n485 = n501 & n479 ;
  assign n497 = x9 | n485 ;
  assign n502 = ~x10 ;
  assign n137 = n502 & n497 ;
  assign n138 = x11 | n137 ;
  assign n503 = ~x12 ;
  assign n139 = n503 & n138 ;
  assign n140 = x13 | n139 ;
  assign n504 = ~x14 ;
  assign n141 = n504 & n140 ;
  assign n142 = x15 | n141 ;
  assign n505 = ~x16 ;
  assign n143 = n505 & n142 ;
  assign n144 = x17 | n143 ;
  assign n506 = ~x18 ;
  assign n145 = n506 & n144 ;
  assign n146 = x19 | n145 ;
  assign n507 = ~x20 ;
  assign n147 = n507 & n146 ;
  assign n148 = x21 | n147 ;
  assign n508 = ~x22 ;
  assign n149 = n508 & n148 ;
  assign n150 = x23 | n149 ;
  assign n509 = ~x24 ;
  assign n151 = n509 & n150 ;
  assign n152 = x25 | n151 ;
  assign n510 = ~x26 ;
  assign n153 = n510 & n152 ;
  assign n154 = x27 | n153 ;
  assign n511 = ~x28 ;
  assign n155 = n511 & n154 ;
  assign n156 = x29 | n155 ;
  assign n512 = ~x30 ;
  assign n157 = n512 & n156 ;
  assign n158 = x31 | n157 ;
  assign n513 = ~x32 ;
  assign n159 = n513 & n158 ;
  assign n160 = x33 | n159 ;
  assign n514 = ~x34 ;
  assign n161 = n514 & n160 ;
  assign n162 = x35 | n161 ;
  assign n515 = ~x36 ;
  assign n163 = n515 & n162 ;
  assign n164 = x37 | n163 ;
  assign n516 = ~x38 ;
  assign n165 = n516 & n164 ;
  assign n166 = x39 | n165 ;
  assign n517 = ~x40 ;
  assign n167 = n517 & n166 ;
  assign n168 = x41 | n167 ;
  assign n518 = ~x42 ;
  assign n169 = n518 & n168 ;
  assign n170 = x43 | n169 ;
  assign n519 = ~x44 ;
  assign n171 = n519 & n170 ;
  assign n172 = x45 | n171 ;
  assign n520 = ~x46 ;
  assign n173 = n520 & n172 ;
  assign n174 = x47 | n173 ;
  assign n521 = ~x48 ;
  assign n175 = n521 & n174 ;
  assign n176 = x49 | n175 ;
  assign n522 = ~x50 ;
  assign n177 = n522 & n176 ;
  assign n178 = x51 | n177 ;
  assign n523 = ~x52 ;
  assign n179 = n523 & n178 ;
  assign n180 = x53 | n179 ;
  assign n524 = ~x54 ;
  assign n181 = n524 & n180 ;
  assign n182 = x55 | n181 ;
  assign n525 = ~x56 ;
  assign n183 = n525 & n182 ;
  assign n184 = x57 | n183 ;
  assign n526 = ~x58 ;
  assign n185 = n526 & n184 ;
  assign n186 = x59 | n185 ;
  assign n527 = ~x60 ;
  assign n187 = n527 & n186 ;
  assign n188 = x61 | n187 ;
  assign n528 = ~x62 ;
  assign n189 = n528 & n188 ;
  assign n191 = x63 | n189 ;
  assign n529 = ~n190 ;
  assign n192 = n529 & n191 ;
  assign n530 = ~x66 ;
  assign n193 = x65 & n530 ;
  assign n194 = x67 | n193 ;
  assign n195 = n192 | n194 ;
  assign n531 = ~x68 ;
  assign n197 = n531 & n195 ;
  assign n198 = x69 | n197 ;
  assign n532 = ~x70 ;
  assign n199 = n532 & n198 ;
  assign n200 = x71 | n199 ;
  assign n533 = ~x72 ;
  assign n201 = n533 & n200 ;
  assign n202 = x73 | n201 ;
  assign n534 = ~x74 ;
  assign n203 = n534 & n202 ;
  assign n204 = x75 | n203 ;
  assign n535 = ~x76 ;
  assign n205 = n535 & n204 ;
  assign n206 = x77 | n205 ;
  assign n536 = ~x78 ;
  assign n207 = n536 & n206 ;
  assign n208 = x79 | n207 ;
  assign n537 = ~x80 ;
  assign n209 = n537 & n208 ;
  assign n210 = x81 | n209 ;
  assign n538 = ~x82 ;
  assign n211 = n538 & n210 ;
  assign n212 = x83 | n211 ;
  assign n539 = ~x84 ;
  assign n213 = n539 & n212 ;
  assign n214 = x85 | n213 ;
  assign n540 = ~x86 ;
  assign n215 = n540 & n214 ;
  assign n216 = x87 | n215 ;
  assign n541 = ~x88 ;
  assign n217 = n541 & n216 ;
  assign n218 = x89 | n217 ;
  assign n542 = ~x90 ;
  assign n219 = n542 & n218 ;
  assign n220 = x91 | n219 ;
  assign n543 = ~x92 ;
  assign n221 = n543 & n220 ;
  assign n222 = x93 | n221 ;
  assign n544 = ~x94 ;
  assign n223 = n544 & n222 ;
  assign n224 = x95 | n223 ;
  assign n545 = ~x96 ;
  assign n225 = n545 & n224 ;
  assign n226 = x97 | n225 ;
  assign n546 = ~x98 ;
  assign n227 = n546 & n226 ;
  assign n228 = x99 | n227 ;
  assign n547 = ~x100 ;
  assign n229 = n547 & n228 ;
  assign n230 = x101 | n229 ;
  assign n548 = ~x102 ;
  assign n231 = n548 & n230 ;
  assign n232 = x103 | n231 ;
  assign n549 = ~x104 ;
  assign n233 = n549 & n232 ;
  assign n234 = x105 | n233 ;
  assign n550 = ~x106 ;
  assign n235 = n550 & n234 ;
  assign n236 = x107 | n235 ;
  assign n551 = ~x108 ;
  assign n237 = n551 & n236 ;
  assign n238 = x109 | n237 ;
  assign n552 = ~x110 ;
  assign n239 = n552 & n238 ;
  assign n240 = x124 | x125 ;
  assign n241 = x126 | x127 ;
  assign n242 = n240 | n241 ;
  assign n243 = x120 | x121 ;
  assign n244 = x122 | x123 ;
  assign n245 = n243 | n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = x116 | x117 ;
  assign n248 = x118 | x119 ;
  assign n249 = n247 | n248 ;
  assign n251 = x114 | x115 ;
  assign n252 = x112 | x113 ;
  assign n253 = n251 | n252 ;
  assign n254 = n249 | n253 ;
  assign n255 = n246 | n254 ;
  assign n256 = x111 | n255 ;
  assign n257 = n239 | n256 ;
  assign n553 = ~x121 ;
  assign n258 = x120 & n553 ;
  assign n259 = x122 | n258 ;
  assign n554 = ~x123 ;
  assign n260 = n554 & n259 ;
  assign n261 = x124 | n260 ;
  assign n555 = ~x125 ;
  assign n262 = n555 & n261 ;
  assign n263 = x126 | n262 ;
  assign n556 = ~x127 ;
  assign n271 = n556 & n263 ;
  assign n557 = ~x113 ;
  assign n264 = x112 & n557 ;
  assign n265 = x114 | n264 ;
  assign n558 = ~x115 ;
  assign n266 = n558 & n265 ;
  assign n267 = x116 | n266 ;
  assign n559 = ~x117 ;
  assign n268 = n559 & n267 ;
  assign n269 = x118 | n268 ;
  assign n270 = x119 | n246 ;
  assign n560 = ~n270 ;
  assign n272 = n269 & n560 ;
  assign n273 = n271 | n272 ;
  assign n561 = ~n273 ;
  assign n129 = n257 & n561 ;
  assign n276 = x110 | x111 ;
  assign n277 = x108 | x109 ;
  assign n279 = x106 | x107 ;
  assign n280 = x104 | x105 ;
  assign n282 = x102 | x103 ;
  assign n283 = x100 | x101 ;
  assign n285 = x98 | x99 ;
  assign n286 = x96 | x97 ;
  assign n288 = x94 | x95 ;
  assign n289 = x92 | x93 ;
  assign n291 = x90 | x91 ;
  assign n292 = x88 | x89 ;
  assign n294 = x86 | x87 ;
  assign n295 = x84 | x85 ;
  assign n297 = x82 | x83 ;
  assign n298 = x80 | x81 ;
  assign n300 = x78 | x79 ;
  assign n301 = x76 | x77 ;
  assign n303 = x74 | x75 ;
  assign n304 = x72 | x73 ;
  assign n306 = x70 | x71 ;
  assign n307 = x68 | x69 ;
  assign n382 = x66 | x67 ;
  assign n562 = ~n307 ;
  assign n383 = n562 & n382 ;
  assign n384 = n306 | n383 ;
  assign n563 = ~n304 ;
  assign n385 = n563 & n384 ;
  assign n386 = n303 | n385 ;
  assign n564 = ~n301 ;
  assign n387 = n564 & n386 ;
  assign n388 = n300 | n387 ;
  assign n565 = ~n298 ;
  assign n389 = n565 & n388 ;
  assign n390 = n297 | n389 ;
  assign n566 = ~n295 ;
  assign n391 = n566 & n390 ;
  assign n392 = n294 | n391 ;
  assign n567 = ~n292 ;
  assign n393 = n567 & n392 ;
  assign n394 = n291 | n393 ;
  assign n568 = ~n289 ;
  assign n395 = n568 & n394 ;
  assign n396 = n288 | n395 ;
  assign n569 = ~n286 ;
  assign n397 = n569 & n396 ;
  assign n398 = n285 | n397 ;
  assign n570 = ~n283 ;
  assign n399 = n570 & n398 ;
  assign n400 = n282 | n399 ;
  assign n571 = ~n280 ;
  assign n401 = n571 & n400 ;
  assign n402 = n279 | n401 ;
  assign n572 = ~n277 ;
  assign n403 = n572 & n402 ;
  assign n404 = n276 | n403 ;
  assign n573 = ~n252 ;
  assign n405 = n573 & n404 ;
  assign n406 = n251 | n405 ;
  assign n574 = ~n247 ;
  assign n407 = n574 & n406 ;
  assign n408 = n248 | n407 ;
  assign n575 = ~n243 ;
  assign n409 = n575 & n408 ;
  assign n410 = n244 | n409 ;
  assign n576 = ~n240 ;
  assign n411 = n576 & n410 ;
  assign n412 = n241 | n411 ;
  assign n302 = n300 | n301 ;
  assign n305 = n303 | n304 ;
  assign n413 = n302 | n305 ;
  assign n196 = n190 | n194 ;
  assign n308 = n306 | n307 ;
  assign n414 = n196 | n308 ;
  assign n415 = n413 | n414 ;
  assign n290 = n288 | n289 ;
  assign n293 = n291 | n292 ;
  assign n416 = n290 | n293 ;
  assign n296 = n294 | n295 ;
  assign n299 = n297 | n298 ;
  assign n417 = n296 | n299 ;
  assign n418 = n416 | n417 ;
  assign n419 = n415 | n418 ;
  assign n278 = n276 | n277 ;
  assign n281 = n279 | n280 ;
  assign n420 = n278 | n281 ;
  assign n284 = n282 | n283 ;
  assign n287 = n285 | n286 ;
  assign n422 = n284 | n287 ;
  assign n423 = n420 | n422 ;
  assign n424 = n255 | n423 ;
  assign n135 = n419 | n424 ;
  assign n310 = x62 | x63 ;
  assign n309 = x60 | x61 ;
  assign n364 = x58 | x59 ;
  assign n363 = x56 | x57 ;
  assign n313 = x54 | x55 ;
  assign n312 = x52 | x53 ;
  assign n316 = x50 | x51 ;
  assign n315 = x48 | x49 ;
  assign n358 = x46 | x47 ;
  assign n357 = x44 | x45 ;
  assign n319 = x42 | x43 ;
  assign n318 = x40 | x41 ;
  assign n322 = x38 | x39 ;
  assign n321 = x36 | x37 ;
  assign n352 = x34 | x35 ;
  assign n351 = x32 | x33 ;
  assign n325 = x30 | x31 ;
  assign n324 = x28 | x29 ;
  assign n328 = x26 | x27 ;
  assign n327 = x24 | x25 ;
  assign n345 = x22 | x23 ;
  assign n344 = x20 | x21 ;
  assign n331 = x18 | x19 ;
  assign n330 = x16 | x17 ;
  assign n334 = x14 | x15 ;
  assign n333 = x12 | x13 ;
  assign n340 = x10 | x11 ;
  assign n339 = x8 | x9 ;
  assign n337 = x6 | x7 ;
  assign n336 = x4 | x5 ;
  assign n426 = x2 | x3 ;
  assign n577 = ~n336 ;
  assign n427 = n577 & n426 ;
  assign n428 = n337 | n427 ;
  assign n578 = ~n339 ;
  assign n429 = n578 & n428 ;
  assign n430 = n340 | n429 ;
  assign n579 = ~n333 ;
  assign n431 = n579 & n430 ;
  assign n432 = n334 | n431 ;
  assign n580 = ~n330 ;
  assign n433 = n580 & n432 ;
  assign n434 = n331 | n433 ;
  assign n581 = ~n344 ;
  assign n435 = n581 & n434 ;
  assign n436 = n345 | n435 ;
  assign n582 = ~n327 ;
  assign n437 = n582 & n436 ;
  assign n438 = n328 | n437 ;
  assign n583 = ~n324 ;
  assign n439 = n583 & n438 ;
  assign n440 = n325 | n439 ;
  assign n584 = ~n351 ;
  assign n441 = n584 & n440 ;
  assign n442 = n352 | n441 ;
  assign n585 = ~n321 ;
  assign n443 = n585 & n442 ;
  assign n444 = n322 | n443 ;
  assign n586 = ~n318 ;
  assign n445 = n586 & n444 ;
  assign n446 = n319 | n445 ;
  assign n587 = ~n357 ;
  assign n447 = n587 & n446 ;
  assign n448 = n358 | n447 ;
  assign n588 = ~n315 ;
  assign n449 = n588 & n448 ;
  assign n450 = n316 | n449 ;
  assign n589 = ~n312 ;
  assign n451 = n589 & n450 ;
  assign n452 = n313 | n451 ;
  assign n590 = ~n363 ;
  assign n453 = n590 & n452 ;
  assign n454 = n364 | n453 ;
  assign n591 = ~n309 ;
  assign n455 = n591 & n454 ;
  assign n456 = n310 | n455 ;
  assign n592 = ~n135 ;
  assign n457 = n592 & n456 ;
  assign n130 = n412 | n457 ;
  assign n593 = ~n245 ;
  assign n250 = n593 & n249 ;
  assign n275 = n242 | n250 ;
  assign n311 = n309 | n310 ;
  assign n314 = n312 | n313 ;
  assign n317 = n315 | n316 ;
  assign n320 = n318 | n319 ;
  assign n323 = n321 | n322 ;
  assign n326 = n324 | n325 ;
  assign n329 = n327 | n328 ;
  assign n346 = n344 | n345 ;
  assign n332 = n330 | n331 ;
  assign n335 = n333 | n334 ;
  assign n338 = n336 | n337 ;
  assign n341 = n339 | n340 ;
  assign n594 = ~n341 ;
  assign n342 = n338 & n594 ;
  assign n343 = n335 | n342 ;
  assign n595 = ~n332 ;
  assign n347 = n595 & n343 ;
  assign n348 = n346 | n347 ;
  assign n596 = ~n329 ;
  assign n349 = n596 & n348 ;
  assign n350 = n326 | n349 ;
  assign n353 = n351 | n352 ;
  assign n597 = ~n353 ;
  assign n354 = n350 & n597 ;
  assign n355 = n323 | n354 ;
  assign n598 = ~n320 ;
  assign n356 = n598 & n355 ;
  assign n359 = n357 | n358 ;
  assign n360 = n356 | n359 ;
  assign n599 = ~n317 ;
  assign n361 = n599 & n360 ;
  assign n362 = n314 | n361 ;
  assign n365 = n363 | n364 ;
  assign n600 = ~n365 ;
  assign n366 = n362 & n600 ;
  assign n367 = n311 | n366 ;
  assign n601 = ~n196 ;
  assign n368 = n601 & n367 ;
  assign n369 = n308 | n368 ;
  assign n602 = ~n305 ;
  assign n370 = n602 & n369 ;
  assign n371 = n302 | n370 ;
  assign n603 = ~n299 ;
  assign n372 = n603 & n371 ;
  assign n373 = n296 | n372 ;
  assign n604 = ~n293 ;
  assign n374 = n604 & n373 ;
  assign n375 = n290 | n374 ;
  assign n605 = ~n287 ;
  assign n376 = n605 & n375 ;
  assign n377 = n284 | n376 ;
  assign n606 = ~n281 ;
  assign n378 = n606 & n377 ;
  assign n379 = n278 | n378 ;
  assign n607 = ~n255 ;
  assign n380 = n607 & n379 ;
  assign n131 = n275 | n380 ;
  assign n608 = ~n254 ;
  assign n421 = n608 & n420 ;
  assign n486 = n246 | n421 ;
  assign n459 = n311 | n365 ;
  assign n460 = n314 | n317 ;
  assign n463 = n320 | n359 ;
  assign n462 = n323 | n353 ;
  assign n466 = n326 | n329 ;
  assign n467 = n332 | n346 ;
  assign n469 = n335 | n341 ;
  assign n609 = ~n467 ;
  assign n470 = n609 & n469 ;
  assign n487 = n466 | n470 ;
  assign n610 = ~n462 ;
  assign n488 = n610 & n487 ;
  assign n489 = n463 | n488 ;
  assign n611 = ~n460 ;
  assign n490 = n611 & n489 ;
  assign n491 = n459 | n490 ;
  assign n612 = ~n414 ;
  assign n492 = n612 & n491 ;
  assign n493 = n413 | n492 ;
  assign n613 = ~n417 ;
  assign n494 = n613 & n493 ;
  assign n495 = n416 | n494 ;
  assign n614 = ~n424 ;
  assign n496 = n614 & n495 ;
  assign n132 = n486 | n496 ;
  assign n461 = n459 | n460 ;
  assign n464 = n462 | n463 ;
  assign n468 = n466 | n467 ;
  assign n615 = ~n464 ;
  assign n480 = n615 & n468 ;
  assign n481 = n461 | n480 ;
  assign n616 = ~n415 ;
  assign n482 = n616 & n481 ;
  assign n483 = n418 | n482 ;
  assign n617 = ~n423 ;
  assign n484 = n617 & n483 ;
  assign n133 = n255 | n484 ;
  assign n465 = n461 | n464 ;
  assign n618 = ~n419 ;
  assign n478 = n618 & n465 ;
  assign n134 = n424 | n478 ;
  assign n471 = x0 | x1 ;
  assign n472 = n426 | n471 ;
  assign n473 = n338 | n472 ;
  assign n474 = n469 | n473 ;
  assign n475 = n468 | n474 ;
  assign n476 = n465 | n475 ;
  assign n136 = n135 | n476 ;
  assign y0 = n129 ;
  assign y1 = n130 ;
  assign y2 = n131 ;
  assign y3 = n132 ;
  assign y4 = n133 ;
  assign y5 = n134 ;
  assign y6 = n135 ;
  assign y7 = n136 ;
endmodule
